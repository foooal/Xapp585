`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZnH/MdsD7q/57234Cl62V0aziOXrSWtaOecgtEFBKoAjB1uU08GqaHtTbZOGqsU1Idg2T2s5t8uo
5MdeAUC48Q==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zIxG8ngo2pqNq4wqKPYYh2HaoQdN6vAvjqpmYZ3uXy2Tprlj3Lb0MCAyu9wN7vPf9ZXaPythXTul
dMQu9KCW2z3GRzWYoYk6y2f3SQqMX3t586UyXES4e+Tb+MqUe9wozPPANVHZegCcTzFaj8wvVdVo
pZgxr82lKIl8OqKNvi4=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
k3BHjKiWdqNtPNV7SM4w1K8nS7g6tn0nQ6MkLFZW5q3++f4VB7mfDN8Lo2Y7HmO/HEAzF4wRwTQV
op+YdAf1FKS7zwmOv4RYxNmZfMT7UB7rugmodeYHCMsEDp/91QBhXv8j9JKRZexPvuODKt08oJFi
y2iHgRNdRHlqNBsc6+Dgxpyv3qcBk0eUxa87sT8hYhoXuG54UBP4U1pPF54lCKGIvH/JLf7MxZOQ
E3tQOcCoG8jOQCi6VLQ9E1i/HTNie6E+6K9cpx2SdKsLggadJbKwlGU0Iz5Grc+jjfNW0mExGUHl
7t33kYhEsbw2LrxCx9iUGUyWyssgUhY4PvLbkw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FYGyy1WGIyVSdzMVsBmPHdNuz2ZwzX1qWik/O9mxmZtHKlxwi1gAvQrtwl8VscV0a5RJfIFUNCN5
LCf3iaYntis4U4U/OZ8G+g49CxvbQFacl7LY2b2//CTY88MCE0dVJj59+scRJPwIrgixoxiFddsb
l8Yife9MTTHnArG3IJxxAIsgEsP+4kbmrEYnmyLyxCOsAvm26ADsxq4O9e8yGWdrI9VARnhENoZj
BFeIzJq6XCff4hJxRClEQkdv3XXkeLcweOU9QyzNFckPx9vDEZW+EwFMo/kxkRCeRM7wdGybJI0A
AT4xg3T6bDEkeuWFIECwb1d8Xjfl2md2+BC+Rg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qpZA7ND5z8Gx2tha1ayZfOtsQUfbcWcYUyVmGRTTK4K1iiHCwZynNpEIykekQtqe3n8oodWZPv5y
k6F62YsGKt/PxQ/YHoxTcd6uY7kG0Ek/ySLuRprUKHNIuTXwmD45ePTFgMKEqYPWRNFNxI6LKRW8
x7OR95Y2pFo9mc200SGV+UmaGpXWwWGJtSt7h3c+64VhnDLXHgkdcpnJBQcTFB0MIrBGvEh8KoKh
nmkRYvA75qM7csX0Sx4ns5ZZfPbt/iGipZZlpcA5l7grVEX38+FpBNaGW5WguIuPtjLerkSW9xNZ
Cwkw5+rPhVUBPzKyrRQp9Z7Cc7IkqGq07LxWCw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DFZU/TcA0Lxg+lSAdm0ljGuM2/gn/hRLwFWjjY4z8Rv87JqR3kg9NtQ7zyUnJETkLli/TEtaf8rE
VkfepNMm4xL8mu31wVw+jkR9LWscCrBbghGFZo3JxnEaL59zLrfTcCjDNM61WbxCqjX7IPeQU1iY
IyKNxTlRE8nSkW6gwxE=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kiAIS895994Vs0abURhvrUvD/d/yNkCTtC+beXSKiBQ/eMS/mAY6P9OJKNz/iRQfQq0scHi19BmJ
uVJMYr7WwRaxyo+q8pd6AFer7FyQJ0pIR9Uk+Rs8t5q2cAzUMSiKU12i7EFpoDcXLVrEb+eIJOYT
izOkKpKj1w6W0EZ95e0NPReFAvrgkanhyWvo2g+Nhbz40m2WlaRuPnZ/lF055UpUUNBYx6bD7TGs
+9vssIS+swsfvT0MaajoHr6WoaCDTo30D68UId9+pBhXAatBRn6kp1y8TADsctcgC4cgKoS+MfYO
ypvqibZPFuOJLf3w5nCXPqce3YdagQ0QKswJBg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1798864)
`protect data_block
4QNvDAmafR/vK4plCqiuYQVSLs+SxwE3L7oQMggr8/aO8ILTEsq+WR/QfeJe+nPlkdoTfpXcsJeA
Se9ua6IDH1V2wj5j6AjBN8Dq4vycr+5qVd/+7afKd/5YiC4hvObc3/cYmae6ixG3Qp5vwEIofEc0
9JEAHJ4l+te0aWUsxSAvfI6VxYv5ZQ1UeKCtuRoA8l8r3JEvqyLEWI0mmFpfiJC2MG5zNjtF0Rm1
Tuuocr99VJC9vWqxRGgE7OwdT5EjklxC0U8SbuO/kTCV+c/80VPiLO1tpOr20PQBTwlCzBuusphO
PNQik1UtBcsGFYI69aIICMeDF8lEAqqzJxQ4B0O5UqcddZSTpYEgoUhFcsWH6uDNwrV208wHcOaN
5quU+vKdDwWd7nTaMIQyFTTIIv7nser1zhX/cdhoV39pb/FjYgAjbsv9fLltW4H9nxGDWiI8sAVY
xUUoz7EQ2HJNU04shvOGODWQ8LgtuWdHxol4vQFNrIWbm5heVs1P7vDgFnvq1vDbGB774mDgdwpK
bIWjc7GBIWxuQQOcsTjmQ/fw1P0P9Dat0mkzjrfWwcPKUbTVrNkNPQyuTrDhs/gMHIS5+Xcb9dI6
UxqE02SCQqOO9QYjF9bL8l7+BBZyjLSCSO+WAqSVkaNCaJfmpAEt8C77gfwdZVQUXeOm7uxL10iz
S+UwVN5e1w/E9pCf6pNhEBz+xYubW9NP4sgSPc8u9itdy4+3bXEBvLrbFHMz5MoanvACd5Fi8w0m
cwqri6JJ2E3SAP+FqN3zAwkrZmbtd6q1xpcKjLT4BSaFKdmDRk+A58V1+KdbV/4sGrm6D/2HjQ0p
qKf1l9EhS4PgaSTGkJPHLmxK2x1GDGFPJFHFvlAy224/921mMjVbFW5noJunBYqwlTGSZqSFtd6s
OQwd3wasyu/7uuU4IjDjmu6j1gyaVjgb9kZDWC2yklj/i6wRW716tlxMtA7+d08wtlBmcPwRocHR
Ca2bh6bNMDUBNTy8piQbu5i6OlgQte8+5xpxRm4gPEx2IBN4B79lSrKTmGDX4t9MWYbRiyRY+bVL
Ah2MtCV3yRsqGPUHa7/NuDfpWj3wkUDsqp5sz+RZEMGoSZ1n+dttVdgJV1LoPYDccVANdAF/tLvL
jJwYqioi1JAEQ/9QBKk6FYQrTli4dj85Okiut6mBxAglSc50BTnUzQftwePXfuBdFU8RSyJuqAZY
ADvIDO5IF85nVm9i26zvEqL1mmGcTG8ckiRXPkOKBIVNom9ftFHoIHBUcPI3j/HgQ58If0xrsuiH
rP5PWFTIdfcK8BFvtq+YvnSaSWHcGDqkXD4K5AaHBwc3yguDsoBGwK+UzVcZSYOGFgMu9sIKqape
9kwbfycZYzeLxrOQ+LOLy3tzJWmPZv7m5B3ERvViGySG649Kjza2PmBfZJBjNzSDsS1+FQ9L1C1T
+hv2BzyMh1wrG4DNI99jj6D8XMRw4rS/qoAaUjQ2lh2D+IzaxeMwy3niZBNn02scF0cehsRWM6vC
rbJvtRYFx0f82yG/WdwIKbyUD+qCXvg6aSVBE7DlJnxt8mYrZbQTBphNfgxVtOMmBaTYkYHk7PLY
CDZPwemfFs5rdMH3y5jobO3gs7dPoIcYGjgFDf8RUdQuwkvWuLSnWs5sn4MKZt5En5TS0vX/cS7H
pwv56GyobgLWmMGiJy+YfiO57+hjaGOtf4TdWIkOdULsdlI6dGLPj0s5DXNW1QfVZ/rTP+v4i2T2
+Fozu/SN/YgBFLGdBQBKZlRlCy+39DSnkO8YlhIlkw0d/3TPBnKtYRRdeO5lF9ZP8VP0u9pDW2NV
5O7c7AYnbgBNzcLW3AXQWRr09YCjCLUCmEyLHfB4AZiE1C80bsXJ7QFXvD4xfisshPpeIEjiJ26i
HGU4RAajlHmSgbFtPsmwwIMwZROUYxw0W/o4zCjHUImPilqXI+e3sYI12kHaKznGt7EOP1K48eiw
tesf/px4SHy6XSFoYI5JQyquka/syxdN4EQ+BCv0j45TBQ9YyBH7vxnyKrbVHJgxAsElhSqeo2XT
cMKik9DOYINtCx9EBd6mionrtcMsHiy2E0RNY+LEQ6O9tVOLYX6PpDSJtytkey9rg5cvNHgfSTJv
cwuPxwztEudX2oWJcuUBI89ckV1VwkR8Fk1wXvBcczActAR1XsIm8v5nyGUsGdUgBlLnqtgPUbrv
ifh3nj1uBPD2NU7buFKZGHs5c3FugrsyJeVKjZlmvo5hk6e8BQUvN5ab9DEzKdtvUsytsmQoyO7H
E83rpzBu+SQspdIHm1fQRtRjejcM6BIX2PTXADVJXCWdAzZBOc/82cl394jnPcXHIJNBK/psHN55
h6o0Fh2fMV/u1/ANn/cdrQ53Un18OIN5OCuV7lpVN44Q6yMkYcdH44pNM5//IuosOmzSDQkGQiBP
AUXlL6dDKFLDWhhUIgDexBzhj2nb9KNPVRidWARHvOVfHtxe2lYwhGc4BGyhfCgxrxD2udDe6wgt
cGxtMvVc0hgXjWhCM8bUu2koZqw9PJwikH8LXbuQszcLF9GgQXav24jUd8ApcTboPmRR8Py6jrcJ
Bus3fB0NReGyYi7kU1axu48kmc0xJ1IOnPHAbw/85EmhdvmqnaV39f32OG7sa96T5kiZTwmlsabj
9cQnCVE20TICRKMnxmAb5xo/MK5JeQTfO4FzxE0tKZBMuvTLBRDK/dX0xOprZnK+px+Mlm0ADj+r
dm1P9ai5eQe3WkOK7oAe0ftzlJkaa6o9pUqJ6SQH/fNWRcyFvbQVvOJ/APG/TBp5e3mGbhAorJ6y
qcsbTQWWWNTKCAGExT74DjRwOM1F3Z4du7hBQS62ZEIvq45hKCeuf/t5yCqhrfC3xFx2pZ8PW+WZ
i9vineRHcBbAQieQsc1by53r/V2RPEVPxUKtCz8tF25EnYa37vT4WK0ZKo7CmNBnmktXvpb3yaS/
lwLr8IwxC78S959zwjfosbs9CFBC6xkVkdl7O+G9AbYzQFWVVyYq0l3tTjLMemWbSBeUVE8JoZbu
CP4ukghbgmiPWS15lGJtTNYCpqooxaqjty4NAlYSAQjcHl2H1fBs5vCr9DvCSLoDuRbM8k68wvGS
e7uwcGQApeD3nc34E/0gtMBO+DTuoGP/jMg995VRViCDj9TzenrlJXk79+8Y7uqrYY3NTcmzmxaP
LobS01FQAYziezKRjL4k6WESNDWWVvZClo7+F6gyQiSKCeKtuOqr9roCNplvMHVrrRAS04QjIuaE
u6aDD9KF1WlargapesnObpJ9W1gLwVCwvjgogsS0tyfRCLPf3y59jkt3AKq5legVWzq8dCVjcN0l
mugq62ro+JtJPHj4WKXHChFxwYXLtqMHgOzGMlp2lQCERyJ5fplnFV9zJ/lmy6JMDezle3mqC8zv
RC83MOBY9EZ2BMpR55RoBHcYAqCsv/7+FHfkR/U4CZ2n6eyFMoXhj5D7S1ecFNO/Mgs2t5BOpLBh
7o/YDAbJqwvQjoO5nS1aSrI6TOxroi9UehkQxvL0hMYmr0TBAxr51toh9U5dI4sBYBI3aKwFvc/G
dCG3utI1q0uR7QqgLDf5J01RzNNcrahn1e9Euo1QeTK1VN27F/8tCYfBrA2Gd1b4jlj7MXWGKWA5
ypHu+MBCJAIv+ZPAxE0xVyY9ws23QwTPa15ZybS7RCiAv+RciluoBsQ2coGIx2kVUFVOzj2oHWdJ
yaXfkw2QcVAjXEapWZycyj+rOn6PlFuKot/uEEciFG8WpcfJ3OSYarZl6HD+IOkg7kMT+A6Eb7Q8
N3DWm9gHRRvRpVnzGdWoqTYpWSras9uvKtfWNRAGpf5e4rGKGj5n7+XNqXNcWKENeljyzln/kFwa
qOS1/fRuEdOaL32hbWCf0Z1Hf8iGJvzsjaidG2DTU3OwJF+HfudM+wM0O8fU2t2ZLc8lgTXL0qbh
tZ3ENkTkrHOUPSIBEOxfZQGqEkwWwCOJ1juadOGAW2/CRe5TmLF8AvXVBvw5eJ43K2J5haqlwBzq
VLbgqp0efI8Ts0i6o39JOKz5bZsSGES7sn1wVTyjq+LsTSxyPy3eTw8ezck+mHn9Ry2onPoC0Yf/
MWyeulTlbb4V+Rfwklu4pTxuKzOwQsncW1411/I1dpGx8O0F95DiJthSTpOTea+VHJgbfb6NfP1d
smFS5rYwF83HqYhSDNXMqpqFmNSl+kzCy08TwiKmazHuVsNxI/Yfb6q1pdgKdG2EZomYYYzGldVa
hTlZpzh16tzY18Lyp/9Yd9hHsR/Ijft55QuXjl368HvtYv55wCuz0vCHFHaVyO0HFwJxo3cU9DBe
t/toPkkgJ7OxsnCKxasVk1t4tLqYr3T3U4wmS2m0RHss/zwMp6ZfYqlHMHGP44IpJ5Dl2bSCt+52
+CHachyOX141DaUUGK90Q5MoDWfaG717xQiQ891GALcE3IzJvHqY/SQqjfaOr5upYGCXTWq0wOk7
DnO6+9229Lh+ok9ZBeT4FSoyRbo9NYDPr8QwstvAPuNbGaQksZoDkRmZgAucJEkbYZR7wHkaqF7a
E64rjKG1kXj9LnnbIWpJbBrZZ4C+64iXI+puE/Fp1q3Ws+LJxZDMsW8FpKJ8OrdIt/Ctf8NyjDWw
44H/nhbBT+PfF3+Nmk8rNGSRx5QrpPgoJlj8ZnS6vfmDh854NIwndbbJrrUatOl1aIRFWHKolidU
5RAZ2Yc5xnUSiq3zIYMWLct61bzTWhpjiV833OYR/C6tKkDL8R0i+jhpmttl9PIidqlw+yLmo2e6
NAiOgUKgqRxe6p2a5zF4w3Dmih1ClClBW4+rQQeqc1FLClpiIIhCSxubmGHCmLUblnB5yleNpzd/
FDFh+i10xrCaKV3k5Pgnv33BLUNqVD6oJhX6Ll9huCRyQFDugaWUJPVUi1W/75nsEbPnFs3Vywf9
wRE68IJDWUn1NuAJL6ZB/f8kzNoo5OdibksPSnNHL+eByVOLspN1suEO49MQhVp52YM7sL90eppl
4oLugcLR5Fr84U3mJVtwKEXl0NwPKIoNfQa7pkFFo9b+MfXXRfGNyuBhQxFglbJSoTYZgAJANnoe
FjN0WRo7vedxy/vHL+gF7uj7kbbXsnBwWD1S2ka/AatE2RmzxUDV+VLmODZ2DcfJJDKOJE7riOGe
SIDm3ET48d/NDWiy0+vCA9CyiUKd+1QYaNpNEsDrS9Xf2YYzKUKRZpJom7F3N1Bso6KhEYVxQPwI
XHOwYykHj6jz2d+5G3ihwOCpy+htP68jYXdDofyp8lJ29NEEqmp8127MZv4Te36AKl0k6hRAdBPQ
VYgoEULTeowqALRCeu7bExkJ13ybOEIB/ckNUKFq/T1l6131eE562+J5cg2KOo744jkt4+GIJH3q
tTSI+3WCcwKvleIdqlBQKAGtKWHfnVVSuc95Y9Lp5fD9ZPwlXLK2N9M/rC1Bn6GJ/E8S0T4URIDC
eM2AnT5l/Rzjd6mhT4/omNGZpEOAJc9sFyr/2uiTPR8Drax55pSgtEl0l6LFwmWHUQQKlnG/z5mV
xvkstW6EWI4EUGyDEa6zR0SjvJwdNqlgFLiOWlB+Lr0X8FMyTEDi3kSF+iDGk8O/CJoQrDiobDlO
N6TglAGI+bQXA3EYeB2H8M9uaGVJd+QDjXnL9C8djgZGgWWkv/nZFQ7EpcUGPXIne1AIyEEVFY+B
o0FoxNA0INOdiwVEI7OY8uleiE4FOdN+v7Ud9nhJN0LLI6bJ+943y2h4Hx1ibZo7MQYQaetzHN79
8l0JZ3k+GDfGkP0ouBKcgWbedezyDDF6b6U9NQ+PytE5Mgb+cmSIDXMbrW9WACYXxpVtKJOi/3Gh
FNahn4mOkoXjXSQ5ooT1aKmD8LeAiDCs8Hco6ZvBOunGxgXGOOcyZyj4Ktg0Z8I3x7xitHEPtVbT
ioq8Y3dv6rFYkK+k6W3axANLXv5ihSrtoXvx/A9SgqanCr0vuUv72+84y5J8g/CImoZ89b172Wru
pZ5MhEymg67omg5xcv2O2Lz5P8f4KJyq1iMntdDu7HCPfu47TQUqS0z+eZbfgDk8jwQLlrTYJpss
b4iau5BzfIeP8+qFkUuD6acMzVhNiI2GCqzdvA67wPkS9VU+UJkXxNwrOc5G3mh7GcnF3ZC7SWZ/
7DR186jgtRtY5JT2Q0dFo/mZGyMq4cvQlShZMpByYm4ewKXXHyKimRqZaiddlvmcnsEkO0vPIRVz
e979izLaS/ESBuUG2H+3V835M1QfyVkl8rNaUaOXDYTMkU14YvyYARnB3kYb3bghCPTZ9KyW96Zn
g7mwgUnzxbjK+61YPq3CSk7aoJ71LePkg87STa9iKy8m+KcRQArQ/lBrQbJhaUlVdpmQ83uCq8DF
5jsn6+oD7tDwtEsOtkZ1aavSVxJMmTXr+6LddOLn+IVXjjn4e5WRhg8/QKuKYP2bWPmW1xP7UK+O
fvUuPKIXoli10tfcC9cu6YVdwLLhPrHiDlgE/x9LgXx9KHipKYX6UKSQHl2E/Ml5/FIvQYBUm3RE
RpaE/aqeFzD+2XEiZNKJSuhl2x48B2ijBSdc2x6tQKCVhTH5xtxgDrlr8otN96oYVuWu4F2VOgw3
wtP2kZCX9pezKfU9OyCfoWDDLWMuzpFk8E62/VPEYsWFTqgJWLGmYne5Y7LhTYn6q8Zv7/6WzJFc
LJxMSJXnZ3zhFWdjEIJ7HJmWS4Fb/ahYi6H+N0FOG111mLn0c3DQLJpP/436GYFD4zTG2kDjmex0
+4SyizgkUn3kPeqsnXGOfCX1BMFHF45udRn8r86NrkL2NpVMQ+8O+WWTysA5icXs7e2DAeoQ/+T0
iMbchhOnjJxxmNnDWm9r1FUuJH5JPJAu+MbB5HnYXQD+U/PElyuYx0KK5ZROsp63NBOk0kZiSWih
mqlLpWr9BaIcERxSrSLqalDjZukjhpqEu5nWR69tV4iwgzjKiu6bq568Ja+U+bGOXYIaTS9QVfGq
iedd1NPxWj/MDap5DCLb5TB/umrZKCl38yeQFMnJL5FWe5xt3uxTfk5jfn9xaqsfWQ/1CFzRH2Pj
J9RwuRAWg3wBZoJ8yMSD9+QfJfBPSf2HwQVHKNVa55Q873WTn7mw2SHeumfYx0KMRl8niQ9xRrrd
+As1VykNHJ53XtxxHHouBAqw3NpMmgu/lEaxabFAhpkQEzVKJqIm6jPDGmLF3sgAADmTY6dwkjTO
0yhFqk1nwexA/Oo9wADXwfZpUrWaAQYaolKIdg2TxFuzydMVm6y/wn0PwX/pNs4n6hn7l7upWwhw
Cdhrz3jsgSIFujIbVe0WRVoKuMzgX/fr5sj/Wt/TroP4ks4EN2kG1FfUpYFLPhEA60PlywFG7kiH
YXfphyd8yB7uYltssShVI0G3Ra+Rxi7H4UPkfSYI1LbW5chG9JZ4JB8Kza6bfKf0x5MieQaKD4Va
WkWOVnPHc74j/d2EzIVcl1Zbpf10qCqVWXUrVJiWRqxaETihIh1OODgj584kaPMqTt34LoeLge1o
522xv7TWKJvTnLUj2CxsJbUvxjp4UN9SDBaTgqJOj9W9GVMbZ0zjzqjcHqE5OLOa48BO7B4Fzj7S
75U7jPRKaxU9Vb6oRV4djP0W+6Xxo1OV971oV8oZmxGf4WmvWxb8nzDhhHC6QsfZ8tylVJ443Cqc
wMZ1AK0/X67MmUV7f+V+alcezPCfsA9O+bYX4ITz8L0NJHoUhmQ4FKYL8RXBwADIeitIusW8bZVw
iju+YgRecgmPEfUKSEjC/X0Q2cOJJH+aLgP8Wb4xBazAFjMFzDxRZ7dqEAua2O7T0Y8EVuobFz8a
Gyocy1RrjZP702fDM8aDVP5AQPREjM09M3I0EzQLZ53XwYUGnVeamEJS1MlNYRmcZMeui/Qh34+y
FyIB9Bv51q4wrJ2t/i5K8YDKGwdBo3xbiI7usHG6PMXzcpccTLwd+Oj1ZYxPL2sye4NUVMqLP9Uv
z7HzNTY/FBdtcI4MgFv7xvJ3fK/bfTpBTOjnjJB0x+0ShKKU9IKU8UMXfQqageo54jqCFgHBt5Tb
oIv23w9AZEGGUZcsCEYJZjNgke06R2kqjOkJO5kFZLYYWo3TxnJptqOFd0cu9FwDtfBrpMhRji2w
NknHKVMLAsaGca9CDgcA9F59ZtXZPkWWv8j6owV2vTHDIvHKL5/YuYCvxzjehmM1M3RtpAZi6uqo
tJgsWmKWKgmt76ug0nEF6fL57Qy2kCP+0LWwZln1j4n/9rfxxkKmMYjhyGF1cCAinohUiCYJJA3T
9hnghiOvG8c2VeYLsS5KPsx8+Wsqj50JMrhd/ufcB0ArIARJ43ZMmZUGoh2leTdBr/Ou9EL5nmQJ
qXythGfDb9VknIxr06F7hrJ5reGvR9C298v6gCLZk2EvrbZAG+gxpDCXNzCMNuDMtYGgQ5ohX1RG
PoEIpBXiiZ5AikTWgkX21xagYv+ZmExc5LZdJi9AoKfHeNnkwiZl6L4KAcMaEROxFE3WqpIcgzDw
OAdoT50V2m0e5SiiPz1M6/ZZEIed9YWRY4VRfuIXhgHBfik0F1HzV7XUz/muVI+JLAT1r+BlxZRB
kTwVI04xdihIFjNrvka16GMhudEzKQzlXmvVs3mC43dE83ah1MQ8ujQqHLpahliQPiyezNIW+3Vh
s/JkOp4VxWQ65y4pzvqMqHxnDG0vqyTWFLvlz9BAAJGA4cmj2pAr3CQUAq/UHanG+P+QQL3cptr2
6fnlm/ejHbsqSzuUkEkXWHKSo6lZAv3LhCcb1NNoySX/kbOFkJNsh9K5qVui+PsC79SrCnByj1QF
3z/RsipAw/hFJQpI/m232W0jA4JKfZZwDtJL6wxjHis0i0Yq/vRqo3IGcUmE4smKtNlUYytE+6jR
lBCygDIpAbzdH9QPXJYskW3mBAen9/2oh2q8nzqUM8rnJAD8h7QP8+H1A7Cx83nvtKJ8yevG14zD
qmEeA70fdWHr5Gmni24DsVmMb/FErUjKCWNelIEjzDq4yn6UtuUITiKUgT7IQKo4UVkafQIrLkg3
LANuolue42rtHPRCO4KJ82EmDERu2+cT5k9pOyaeon3K/yCY2ScuxNNy/qNjf5lXE2KeZ87d5RyX
LTlRIQyBfgR6Xg/uYrPZI6YHkN0kYXMhUzJpIXqTNFJeUJ4ndvtaCaTRkhvprbmPHKR2ep3vkTWM
9hX4axrTJlmWblp+bK74bowSdh2gDLaYxW6CK9sYYLvulOkwq4iMswdoUJUYK3hIb547Vu351M5O
hbQ+6ZScBJMUjFeomJfU+NaL0u3ofA85L5+GD/F/TaD1crL25KbDMd84VE4oMCilr81eDpJXwv1k
13c3U58F7cGKGDYBaRIq/BlGFdIiYJ4/S6ldgpaWC+qoZR1XcIU61K8RauuZ7HzoI0kOoryZw0nD
G39bVATtX3Btd7BnWUSGyd/RPO2cMV27myHgwY6cJs2+DeN/JRwbpS8lM7dEQkOFpOIyiT0btzjs
r01C9FJNA+lty2hP21Y0Hm1PJ9x8D3U13zGkoN1vSK5/WPBfetAs4vy9+Ax9nzgZedPZK8+H3muT
fcRYIEKhkU5LC/aDAT+jjDP821wmpngJJGbOpraU+7E8VmR6hZ/OgqcDZOIIgdotUGkffunAEqgE
lXENPair9YRaD/LArWDEpUeqyf+M9oF/CBCZ51QuioRdS3ijPcIdUjbPzRUqcVtmoFKDpCL6m5q5
+Y3MhwmT9NFPnNg8OVZyvlGZYMcpbZCVkZKUN+H/UK+SYPYIwdSavqU6B5pcBOGWC5WsesXG7eG3
oyYYTOSfaGp7LWdvcLLxWtzrmpf9+iqM/vbHJWDt0JN1pUtbYBvtIL2eOwh+V14jEO8GCGn7xF3R
NfCi5UWYbhJVdcB0+SHIiIm4VzsLi93ob+UuS3UhM5zbnmhpfjn0Ibew+3ETJawyVruakwRWKbDF
a4V18m6jgqZ/ykuOAMkxSYL1LmJZQf/qJi9uPXZgXDRJOo3DleIq8F5GoUQ73OVi/2WWFoVOBVW0
Y+Ulz0zkGSgJMSl4Ozv3cYjw6zcuymUX0+RqlSv49Nk0dsaeIwweWYbc67jkROyKMDKJuhJfV2et
kTojLAcHPBkiRlLandBmOLJ9MPoTPipOsITWAcWzo3yGS+yjc9giXbxr/QseGi5PUz+YBpXrUq+h
xNpBBhQL2XTUP+ludvNguT+9JTtljsBUsAQMSmZ9WVlPlTg9/arYYaP31LoJ8SBUKL9U8B62GufF
v5JmHQef64Uljw3/RalPrE60//J4smkEO6lvdwbOV37CUvh4JMQfA704GwgC00oMVD4CkP7V73cK
pSfJanXzcHfSUwRCm1lyb28Ac/0fXSxWbZPCyFn9whHJjvr68NF4gdTZs8/2qXuQshneRGXtVf8b
wRVsNn9ZDqsX2W4JgUlsm61GNv5FVwhOAUiyQDPOIPkn1bSsufLC69KuIGRe1ZeBJzybQNUGl3tx
msimjmwqWGw6VIxry+D3MclgreLAQsK+B2qbDX4uG2XZuNtWcHeDIq0nSvhTlzft++dp9N8hWSg6
Qx2HzXsluzot7ockMaswqoxfkLCDAAKlD2CpeRRFelSYu7/kscIXROiL0yYX6oQz7wW0nW2W3ZRF
1aTb8CJ0qHnby0zQhTnYaDVM/Q0KmWtrdqPjKlwuDEEg0ZGoWYVMwEetA1OLHHCIdjGlANC6WQS3
XYKykaUOFmDOhVNIp2NYo86ED2dp9GTJXUrHlh3lYpxZCNiEmneXjDU7YK4OBJjAoHMzAm8d42u9
5q4a6G4gCmH9zsE1uJfBHk59AZY/8y6DTF+T0M+N/lcvAGMA0RxscriZjB9Yb2vJzo76DuwDFRDZ
E5seXER61M1W11OFsld7sSUwvlKIX1Kbf770KPsS3IeOuLrWUqCf0hU7TFvmvkMYbyxglMG5hY+4
zG3B5YketSQerAUgLxNBXzpeMzyFZbe7LUHEy7v+BpxjJskVmvMgsRf2jTiigb9NX5k40EbHcjPt
rxYnXyEn3oFr6M43y8YgkwbEOlK1eYCuM6bwxGDcShDElzPrb1CM8ZcCVFQi+apxcNoaodrncpiI
WoxI4X5qpfYZu+BMMKZcq2noaVD26/PeeWzKuPVZe83TPTvRh6zyqQscGAvcgEwoJVqPqWVrymZU
Qbs/Wo5pFhtgPCnB4orN5ApNmuIYopdsFCWOh74jwOxDjoT/v2dWvoaTqle4fn9OA3cejSrt7sX/
BiQ22BTPiyRigiI5lcnhEy9iu+zPYOTTpjhqN/Kk3gB5T6+UexBXcg+GNeUld2PDdnC5o5etduNo
ctCXD/28o1nVVyv0XZ9Jc8vEf35mv+zh4Nl/c5ih/N1mvuIjGcu7EmzLSbsW8vr/XmOzCN3ayFAc
8afaltzfCDqtoeY/Be2og4Uzknucns/0pTDL7iZJLZ0jPYhUCLQ14LhA2foDvDK6bQ2opynGM28x
nP5/6tRtfsXPWZHoG4ZDuah+qo9GXA0oNE8tY276qXy8F9PJoH2+P3Iv7sdNaua5m2UFhsZ7nZDt
ykaDu3PJyCde73+Ky4Efdg7TMWWAux+Qa4AN3iHo5gHhKQeh3XAHxCPUx6gT2KthEmrNy/21w7SN
guAAUPTKk9HmOTi9jc9IPt+EuzJt8a18+Q++9qt309Uw63C5Fb2JH1jU8f0JH+Posfha5FNTMe81
QD8qksrAb8G42BZoyQ6dcLDwbgQVALl4hBpwNln4xBtQDIUHr9PEBuwS1C+Ah8RGQPtZkXEnD/YL
uqhIFpGdSD80K/UEo0gRjKRaIgUuDM+vf4qGK9vQjQWwDEy32m63yDMtAY3VPWFMRcqqpEmHc/Gu
bK4tC9tYitmD9NwOwMcoCS1XuZ0hKQ4wQzMcKwhKto3LBTkkyTRhrq8p/xDTiAqoCiseIWX8Bsm/
m+FnvhtMysO69MoEcZskPsfA16Dxi587j232BtNwaj6vZqbSyuxeCmLYMcH+YsfekoHIzZ/VzEE0
dm1V03NXtTC0pwAeqFc6n1mVSH1hVZKPzmxr5828pO0r86Tjgc0gUOgbIONNtPWAVRVnd/KiLwtk
N55fWHuFu1teeWo3sftKOYBHG2bh6r8Qmw2xk07mpRNl+d90Z8kNPZmrAm83gKbrI18ACtR82nc0
KAktRljqMUZGh2q/WlUrdi45yT3TnOqD3VXgcMxx9WPojzvrwdk3u0nsBofEvkbZqGDpy0JCcytY
tZiVeKLw8COAusH4R/Mc3JQuHDS+jikrf1X2z0tQ3lo1Nqyy/nF6/7YUdArhE4Rf4jt/uxYTo+/z
eOdtwDatOPenMCj/YRFV7UWf7m7/3R1Nf/e5D9OrLQ0rn07TNG31x0PenEZwsJ0E5zjZF232CwTQ
ogWZOpNPLg6CxbPwYY2TvZxRp9Ll0cU6JpfizgqeYlLVAHHSI5hlIao8DTmis+7B3IsoMQFh+Jc1
I8haM6TTxWquc1t9SXuR8JjpxaXFHRdopH5ZeyNawEGHQ3WI/9eYqyMpdD8NeDKfnxRG+Tj5TnRN
VsCRsosnkWfdjQ9lEHH9RT4SLC5jNEv/KBwBtuu+CiBI99oqHvMNzF538dUbQtrC1dyMtiDACDJI
QndT3wzjLAEaGSn3y2Jl6qyIfLCrIZ28MOKhudzDYH6IPUhgX2kR6DTBGMkubGWyrArZI6vJaWKv
mNx3kDk6aTbfZ6Dku36hi8pr0Xecatd7o4WfPjVeFyER+kiEn5taOXPg39i59NXOZzDUuPJyh3Iw
Ucbkl0brX51L/m7ohM/RPjsm7OIAqeKi8wX9x5KPuLwvqayv7oqijLVCqo24KHhQGg7LzjanEyg/
I+bt53emJzHmPvZ5az9GVrbJU3eUQVo4wHbr2eAys7MEZR96zHOkNKzXj0ykeenRcEuyzdvu+9pO
S5o9bGS927BmgHbg6Cthk2XXZHDhAH9rt+8ZrLHAYXzxt0oBRkTUPQM/e5r0FET36opgkmqn7T2T
DkOKgdCyOHi2//rMBjo00dVvIOo79PEi235G7pVkSbRSX5/ItMt2f7C+Yz4kxZjttSMQacQKG3hL
4XSCTRqvACaysWRorzUaL11P7EktS5/070KYkWQ6PYzSvUGzbj8YfVvzAk25IQsq/WAdIkMxin6H
EVuX7lPpCK1POjPxOOf/4XVdJIN1V1IRY6zLLCAlqxzHVTEAb9X8khEv7MsiaGdaFspvss1VsEzk
D8lvkNhNacs7UE5HHFxBBxbraLVXp6NyO1aX5z9+1io9abeD1Zj+hRYdyo/citrLHqJ+91bN187q
4ZSbReIYS7lzGL2uFL9gXtFYdYVbz/He9tSuZ73a6Zan5i9znHEQ9Fc85EY4PmDvBVyzSDZHl5r/
EUR4EpVYcItdahPKvHhfH+Hj5TfHMzsjdi6aZTCziH/TQpQXB6f/25Yn2eQApxZJg0bIVJc38rdA
uo0KkZGCVJYxaDenaRP/Nazer4+dIaaFvhu41GVVfkj1rwrWAXGGjvfbQa0BnTmjMtsbtHR+Vuor
vv91d+8+iOkXxd+77mVWo9+IjgDhCNOFGFt37HnvFRmoiYGp1NZn/Qyf4coVslLZzM9L5o8uHReJ
wwb7DXFDxk+YxvHF6zlDZvnWOg7z6w2etTJpXJ0zj2NiDg2+b4wWNPb+nATWrncQac4YViCqHPBn
zpPqmbEXBLgHRnlNK+xZ3IOTYfZi+aBuO1fMDT3Qz6sw5vet9+V5I6169IwlnvGAA3JhgJjZu2GV
HJMWKiJNgzJzC/pW941xNVYDwg4zSiLYXCCqb6PBM5OnQjUF2LO+8n0ohMBcLa5MJGs11/F9vO+D
jxmM+yCjkXNibxYqedybrhVNUIGpZg4hq7krms8DFsvGhtEmmp9Y7oy7PSnOe5PQ9XmzbeRrreIu
8xDhediSR9bgMaYeQK7timUFWxs7ASFH8FNPw+HgEXxql5JJlKXctD6+tPdJR4ANMQc81jv9pknr
BVbfy0JUVJ7ueNYNVHeqhl8eVahTwEpyDls6sEj0jGqH47gs5LsEUxr6LFraIpjB014GBsdVqdNg
EzQ21R8OHRe4ZeYp0YTF3p1NqIbAk603H8vYIvwl0M6RpEg95yWfrKHHw8a0O0muIOUmYwA9TVbU
c2EwPLv5VLYd8bzxzN4Y8O76iDGO68fAEOPd9OcnRyHmRu0HoknjBGL2NcTfhcUvzKNnHPd8pEJT
eLU8mp+DlDrZDBmtk9AAR95mbec2hjT1kyh0Ki1rMmTrEVNk+P27tcwK3TBsNSdqp5UqQIiZkPLh
9ZAOioOqR08PtAm4Br1cn0Pn6lNU/1blfEuiEdHgnGjNZpolVw5s6asCOhgmGtK8hjnHy/Ibj9u2
aULH0ZKnouiLdixFqV4jZiQUWXH0kwAF1XBuwuenhZFxoMAfgFqycFxWbpnf9lkfDZX9Nbt9FoLy
3nBJUTo40jKVl5J2HcMPRrKHkpi/t+ofilUWAcyZOQSGelX4vINa4QZ3kVBwNEGOLig0qwF4oSed
CapTVsAVVLcLxScHkavYVFgEjRUe6hOhN+TD5EfOlUpcDBAH6s5boU10pXw/68HQlATD1QqEPCgp
AoMCi+SMJbb6xMkK329hoM5Uz1yLZqc++e5BYUKLXQl1LcwKbWRNy6/xlR1uMxg09amyVL+dAe6y
go7Uu/RxwRmc6NBPC/6KbRxmxgKBNknbXsMKcDpcbJIElejPlXVrErkUsuZ7RO3J0U3ysh3HYVzk
xtlvt0qzXnUUh3Yc4JiOmtH6aQRx1ro0O9Rrz4almyTefrjUb4U8I8BTToVZ18X+m7UpVSsdst3s
WCw6YJ22P7uv5MZ3+i7cnfSW7kN3MZkc2iBcjRJFN/f1TDQWUeSgBOBs7nS+rwENtEXs0Jle1zF0
OZ16t3wUphoytvrDSv5PSiMOnt0XdRoivLgRFUXVE+dhwgftL8p2Lsq9MT8bkJRYo3A+FqcBPxfb
qsXBDFV/Eslg0+2xzZ8FiPnX3agtCsbVNwyX0b67FrMINQ/fG8ygvN4f+SRwNUvprP+sXTVFpwW4
A9lGlA89RHe78/QKA+niy/RVSIfr1E74oUg7u6R898LwbJfsmXvJJ5xw9KvPMjSzpfwh8dmBMi+H
11JPRal63erknmUY+8mTQ5m73DXfJ+ILNWN8OoTsOOOVeLw2/GipUAS+ff6cUGtf8h2pJopd37bh
o5JEJfhUcZXjSotnoBYixwra8fnBpB0lDrxJ+oNH1J+uhqtP2r99xl5tq5nvW7ifhMuteQnxi4MR
J8MRtKH75d7BvNxGi81KUriUwBkEFKszyYuTGsDKmO41wj2YoTN+h3Guudb7FTWU0PUgfEZ06+/z
wBovPXdLI2rCr5vqTOfXPGPzYlAD7n+LWkwLQObp7wA0sXFZiB1JlCJYytEOfg1nZMQCvAQolpfp
8rzjl8w0iYgmc1cFLJ1cD2dBNKz1x3KjNl1mloaedN32AHZYFuYVJBArK8UllW5Zd/ulpoFAjOaU
aeeDfZ3VrgQyNLiw+iHXM6cDKaWNlcyNY7sAPBEp1e2i5u1hslR7lrD18muq9Jfh3jWAmnBPgmhA
Qtmv8D4fJ7N56KxxjWak9GiGsQra6/+2SztH2xKXvAl/4UkxJUeUEoTq7H2105re54Bfg/Y0+MVQ
hi+d97Rmb2kScC+1fvQN51GMZdUoeBmwqUUYPLlwAA7vFTmii7CEHXTw+LR4cx9iDI+72iJD16hG
OdymF2JWmeCxhEWvJIh9MtZ66QDw3DW3jAOHr2OPWPwoojkxSyKVXMrkMBAlQbsWAE8DCntvcYpg
DFDcn8EzpBtmSmLAmhn9IfVl8gIb8k/LFVI+jQ7OE1YWTBkiuKHPhlY+0jBsKsqkFZgLe7rARtKm
BLOfNEWzmyTI2hMXK7VH/qvV0bZEny0L81f3K149a8yPk5avrbgxUh2ZsergqQeKvqagiUpCkzjI
BCnbtHhufBkIINyep5tGTQ6h1AoGOJt+VPZZiTgSM1WIgxKHnQ6mCOEcjVhCkTuQuy7fdpV4otmP
uR2t/BfB4Ru62LeHwwfQaX7l1u7KwAA2X+MpwYf3ks6BwiKkEwcaufc9NfgRrbOwzCUalh6tbZFz
MeVIG5460iMPJpJ6SLrIjqs2EeZJEJ5EQdlxJvOV4FUirphdyWtOg/B/me32plWc6zfouf4P3ukN
2P6K0MH2LDdOyKIOO+p6cr4/Dlkbfq9cTKfX88b36L5LaJyG2xOzJlTF+xeozrryP1yCd0g8RMd0
XQ7UOURt6Ynh0ZLd5WDZDpWGalfJgfIi5Xay3qXzdOYD1KIZ3h6Ow0QxM/CKxCSq2vFHiOPoMR8R
v3SIepHrNPzqZ6Qy+98jk1et83bDZVySq5Qc10Qq2EFpFumwmq/7DRsITtvT2q3MZopRR434jove
T2tSJ8PdtK7rWxvEC/v+P4MQkgClz2e2s9YBF7zi0NWuCSplFhZ/3ae/H8bRvJat2Zz9TT1NdDoF
sGNCB27c0RNVhMw8ekWgxQFDEFOoVR2dIMp1FWOHdTZwO57NlY9RPiPry1AwWlMIAyn0Tqgzppzl
MQwX6XY/vXutBLPGZkPANeK9Pql+oStuREMmZZvm2thx4uq/QxJDmRERxVlPlIm30KgaTqLvs/E3
J0hQCLsCpM39Nz03RQdCDZw0UyZxZUHyI2/YaO9ZgpyLcrm2NgnnHDErHcCNvdIHbQJFrUSMQXD2
+tqDUUZWtPQa/ppn9rGOGYo/TGoio1Tt5bg2x2rphr7QD8DjZfQT6cgv2npw1JFfVTiNGDKDOfmc
ZfTjdvQ4IJF5o+jUJ9DdiERo2Wt+iWzRq/u9HSmRIxOOA6RWxS/YMLjERK+eXEToISQK0t1QcdYa
8IIETGUvmB8NaLFXTA0+NZpFtirCdKuG+kyC8PczNd9wzLB/DFjthHUhnyjOiH93em3mAQYZrcFO
5/ol9jj8Cb0e3zB6+xAvOufBqX5yzGVuH7WGlcYqXLFTC3LYnR8nc0TpXLPp2EWxo9Xrjq4ZBCIl
HtTmfmkrLV/BFHZbFawV80CDX4PfVRVad3akzgVJKF1BicNpXtsYb9Vp2zp6ILk8Kzq6bAZSgdt8
QFxUiEBSgmbd+ulhLze9Y3AamK/vISD7xrxCUf4gGAhfJcMQ0eRweC9W5ej1TDOzOjxoFaVdj97r
YY4BAcBYXH+q+iA32bO5MY4QZbJgE48IuGyWr1m54u4VPFiFYbYHfrngtHYWyzv7udETHYCwLcyb
Ee3O20+QfHcseg5aOKeligw577UPUGXFjopI8X1uaO/sU0R7Pg+hhto4RMc0UBfesEai2LUkoaCB
EWI6nYxuc48pyBNKEYRkwolBMT5WlB1I+0gL84QeDkhRLlXyjVydlGdnX23SlCTjwbu3U3iuccoA
tfE3aZZsHIhxs5FzKdV2yoq3jVwNb1ZKxEyLLILd5HcX4wvmQH0IrbAxtiNkaPJMzwpFBb9DxHQ7
2c3VsaybpO2fbMDjdr3kUGsGJ5P/VPcpZtsErtxD00AfS055QHmac0aftELQjXRphDRWMZqzn2C9
jkmLGmhckh9et/MjPXSTuj4qajzUHdSR2pJjj461ErCEppWRBkVwJuciD1aQUjU9f3afqdSfhNzh
vPL01Ea3gfUPjOk9OwbrpDTU4Emo8Q1Btx8xdUYgqLo1XbU0frEXTLHXf/yUOxI5qnqxfxop2N6u
yXT72V28ucMAYxXmmUhEJkRiJPd+DzuPY0n/kwE+hAmWeUTvE0iGJJDc48CKWSU9ofwAU+K2XzKa
MZjMft8QKuO6R8AcONTzl1vU+SxGLV8Pif9hcx8zoYsiJFHxWts9Xwdm68kAKASV4aUj97Wlp76p
mDiu1gNdI7IcxYWWnIljSEqisJxh/spj9bJg7mYVzzMT43UdAW8euydJTauv0QvOGse2D730sqGm
fB8dEmVru5Sb56ozviJo9UASih7LEyn66U4l9U78XTrreUEzTW5BiuwI+/Pzq8lwmiYeVvQrFS9O
j2LjpAZM01vtm3ZQ8ewO9SqeTnLjACMbkVqSZknZ5uNn5woaKSSaEE1JZOjiK1jjNLDlUv8jxrZY
0us2x0ciPHe1e1rTh28UANo6CbbD5K9RleVNUpEh8L13QVnGgvazHfqQH+vlkFSG9Jsh4wmTS5cm
a1DigpfKGYPPm65bb6rZ8jocg94rkx7q9dlNaGmuTfI4/opLGHfjg9DeiOrkieqJfxpsZTIGMJLf
lwJFAYpQpvnQbdLv0RVifnUoj0SNX1/m01F/HutQ9WqWh+CK7yCBSMUhlzxe2R4WxcBdeKf+U/bp
mNbpUH0yjeVcEPCHNsw3ZgTZmhij4RjxvIFKNISk64upf4hUs4IYOde74yXDjUph6MtfaArOVhBH
hqP5J3yeSjqCIW8KW0NdkKNkihFzjEu6NY+6HO84g1H3a/KOSBa3jXyVOhksS1AOtDFNYsqQtA1d
rMQbV7HUN9T7l/d/y+IkIKjGIHNs38eWB+JhKfz7ERwEaa1kyeI5OWYaud2yRLUaz7gLJeS8zJFj
SwSMq+OO2WZ1FzOm0DkJ7tz7ohwEb5yGD9Bivrdu1+2+7/oxw8tdnonuGRDzDNAfIhU8E0Iu9Ojy
PDEVTl/m3pOw8l2zxYAgPO/iC3ZhCCTHa8/nsFDiCGNavHkg6P2DCKnhIXZW45+UJVyK4Mml1TFR
pPzffV0i09uMEu0ks7E4QbbfbcH2TMqSnKY+IdXbkJIZ1QNtytAN0UwkTy7eYpQAbSH5SFHxzp7r
1smIwCzl6uXpIm+qoWdxTwHO6EpQedQaOS07nhzKjnUr1IJRtBxqFv52wH+IajC0eUyEmw8Jjmf+
dWYs262bhbMhEZNfoE9eNhYyHzts7wqc7gZv5CnG7RXBloxavay+P3g4eRYkZciu1PbMN9BrO216
Zv2cznSq42fgvNJNe6mDZxvSji960+sNXIv+L4IC/d2bzHdMLtT+RU9SzdCg7mNilC9+/uxU8vjl
cv+jl5ddsK667/XT6l0yvM4FqKns8U6cwtN2+0KAqDpZ4Nwj+/o7XWQJdddPbg87YOJy4IGiDQRE
CIA//H0DnDE9BMatpjeWtdadRY79k+9EHAlG0rHGf3XGKt4HCDt/PcTBrEZGtmnj8cz6kcOTf8ql
HUKqDYzuUovVnV01biNkRr16h7q239reyXZQnEwJwMu+RdtvlhIeunZLgvtj+bU0aMHTP7WmybWV
HCJB/BLQJWhrHdSUI9h8b4pJA3hd7lygOZHRq5No8N26SYteasPRHZ9J/XLY3JcaDMGIdkE9Vx4H
pHWiQrulNR3yBPLEkr4uz+cEEG/SE9OaadD/KgVE5QGXF03oOHMSz1Fq8QI3AmOGkkjFLE1GjQ1k
rv81CDwyq9upn+Bnkf8zWU0dH6Rv8s3f8OwVpLHJS6lYwQudpUMYWW23HyogkvluYuYS8tKXR3F/
aOUwApD2Ok3dPShsJUbsi0N0fPiX1VHOxqRaeHLBLXvNoTx941xOoYM6WmRs3LI6rmkziAr5C2j3
eroam2DuoSwfhJsEoogDLAHPqVektLW95/bZnPIabNarVGar6/unZphTHjN5/33CpmgWezeqb9zF
uLHsfLDG3uLZgNth/d+SnqiymVSGegf+z0O+gI8KRRbdNqvsBPVBs97R2NbIoRmvqSBs884D6GeA
pEkKGWu2sL/PEvvmAV1zUz+UDObUfz2HUnKHujOCsOzMCJXpYjQ3wOC7BndtvFENWhoyvk2AgQ77
LoAjMp/6axHdGquzxAay0bv4RYOkfoxP3Ud0x1KxEUm0r9oPO138Quo2memZfRp3c/68ly214+9Z
uhtYQK+HnrSE8dZgKTCbXaMINh7ZleDSO50XVG9aZKW2CthpfIsGlp6gKr5zHv5a/+6sQ2+CRwoA
c96P25o/BkWvhSal+Y/kXsZAUlVgqxH5z/1+t48iMfd/F5a+hg79mRBsoxxvTi6//LueuH0ihoc5
+L2ZWTSb/AArz6nH9N6bTBTxnsw+3NI/YiDx+M4qnjn2NU+6bVbcGYE6v+QpaD04L+yZU+lfPFB+
wjOQNyNF59SOUbOakRB82lwQl6PUOdv5SjehjA+P2cJCIQmwRPUgSjXuXSquX9rAw/t+3xqimkJV
6RkdxsWto7ZcDzEeDwLSHU+FvLHN4z19f74BrQzvqe7j0LArVGMPWDoIf+1zc+6DomHzYAiaM58R
vNvREmt/GNZdUAuSFpmVv7ZFORHpiIjh0RjcDQDbOqnPwW7Wo0y2HgTmcHVBt2Piq/+rfvMbQkLs
6qBaUTJNjdD1rEYBHcC90wsq7p4QMScJCGy+G8llXBocEdpI3EpAwoopRmdSkLN1OHqHhGgDy8RE
fEgeRMLNcOdTesZLRhaMzOsDqjeBrMwI9k6rAWa0xo8EW8lWldA9TXUx9KLQpCi9GIznijn7DKhe
Co+UluP8nLZjq97KGlxkHWiotHZBn4IaRcCu+oMx37ZeVFiFKPSIAw4bBp3YxB2Ubl3agUUJbURX
xHyRUjTvMwaa6mnLhlMn2/uUjS5TyqspKUNNG4z7+OP92zRnfNyumoD3JkckjWFjO1gM/mCmKVBM
1jvSHfTIPJtY/rUEX8Serl/1eEz8Nd2o0ShQvVpxXuZJV2p9gFTzYNSkOCYX9yd1dnf+g3ZFLNKX
d4t9beUr/ZEnkCS+uaFwLionEZyJhZKFvAtyrM6qM1afm8vAuKBlicW4OPr6zt+gDHyhxAqb82KQ
zKN9CNr9leNIa2/kh+aNbXnUTB+TebV3OJcNy2prUe/QAuGO0zxt22bLywcrQXshmFlx8B0vpF1r
3gUvXbkRLXMLvRNliFHOBBPG9ZGamPIit5y8LsZIbOOWVUSnxTHYKYo6/MN0mpjYGmAbIPbrtZQV
k2Jz8lLOG1w6VaO0QPjOt3HaGfyLEDbCXe1o+krlHYak4tc4sznCElZEywZ4R/3N4lJYa+dRjw1e
PXG93bZOPUuzfHP7gi1lH/GcCLzTQ+PqDFLS9rOgN7rUxCOVM2tNnBoMLKRaRJVOhThskJCX3P4Y
/7IIwZDGhpBnWs5r/E0aEk8AColgN+xoZwCLoa2qCzXRs01O5643xLLSn0ZLlXW/ZIbgJwZUcKsJ
EBP2xix9n81kZJrMxpreKWgL4z1mNcfsxszSmF5NJezHMWWAs2OkXH1UJt3Q2aUBWIvYFwCwenig
i5Nd2SMZeXZQAkHmXkadACMbPYYlvc/xwLpZKMJ5ZZy5QqiOM6q6bdGBSOeAN/WhUwk7/Z8ESVRW
ItjXP3ChZgEF4FoibA85Z+64ujWOsWLrmTPFHwBk0Hncf+Csv9/Kek2pqqOtGuHu9aMd+6lRhTuo
YuS348PLR5k1N1uSE37W/UyqcoSNslJvDRRrqoQ+GCAhzKDnmdaXu+/74SPtDzSZaBYIZAiRhk5V
umtG9adBqSTFqYGnwJTf6qdd5u+FVYB/gguTNX4xZzbnjJY8Tn4II7+3I4AbPsHW5ADFP0ZQGf+D
5ex4AIy4XXpTXjP6SofoaXzuWH8HZQKz0r5SgAm2f4D4L+MX1umgih1t3v10DB1lxeh5SfNo/lPk
LmmgOnjUdbJhRtE+uetYXWRdS72Z3edcd2FKBBrJaxMcYaByyoja5gETifAgZsL+ABvLaj89cVO+
w5vMtOceIRmFUa1Loh0fOkw77H2h9aVYF8LwG57VIvNBTu5lIJ6evLa8dUpJMfqKwSaaAFdPUCSl
CiJYb8fglI4MFjiZad9rjBITTGSBUFD+ImYW99IcyyK1gIwXy5TSPDQYeLX8XeGmIefV9nbtSa1M
rpeJOocLhzv2fNKuf5HWuMQrCa60Xu+y2C2yY1Ely5kI+6tUcBFzMFb9lpQtvxUqxrvga0AzkxrQ
Z6zX7gO6KSGhKMO+S6B6FWbOdzPCNhfigH0U/4IzAYHp48DguJu4Br7VIEmdXYiHd5nrbhM7i0qs
OpV2M9a7QJlUW9XibNtFp7J4jZzJGj79GUcKC0TayvKBKu2mQ3UgirxJVCNCY3VXEHeyM6m4XKa4
383OjWcI7+bh5yoCG+C50hefdXPNfScDy9gC5f/nSX9g9k6Kx5U2Pfen14yrSyAGu5KQLNgq3m+8
xOPFSxJVn/MxHIdpE8YgE33AN1qukRen2rJdD05R95dBua35qIOE8CAuM3xkr2+Ajv6UzvFq91p5
y2PQNccw21jaDb9E7HAZRowDxObgzUvrZmfOMNHUgjBzHU/6COVyLxF3z/8ux5xGJI/HWNdfs6Hr
eFzo4bFLe6SaInuhyyPLFGFmHkoshYYhyKbHURRRp6YoeC1jmZvkRKxhiKyi/86RdcvcU1GfiGyk
UBEOcrt+B6U2IrbyM35GbTLGpz8lyluZ4ev5BxBrDzwI0So9HzU9fYg59FjjRo6grQ3SfiAa/pXi
8O0kl5I7o92vqPX6b76UqgMdf4lDXZEbL8NoM5hOdsJpEYZS0unAkQfyGtkcDaQ813rQz69ptI2N
saUmYxpG7ilj4S7FpRC+2eS+gyX9xk4VxNLivIcsXFwcm9CUT7BskoMa+kehYf0x4Wnb9/SJkVlB
nd0GTEd0ZoaYDLOeX4vftU0JpCMwYn8udBJzDEXdXa4gdPxmhxXS24yAelBE4QU9T3S/SCkj0NRw
/wVf1gK10JekIFpG5e68iq9LKKglj9UAV+qrsGVz1jwvWL49TkPA92IPinA0NHOChQbiJEm9BRxZ
3lfFn7OlrHspCNdVGwShpxlyZLOr8LvQmS0QPmotcK/x7dguTCLIb0d3ViK2mXabPBF17qx0ksb5
kkMgB6V8a4Voax53/LvVGGV6ZFU+8SvpKpXzsDl/A6KstpZCmk3eibTNZchrpkh2BkW+xGlqxNMS
vJ3AKHqUS57r+PkrZAmV/iR3W48fMl4RCVKOLyDPeEal9u5tl+J1ytg66Am8FVI6IvLZNth5kBCl
DhSNaDS5WXSskLvwQtIlCUw4FJDiHYER9Dlj/KzqaX9sKY9kW2iC/LOYUrjguu8+Fdo4LgSQxl+h
gPwm6nev5vh+I1HPXzObAYxZOhRBsY5nXB78EcgGZmxgpP3ygemNGgGvtsWSD+1FZhlLFDD3mwFc
6THIWYMkbxg6hkYOIc+ggcZt9bhwlDQl0omblFoM4m3ZfNCtSsmehhiep4DsInu8jRMxhajUpUKH
/l1RHaqIZqHrW/VCG26nDKSL/D2wGHpDDU50VhVO66n6aooxlVeyLeEy6gVOWjCl0Q1btGBWGXx1
Es+MYoV8gMedOqacZaCe++SiuKs4xNlRjnC1H4Bdy+Zq+HuYARayQDACNQBElgznjtV91ZyLgCl+
y+jA2Ph7T9EJ27TtLTbd51bPintiiAivNyCCJ6L68me73hjSpE8QMqv9t4QvMQ8cG4Llk9HIVCcK
rJiuYgxUX4reYVfU1rRlqi4Qd2A/z1xFEN5gDxtAiQhlB20L8OQ6VCVLguGthYAMDD8Fe24WsabI
5FJVCsy39Zy82OlYoarXudhxHMnABRY42Fl58QE2MuhOucv5qkfOcDz8MhgX8QXvgoQA3Ze0X8da
dQLQQ2/HrUEgp1lXqPkvblqbWvFKB3r+jcBaDIy3PabaufR4LfgwEZPTuvIkjqdCxOuQE02wMLPa
2OXOdej9MBsgcrCcGhO8umQMHRqQlPo9RlatZKoMv/bCGF01Bi8xHS7F8kJ/fUmMcy6RFi4cJz/H
9AOP4I+pR38c6Ok5pDo6EnWlYcIJaUUEm/GwybWoVn+yGF4l7p9hOvt9Z/MiFAjybBaSMFIM3B0k
c9cuYwicUx9Se/ods9ZdkG6GOq7fLimeaFTJ4snJZE+tBRcjMv2rOCxpm3DnrB5FU9eteBLu2KCz
oWLD/xoV7eKp9G7458fSr4AO9YNs287Yvy1jEHB0sPMp1EfdPqPkgAbr5jGwQLnT81lj78rq3OGe
kFrlw12/Nb51lcRnaM8RBNry+BfIrlcrhcP9SncuY/RH2dq1oK6vM5bk8ILPFk7fHZMionQ6Veut
DRbkcVB9qZ00/wM4zBb8mm99J+Y2hjOcXKjB9k2DFbHlu2xxstknXQfWY7htoMiq5CB51AIMYCai
Biua7wCN6VnDE/vl4IEmV3PpUG4F63jzTcA0NrDpSasLzWAxY+2aL+MAghZy+/ZYIfUEopxegDyu
aQn3RE5YxNfLE5hl4RQIPkxVDPTB6GXHXA/6MMCOkvIh3uWteHPyaeP9orEd3K+9rnrpKzDpF0ON
KmDYuGDOvkGdCsS385XJ7HPGUkQtc/pvXaWjz5DYG7Crb9l+BMbCmKOmeVxjg7S/NgYoq6unCtlG
ctBswo/zlXzWv7WeNOjBgxkPXVbJPizICKb/cvsMuReTAhziJ7I+4rGKb0D4LkjOv+vOiSAOQ2RF
zsIDLn/vkgPnHkNRknh5/LVoW2OQEKMaUUdBoNfyHVT4qQCaJls9o2YgBhi+XrH9hxyNJqUkx9nT
OMzJu0/lB4rSyddf6VrbSM4/LYR4kin3e2kFcyJU0M/kqMSOVbOEpT+mP6FRXXQ/tiMhYvEpAPZ3
CvOfTaXOC1O+csRc8jo9ZBdhzaFzXwuHPk9XOpzizMpBZEB6l4/+Fc1o3rqZ8tovT9hLFJMVNpSy
iVutE3mFpdhalrDZhUN5hyneValbqXMsxuf+9wPDXKsJj7XIFCU9F9GPGzylqNbeI7lRG9hQNSsE
2Uj1D8KUirE1uXypurJS5kQNjzEaUqgUf84RkJaGMSGsZtI1GZbxPlerc8U3Du/2MItmcSVfnjyn
iMaTXh2UnMMh7ih7sxW5k3y3VmB07tf7FPARkuB//gcR58OKXIn6nITOa20SSfkiTLEuMuCkza7h
4gXPVlVYfYfSM3YWgKG8LhKtQ0azhahru/YnxYRb5h7sByTGQU/iwMU7MeE3Dh+NCE3hOgww5toN
TmMucCxTQHPEzg45heTdzjWJhcUznEIJrtPLl+ZIvCpuOw1iH035Ex12t4azBk6K2QDZaVNHQumh
fvCKydprm+PJKMQXvgMLZaiLUXsNe8x6hnpjGBY4L2JIB3aPyXZl6cmClPHdxUZsfzm7mUD5YCPB
rBvriy8qi+CAj0w5PWsl1Cc4KYrfMhqhfAdyWVWOx9O/tkR34P1MRe3m9l4WmkeXwVxur0oP75EX
N8tKPBcUhFx9NCDth8ORR04y4ITV+k9qnCsKr4AN8YmKE8DC/0o+UI8s7sHE41eLt33DDFjL9TvN
cyG0tT28/ozA4JPceUpFfNyGmFSU169cacFRprwjnMIwwWiyrxDk0nllFfLx7E6F6M1PT4F8meEU
MJabUEIxP7PhQLf5E7O2JqxM/9YRC9zKgHA4hc6ZPs7iug4c9b2Ak5EpxAytWokVwy5hIf0I6oDw
kUqSdoUjXrutnH8r6x7luqbW0/mdQgPF5Sr50oOypgCnJaMdcsTtsowp/ofvBsndJiYrlhr9OChM
5N/7yaY0sm1pp2+gsbAut7LvfI9lInvIxgJFMSzXd+lbYa8B7SJo1ukTVTTbXZWKX4JMKhvtG1dI
4qOqTIk7oIAQJfG9C+vhvJR+5CeQva9BI5jh2pc9Z2+GgW2AE3S0zcC0KUu7q0mpmvmVF717+JPc
4V5I21m+xgKglJFoaOaPK67pjJRF4w2WgT4Uha327IgpcSRamJRGLh/YhOiVX4LTjxuz0GeIVars
twvlSkh8QaOMwy0UFg2WsLSl+ANc4HMm+9BFLnSk/1oimP1s85VEzEY/9o39742iumjcniaNECNF
nRZci+RJeMJCl44mkexOQsvcHjIe/Q3BTOrM14/wRpe9HvIpSC9XAumc1DEYWLq5+HTvT9VGRb6h
yASXHbwMFAoQMdoFr7ZSR8n6JOK9qZDo98dR1uT1b120npU81nJkcHa/Tz+1My70ex0C47OSLxx6
zV762p2lcwOJgyvEkSyh3s3m2pHwf+mfuBIkRjquh5vvKZDZSPhxeQFPLkm1DYHRnBHiXd4L9MmM
V+C5tbZSQcWUGSOScqzmmBoTXEUHAtb4FM5bt8t3RgRPzrBHbXgrXP5x91GQ53sxaTYl8R6vfOw7
YaCT9s7fh7bq9vEMuf5DkX1SQOqJGF+cL58VVnSfac0Oac2DigrpLeurzmzvLr0/20jGYjNvHley
zholzFBzMWViDOD782XZoAOU2IV3o+SDgiC7R3Cg+Dg0VYT/Bc4VSeBdoGryPaF4f9aC2kg2fU6H
KJragLe0CkTFhqWLRa2cFZmtaoLBsCd9Z9lUHsKyln9jGxG9bAWwihQezzftwgY4JskFFpoHueDM
FFwL19bdtL2jMICzAcPEeu5UOi3+kZKgbM3oOn7WxpMfCzLbUK2lALpw2ZkuZKjzWDIvluJIbebb
0zXRgNKFXHOkjWY49F6N1bVIT8zCjcKSP0o1ajbF29U3mu6j1u1zkLAD/7YK8XAhNHXj6bd7V83h
7Lcd0drbLx+kuPWVNOKlroe+CEiLe9Mv6UFy+GmVIeMqaFh1rPMOEJn5g04cJd8zqS357Gced6nR
ikGT7pdeHSKepLP/rSp3mFHs+pJOyCjMjxsaGD/zgOT3LttVFyczr22mJT9tivpduFzzGXjHUoNk
wTMNjQ2R3WaVM5CLDyXOQus7XKyTnXdY6vPrV+ZVL++cftCdl7JDf8uqXNat8bN7NxyFLjNt3YlZ
mnXo2YX0MT3lQso9J4SLFAujC9fncT6Vm2015MendfoU/3t/S4OE39QF5r8dShmc7pyjGKdkYw/i
JndLBhIAMjvdUpBURkp1m2I8IvSh0M8qK4SXIsCg3MrB55i7lg9tuoUKV8mMbRvvUs72QlJdmjor
NXJpxYVQl2ziqe8MttzBXUYPMYeaPhPovXKa9PHYclEjnIoV53Sg7pmizWzhCHZR+YtUhM11GtWi
ps1zSnd64oaJirlIVZMfnPISAeuArP5XOn1zS7VMtgCAE/ELd6ekOHX9lEgqRU2GocqDrrykH81e
8Mwazt44REtPLZxl4O7/ibbfbXAsX/uWz5zFUqlYzQRGuq9erk4FF9fO8VOwXiborzy9dyOz+VVA
THNMYus/Ax53OjpYxvUT2YQITmpvcMGdCaAXn7tg9GglumeYd+CcZR9gKeMTpf9/O7WP1TH6fc94
3eoEqOlplBhFNugA1t/FYrHWXOrUw/d49p0DFHaLqy9mTKTvr/FtmcKNZU+O6EC9XZfWQtJgCuju
HGcK5eEiZH3tVGiEbS6mcK35UxxwDtnvuHrjqgRluCRWdGY6du2A+5LJoywiZqw59Lffk8I/nOtX
pSI2BTyOB2o9x3MtbzjkKsdkIdi1KBjlgvdvYJq0Mdm0vaBivd+1E/u/KQFQzhs9v+7ydfyukWPo
4UBReF4HcSy50XxX7TpHjYFAoa47Twm607Kw9rIrLGeJrfgfqng/fwpKJZwNxh8L/vEGzjCutSEN
c0rGMDhEJGnPKltQk3SkOkay57JHzqr5NCx0PLeDm9RJde/uatQGNpBdppC1ojDHcBXgI+EfAHTB
9zbuRZTOMxlHhdSUrctMVRHeYZwOylKd16RhZes3ln/m7T9yRl305qNgz+c60AG9+KF0RCo7Fqv6
O5zQ9yn4mfEhRjpwjUuHDvwrRFU3WQsMPWbnXN1pSSSKRdLLT4gLa96D1WnOXMzvFO3/6Kk0n/06
R9BMoUljcs72+udOCyDEo/1s16rRk4XlHY4tNY1LjyrOYiDpRGGRP+qFhyOR9lgbTSS2HIic40eT
0cYemuIxWRc5lb/7a5v1E7KSAobPSS2UR5e0Moit53/H93qxq9tShrzEHvX1C+tc0gOuWIJMR6rJ
mfQOoSdTC30SAol+u4m1egusfG1rJ5EFzPrAf7LMvo6ZRQn1oymAgbRKaiuUgbapbDjdWxYFY3i8
/0aeC9pB6xKPJKuaKaKZi5G/vS55nxJR5HNK+jKZyG1lE39UgL73mnBw4s/h5Ud7VzRWmmBfyxoC
eurGNTzj2D80P0QI9d2YxdlD/ewfyKdHVpwwt2eKKqC96d2zAcBa3OMu2YaTMy8jE+/H66U8hLuu
YMg1tLd8sBw24fM1wKe0TbtjQyP8dZ5Okkewd0r7ASYpIup1F1CBVb4yn9jx8J1cd3JIl+Lc8Mg2
0q9T5hbmdFg98TIGoHkN9Zn1wRHYNePtFjXx91q582tvIEOQevBl0gvaTx6icPbI/fvyu+5urbMS
4emo1wRkl/c3AbRLsB/vWv4UTcvMnolAS+VmHzAmv59/pUcPSENSp4W46K6gp9hlckcjprdSCpKv
F1Z/1ahYiRWNLjUvUgjT4WBREtd4beWuQOjRnylH/GiBIrEd/ZzB+0zoDn9t60pZobLlqyh5UlW/
HkL7tEYG8xU7xqWxU9Lx/mflz9HIVzkVqiSEmQBdoe0LjBQAcbVf4+QT3u6TnkSy4jd2+Nq4PdGd
6Jhf9eixTF7KKZMZeDBRlxQRVfctNzJqHyoNOoHoSnyYgLjtGzWdDZPGGP0flZRXK9tkPDnUnPYd
/SEcKXErkPLPGcUAjFZAeLRrk3eLfnQsvPgJwbQhi7U6uEGg2AV9DVCyXPHNIp44kE/n0/odMh3k
2QYV+pzscuJsZaF56Pp1uiRdffDHvh5w4FyBRCf4SERZ5jDxrgmBP2/MHxLmVhtmyozLzlTDShEy
ntWWnbFD83EhLaweyNusT+NLJxxh5D1sR7AsJ96qefCAnDPQ//Is4X4GNbkTJ35hpklgDe2YxXRb
1UY3h7TWay5OCMUsSTdsUJ1MjtAaW0fdF4IbR1vMHSNp1VvMvr1Lfjju0UUjJgUpjLQTY+qB9quc
uD+zHiqotZUgnRYwZKwTWQAXvM8IEPPiQ0lILyc0DFfIP2mKnJeuIPRmDD6VCScV476DPkdgYxhn
SVHV08GkUWxyotx4kudHkLvzsy3oNaL0xAutvHUGVROq8tmRh5aF+s+Ml3o/8WNeU6m+9jKqlp9h
cJ8tv2ZqOWFOLsT9aK6wFYkEshEZcL5W0sZmAxYLRQc/HVfZQa5c7MuHAjoI9pHmSfluZ2L+2nUE
mQzrN+wMCQpnq5OAHGy6BTL7MPLQJdDDKvs1dGbJbHdE7TJCiiM9M9n9exdMXpDFh8S0J0hPKtzr
2PUGGhZ+RFpZJUDpiUNGlH6A/Xo5k0y4wjVQ3Mxm5kl0G9+zm4E2SpUzdQJflFRs3zkDoPddbuDT
VAslNxwzSQrWAICiSExwkf1jpKtpTbLrN38AfIOb2EP11Cp7h8NPklv4DhXltOtXUWd4Kb47m9Ec
RbYdb9sEEzyET+QK6aloP105zIBjvNJRITflBA8JH+UGKXrmTKIzTY4HGdHCE0liUFFfvUawRQiC
3XkhR1EhW/5Q+lF/6jenrWteKvxA8gv0ESR08bTFsd0PUCCek6I+HlYJfBpFaUEeG/RChqCVRciP
87erX2EzZOCJaa3AV6FgLFDtRHRyNcMEN0MYJrNaQ/mhjp3z/RldHmOX8S4Xo+R3dICk6ktopGdY
+gewawviNCY3pm8MTGAuwOQ7K0BjGPVr1gtuoCY8MBUzlIF4WNfsFRKk5wXSzebgLHsahpHD75O6
GBMHIXOiNo6ntlmhznDl+Pyt2/Pwgv8lg8fflJEmQgzLjm0hgILls1fl27CDEEl+Ae4f9H//xBfr
m96mFEL6nBIdtRpkEaW1FLuraCYGPU6vTP1St8P3vUrb+oH2QsiFpDdX7UQ+UTKaHKqLKtS7Kv7i
0+2X9zjS0/zg+G/57YEkl8kXWXshHzYmccMWzqqHlyS24C6DfcM2X1w7Sc9eAml58WcNvbwIG56s
4IFxsMGeRgaInVaD5bxveQSpsfF6ZfMJLrwhq0LKAJUBkANio6s4pAdVsm8vOeIAh8c652x3Tam0
gYo4NIFbMo9dyWqtR9TwQkKdwL42ev5zfb8dnXcjQ0j7BCZCAhkti8aFw8ASeYqKP8QCjIKCCqDB
61pK6ev/cBfB7Gi49iFKyeyVntKOIj/NlWUJfbWpIGuC6B8sV63xYmugOC0ZvHyVL2uu2YeXVJwc
vFSgH2NHD5A3phiYFslWFCtOKUeLZ+gzyUWnOcTsbXiHPGa9BVookDvCOmu6KbkAHNhzTKMT0vDE
646AwCpuhk/y2RWaFhCsMLbxJPcWnapFhEqoSAjUCaCvrschIXZzd+/wfGX63f98drtG8HtQmjsU
sdA8pbbhGgMOPNELxQTXqYdiuJeacrzRW2X3V9f7cfAiGcUVu9Bcn8kJ6mD9JtcXfTm/S5eEzKTp
AnAlqrd2CprzLwxfH/BL01E2kL81ag/iOh+netr2PmCOetj7qMSnfvfuSrDbJWX3lZ4udCV2dq4U
y4tEi/MFOaipWygCGZoXPrMsVf31WMfSne1oTqQwcm74LtbLZUpce0i1+xNdmz6atlS3H+QNH7I8
vkBR0s5GpAoDDO6op4P3yCbbT7Leb64T3O8x776XVnNG9tcMV2+B6iBwbLtR/GMCoy/wjAjoQPVc
u4DdGhTjyUs4sCfIFNgELXzdMI9C20fPP/5sK+qCPCUpL6YraHBOHQWGmcBC55GifNj444vKJs8m
RB2jlxJd18Zfzhm0GqUs5TQ3I/5v0IRrapEp6Zo/MUKhaeqFTAi3NF4/jkA3R8mPkIxD+AiUBsAG
fxIhFMl0zpr9cqCAkvKnyACzZeOEK9ye6nufrJKHT6tdPSwlXwpS/iZvrt+ycKQi4J+1IOBryfub
1/oyv3tRpVO0iSsINk1BvFApGGd7s+0Hd60jO8bTU6axRlerNSunpvB92h+fQ4adkXMpypjBt2Bk
p3hZiHXl7/sm0/RqE+MYCwnHjmyZf7Gbcq3Da9n+cYHYSa+Nq2DHPIk/BY4vza/iZOuGV8b2GWpN
M/SP0uu+ak7Fq5VjeCnVUJl49Iu0vfV9VvuVO0snlLln0nsl7WtZEnMD9BcE2W3NjgG1olueBAT1
4SZAWDLzBKeYpuDrLphIPp1oHgW4Vx+PJxZB7mzwIFiTyr+/lNIH2H9Qzv69KSLebb+ORwJIlrKp
kaiNHqsKfMJo0UY1coeGBOfXSshSYhaBJEab2tC0F/grWeffJ7cI5oOMhPseIUqi8b3FSmpUhjMK
KJp7+fSMPaa9qmCn1jBNWtoeUBNYzAHCF2L7G7MojrcjstCzvYHVaBWUPOli+JTxjW9zs5IaFwIU
SQ1YeNYizovF6zLorFBMCVfXUC750PSsdZQJTzPir5E7dc00210pGvkLwa6W4x5ru8uanJX13cqW
bjswokH9qZk3m5F/lzkvI7RPfJ4gRbJaqkup6Dw2d8mGgj+WCzJDTSpsjdvIy23rpEXbNZhdxIwm
OtJHhlH76HiN44xvp3ThndVixaoAhSukgxSdZ1nkyXcf4tsTlILaprb3M8eMN+Fk7H7R1Fg+zavZ
bHGe24DGnrztM+YfkX7i3+g1vshtJXvM0fl6s5YZRAUahHqZB8d/q3gZskloixhVkNaH8eXPlAOA
Neg2I8ZIgLt7LDYUM2aRpErOn4ryR5UMMl0/rPXrPwwhlrxti9WsCNvXSFCMQbj9ITq/aEpWqMnu
xm8TtGaFUakrv5PYFL/uhftymcmeSznlP/hMuDRCkZYQY6l8R1EOJbxdZvNpW0w4banaDRyWPOUA
ArLhHuFZ1Sor67VEOuVxV/XEPYA9TyHg67vbXf81OuXP5Jvc1cvUYnf9u9NSvFwHfS/4UsWNeH81
w5Azb1O5XC9joBgCBwZ0AoqSpcTf55fEqxSIZf+JQyaXVWcmgH0ilZlZGh2aXhmmXS5or4S/RJMT
TUMiVDyCG1Bi8/cq/LuuCQQlXhjkqyeNbdsGPZA6D2dQA2TvQTWfMZsTkQolmKKfgmbo0Z5rCcjB
IeWdsikHWwyX7+gwqWuLKo13Umuc8LNEY0m+vh+h/KoaUKNaQlDVafrdbpHHg6S2c4DeofRJKCFz
azpCvP1jTZq0bvTG07BrM9drEegRQWJ+arQf3GN95IZutuODBI96gV+lhljKoNkx8cKWlOX4vcJK
88oJXl/whxdQ5TgzTlTjrBeWQB4iNzUWW03BFD9X+ALKIwXzTEnOMvmPMFinlDxjwwQ+zscYcHjj
MugbNfbXUFVD45yypsXtGKn/+ilmD8wP7S+lREeV9uB5opLcr5NolavunrsSe5r8yMPTD8Q14r9N
Tj/phsZUNUZBGlM92e2Jr+fNYUtvaP78imuGlcPu5dkLRmapUmFOt6Nc4Jf1ykIkKJu3ZaCaddbE
DBiPhSKE1vzzB8FaNZXhewxwR3JaAoFy4TU+urYfuvdUXtK46Mala1KLCUIz1CywCLsYw8UT6klW
TD55/iTEAi7qTvMA17kVsiQFH1mYwn8rT1ihxH1mETY/AL9hI/dTB3f/Xn6eNfXA+7/MqfpjRGnC
dixJJkaLK89LNP0s8T4CK5d+Iw33MTgKk8wMDjaCsl4/nWtlvTXaw1Ljj1Z8idr27r+ukS+l7Css
8jCFdkkE2uO8Ybl8oeIIuxKqK0553U+/ICNHuerMa5SrlIVJ/EW0fwczJ+yEduiutSHO68WqJB2S
jTyW7N9H5yZ+ToD5yuo1g5boCmUik+6YnXSMHnnDammpbG39zzjpfxbQTjMFTMr348iGf0/RqYFX
BDeR40V2PHtZYndk664uQP2I0sMy9ESUjT16Drp/D0Dz476FjwjRfc+FjqsuJD+5DGmLErU7nLgC
HN/BvlBA1fLfW8zb59tpDDd0uNfDqFtM8XtiCbwWps192LI5ZZGYJmD0XQ4Cf3XKF04BJIwLYGZK
6wIj1ACYjNHDC60DtZVIaEBvF0nYximh4qlm835lE0iEBOertuXPY4F1Ybpv1cU/au2VoRrfaQHJ
QAhvB8zLfv28EspGOq44iQS8Mj38UT91HmlBi7JyKXv27lOrI9dR7S5xMuxUFIw1iVd+npb35AFS
rU0HGgYr4n8Q1uj1MkWszhzhQWnFVJXwowxgXUbzbwl/9vP5xgmNb7yjRwyvh4mEa7kfLPX1AIRq
/KR2kOyb2qBN/y00RE7IJxhZSCH+njEVbMgiA+MYgq1CYAQiSKTsQSqV8/3IwGim9OeQd7u3ZaEX
NonHIQX6Q2zLLScDFy7/c7wd47s6P6JVsMSSqLgsVTCzgWiABTpnfbCYcDe64lqkf4likFEZsDj6
kV8mnJkp6HWC+BfkI1Xqvgd1fXPXpj4FfP2GhhSBPRysU9JAVRlKHL9XImkCcseGWIu3KXOuXfsp
AAbfXHXRCMrKBe2EBB2IZzjiJ9PYqZaNisrkrv8uVoQBO05+6lyRM8iqAyXUAF1hgmib00Mp+33Q
jYOEwYI2XpekMbr56pccd0JZFgyrwUi4D1RtZB/1WjTfH0kKC+Ei6K73yvK7fBehg2Du5i+fs7u8
E57nvGK3AVPNic7SXNNCsFdXmYHiXBS6KL3hGLfGyfYYeAidsPGgRXxd+oV1w7wXPvpA6rOTELcj
jciNSG5L17Wwxwpy4jV3o4+NyGb3SIIeI33IRmyv/1F+m6tjMhMnlpec2wgJLMAj2hFxuzSCMpDc
MGU/SOBVCAbIf29qSvU0esSLNs4ivVOORqMPn3a+CT6EqouDz6HPi5zj3F61haaLJhlHD83QWMX2
KS3RdGJjpr8c9f5guaqjpcmjKFdCzgvhJXME0Ti8jPNHDhLVjcRDdnO+PbZUZbVCfh+fY1eve1N0
aE8xOwb93S4yINuqGL8jhLq8sn7l3oQpheNo3owEW2u8LvcQsKcaf0bUgDLZ08+aUunZZJtY4I/T
la9E0elF+3L1UgDcTFzrjckY9vQAey4zYiP7MQ1t7jsmpVEFFBjNuzky2nIa8EtvrX8hAIHgtvaX
THLwHIcOyLkuVihp+KI2RZS004pt0+LxkswZEAeCZe6cTLKs1/OGKuuFjCxV8pR89GS308owY09n
jknimF3wuaTsGgTL5uTfe1XhFrtQvboWA2vo1b4XeA+bvYtoTGiaPYSMHTqS0vR5iLP8PTFMvgV/
6tYw4x8XmBm0pOvrqVxLw0BDztuQIVTFTqnim0sNi2XKNPk3NX8rqbZTgvZx2FXTG+X71lvLDFw5
XLVc/J5Pi3xFdKwWwPFo8PTFBMRChUeJSKZF8mgbIOPqF/LyyCq/Auz4QAng2L7p2X2yuF/qHUlf
sOUWj9yeO+XWuOrZoxY54xh1r+/iq8oZBlm5NsFNzP2Su5uEsU0/RFcaeuJPk5jy+U2fIxSpfxSl
7QpSrV0g4VdVOEsbq+vsO9/aFaxhKkEDtIBzcggmzVRmMyhVWy4kEm645gLwBOznE8aOUR1Li16v
v2KEugtZ6JBvk+DZaTSVAknShAHA6CLiNXMZANme/SKU9Hb0kUOawzOQyEBDsNCTDFh90tOrjeVX
1h1yf6VfxS3oE3VN2mEUj3CNgYdl9hu+hj8+IKn1V3gmZv1tuC8I6dFqHaULnQNySBtBsesuybv0
f07TY37nYU+42rWFSOBLb8Ewea6G2Ckrvqx7tzFb81VxsUKHdFKZLYHlP+nYytBGa/xIN9FaEoIh
YW3bjnsBwJko6C04FlYtZsDLUiWs2BTG+ZOjrckdKes1Gq3xp9l8pSKueqj5HadUqHAsFKM1owcY
Kjjr+gwVWE//zZ0P08MlIi2Mlb2Lvfdmv/DqGfwe+xAv/U7HPgcYNA1bY3FLevgqp3q7VRh+o1E3
r+nY005OLY0HTfwK8o5HPxGYCaADANy32pUtTuGYY0w8GNKa+o7erTwO2akweDmst7D5PqOOg8AU
0JmhIzhp2MpPSZTJG7LIfkgS+lqDRZvjVZwwa6lKdrJNbUNOlL2/1B8x/2AEwqW0r5R39JIAm+u3
d82wQS9LoB/rKItoVwJ24/HXbD0imieqeWr4dSfk11cJFKS7FKu7Wz4CMT47gvQ8YZzYPQlFnWlx
bVtn+FYHQjnG493YXfycjMzCcgmrnw+RKsURFr5heVxBC7omXmEsr/GOUbhLY5ZD+0vbVlNcUYpF
234Wj9H+7ZnEAN73jA8OI719nEyo0QRr6wu5n5PgoyyBxIs/uwvF5aPJVNEPSSJva//4gqmfetz2
MzfnNfrn+KRQWFzUiNnjuborjjN7k9w1stnKqJWl+SmD/0mo620300WH1QuflY4/jdf7ZLkNe/Gh
8Epe/PVHnP3ye2AJBsVsbIWj2+GoM2j4IK+o7dULHAA1dg0gSs2/cTbqLO+xYmGsbetPFVo2ijSL
64Xgr4hkIKfpPXwH9NtIrZrCO0CRzfUDqsA8Qp+qiOF/MoLxvxNR6YcZ7w+QLkeHwWw2O6pTD8+W
c6Q8aeb5SppyT1fZcUcPys7k83T+Yricn5zMMMwZhwIJof+WesqHAQKgB2DA2Dh+BNulqoOGAG5c
Ee/mlyh2q7gvaFP99jZaXYzms8c1XEWlprlCPUp+CMc4Cgm7nMnxkcUat9uIWu9VCzRLmOvF2lN3
qDM00msox1r90WDJMRFtkMefdORa3ywqA7QXudQQicGhEb7s9sLWl4aKuXLASTs43ytzBFBLLe3w
qc2sm2aMdy7FXuqvoKh/U1SVF7uuw4GfSYNf76r42cW239Hu4PleAjN0nuJWktm9bq+Wlj4U23bu
rv0yGTNjG4M3kGtdTPiuHGHndY489aVXrBHWrTGPaXz22AeuCQmNZ4uCeQYXlz8q6yJzp1dF7SKU
NWAKmWDzu9SasB98MsJlsq7MUbvVRBztxXEI08H1yxX0iGHJH+dxvjpGwFZaJc+zo+PohxF7TT0j
DaiyYvKpNh5FRYTEYj1tpcL+1JH2OGsP3JJGGUCFFfaDqk0lWHVvvRqGxakMJgeKueKO780L//Eu
MFPNxYU99I9JOngzv6Js91PmwomQbP10iSZtLrGpZR1qr2I7n9KophrVKdQ2YpMACTPRXAhKHAGq
ZqmiS3nwsRIUguEL8qAYtLFGA+B/JdnxecW8to1OAQSxcMEocCVsd3kB5suscB8wK74+Sff3anUX
rX2Vz5D/ZiBXbJiFfOXulQdl2PL2+rY0SaW9GAZgBh6b7dfkiw1rNsaAcBhw3DxvlGz+fikmM7oY
xkeR9y1EjIZkTFd79pJCzZEvjZuAQ0krHiZG2RrxmgACiv9XsxTFueGZ2hpcxpoYcMReYO4XTAmD
SqMCetS3rypCvd/U3iz2kaFxHVs18G7vNp0nWEN3BNd48neYyQdmKN98q5BzSPOO/3Fuitsa9EJq
yWd27FYmiGUhCK+IF/wnazPafRxSFooGc3KizqcUUaCx6tzns5LJgVUbHe+E69c4PL0+LGNVQ0Rq
HSKWgfUE22002yGIO1h9I4fYtryIlc40jIg8tYL27s8qy3vzbX3VJwkIVGHnVavnOO9Hr+R/VOo5
82gcTppVLlQ98KCZ8ESfuamFoPe/dsvHUaDJMiMEzBsN5zN5rprUeFR2T4AQ0WDz9y0Y5+gFDEIs
QcTx7Nggj5xIi9nOx+GE1wtmNJaGOS1a9lR3JLPbVHPn2qkLmWhszQ6yCZ3Yt1iLcAdEoDR8fDrp
lwIKvC9RXGn0ndDxSRyPwKRTmpIw0y5UoixJjVwP1Fd75hu4gxhShXa8EA+WDh+e+4v0w4AdMPqL
9Zc94k2u8E+J+AFGJ/VNeGIGb1LYfsmiNk6oZEPHD+BJV646DOD2EoISZrQtw/T6biJFruduQbY2
5/ZZQCHvoREIImlygow1ZRaWjqlwqXlcJgldFR8zcbqPnf5oxfQpDcn3JPxXIES5NcGBfYdEMubx
XHp+Xd48GMrhe+TYSngjRXmxeSWhtuVAptjwcvAkazP4DM0lmdZuI+WAaHWr9mxLAyQ63jtFCR3h
9GDjgTAo1uKOsxS1u2JVC6zpHeBPjPqgvV2o9O+CmJXHpdZHsC6VSVXiXwbq73B6QgfLCSpcmX0d
M1naYQA9vmMo9eIAm5dGMwzDw6awBQfQ6vIiPXUkuhMNSPOrSfu79S14PwJwHnDi3djVu8Fb0JXo
BkJ2nYKYOaIQd6TK3o8LijpcByY4bs9OJKw62FM55BB+hp0iMFFOikehWYub06wV0dsMu3PEEw8K
wmzo8g5OJYYjamkLaBQjd0OXLvNZSRsita5e7yRYBV1syCQp35rcdWa6Ks0d2umVcL9cBBPQT0A4
waDdhcqDnrw9dOhFyNbIFMaYD2oItiqiLrB5qOpAoWBbRcSdVldC7siaaK+QfeTspORigXirMge5
V+inkh+3eQlaYfzDFMsac6VcO+fZkl3aeTyHNgLie41HWqLfslCr0AF3wtMn4WwWmAumK4thpNnp
LTpUPjooqU5V4W3q+GqaH9MBw4lLjm5T04zUBvGEz5rWa7zoMv+lw0qvtVeF5QyIn2cIGC+RdEvW
wFWSYDWVV6Brk0swLY3x+fvNN1LQ2Q+BdR4LwMCYKUk5Cx5ZUJx/off9POhWsKuo877Dgq/Uqm4d
Vw5QZc2tqWFFWjFCrwjEm6l752YN273fDb7Z2eJL6MTTR4gRX9nbqXBaWz1lMnmVqeR8byjbf8c7
0bHY4BPo3ByIqU9Y3iVuosmgnaCp7M5N93h4CsQbVY+HVsaDejpG+oNAL+5KeYRgETECVlLq9MhT
ik9HcMOlzFmi0edFC5aime1rmQXOVGwtXtIXsnCBL5gaUzGocIZBGkl8CaqdVeUaLJpRCu37U0hS
xLJPNEuwsCZDJycuIZJjRq/i00lSmlsXdiCDgHclLOJ7gW3z5tE0/mDnEYA2ELGfCLXv/XzvqcCq
O5bpm7+V2aZR4dNmyGkB9azAH0QQW1+BC8fuFQJtMN4+owMzMuF3+QzuW0sK3j07yzOmun1z71Cp
yejJwNVAl+M3BZshg1zLIztiKXyY85SnzQMRV8+/PrA19YVqcB2a5f2UAkEAzGvP4rqXYRLrfF8r
zUFnDVEco7hfWJUBNLWlrEPSdZhXlISD10j2ShzM54miPoXJ4Qv6ChkUJ0wqiTSZ+n1Uv3nh6fOo
eP0ZsWPSLh12IIAJbw7auT5beo1ogzpF1d2i5QskzKtlOyw/e+kZabJfZs43HoQ6yMOM4nxMOqeA
gl7VIr26JSFGvQunufyGmqq/cOXxr8f6fq8Xgt72BAY0jZycTi9flPqHcqI3OCyeuf9Pvr/V+08q
Lwmc0F6d3cBFOZPjRKKfCMbtwT1nPu+2dF9/tg6SprjVUhFUDFXnMVRi8XQAzUMbuv0us88fFrWA
ZoHIKf2zuEpGzsWuNUdg0G5aFPap1lqjyZBdpZaojgalzrJoc4WdoedcN4qmVHt5b9irBwWVKZiw
VL6Ja/TaOCVVdGfMe352g2nXriEOsGOOD3iXgnf2St4Q0L7RIy0yhf7cPAs9xHtzxKeflI4iDIMF
ZfLLsFU9tMMVsfUeecweR7qEknOCWYa61neTOSuwChHehMZ7q/J42zEKDLwmXMuIhlMgGfNf2zWF
qryrc2mFgL1wK4Z1sl9e3NuuSdVxaO27RZSfXaHQ5qtFU/B5EbFhSIgHkXSCYo4FrDxuh2fMhzf4
QT1pcALn0L0l2wt9aFJ56sc1EV/Hb7Zo2PEtXjxoEQ57oBE9tR/HvBefoPH/HZU0Y/FvFPznfp9X
t4jZltFU2pPL7DBCNq8+5WOKrIWoofRZzxv7fxO1l0+4sWAmqBXkY6RXPzY0dHsSnwWbX8pJ45Tv
BzLidCVC7XWorQAi+utqghLEF9ieuSvlw4EbX59sSxtGOOJkMzuTpN3wv4ODn3wvfkekeqJsKmTf
u7UsDwn5EAtKTZfvPGy3xyMJ+N19LQu4UciNzhiqsOvFismx6jMsipNvqNLJ51b9ieY1xNqAcWXA
o74abTzS1C+fYbj8Y/9ycK8CWmEGOxN2fBAWNEQJBcQtxrIFsIAgqz0Pp3A7o9Cyb7oRqqik1eZj
AD0fdeyU1+AYVuXBjMQuY8nFGmmhxd74+9ikqmKFDtVcye6epO/Pc11dTOOdqL1hA8ReyY4vA9Kc
QS70Bcf7vIUmTgZogB2/Y5jBY0dVcpsMVanulXoZbGGmhkS1Zcvrv0Z8GMgJ1pEOUrfmoPIy6yax
lpmLXRg0X+oBRVNi1uD87+Cafpu9RxBmx9ktALSSHpkFQk3M7+UdHQw20qN1O9FEN9fB0JGxV9Ue
x8lkKwbNywuBxJjfJkQELwCkbp5t2lTRrvK/rRqujFKg6NS3xfIPMRE9NI/HkkF0rHQhW72Mp5k7
hki633a7fjdBvUduHV4DHYiyqjYLdwWTnzQA2o1DGasuxenjDZkQUYQtKssvNEfQWRDAoIG6HQgF
M0Hndlux6tBR6IH+2CgIcjWTwv7JAg4h5/UYuikMy0einu/ttSMrC5S4dIHHbtX+W0ePP8dOybEj
EMZ1+jWvV5ScdrvWtAXYdVvESoLNlWNw3dGI1YzcdRJIaXUW+fyG6ZNl1al7hU2yfd8uWSFOknRj
IBeE5txoasXwQsUYpzZBkYJ3DIpr5/oGnW0JnkLFmUnHruZoZtr6rtyOOMEa1ZcEEiNUzcQSkR3t
JOyu6JaeYHvgh818El9yXTAtwIC1NK+HFZxiYs6iePLPB5rbBUj6XhnHw+Hp6/ru9tXPNZ+JwwUL
MRdbb5/5e4ZqCjk/RuDX1PJH3vrpcfvqjASpoJkAJZ9p7jpBjFGrZp2qWLdlIJ5jajZRgsT4PYoH
e1EYeUE7Gp1gRV1tYUkzpsnoI+SmMsF72PYQY0pIw2Kn8F4EGlTUs7JDGeuyU1rmTXf7V8+0hRpI
MLl3Itr38mSwoX+1+bM3hD21SBU8njSAaLIZVOXx9ohE62gFnG6pyPZ8cW+QKtFVXnRHtatCyHiw
Ye2ZwtoaaPP8psUQglyItkkZ2gpq/1vc7hmf7K2TrUw9Ny9c66Fab1nskt8hMe2F9lfO6Z1SyBut
lY2Mu3orVESnb11W8qbPI43xuJIMk0SMAeyeRrrYV3yXKUD7K7DEzfa5PkSFzyteWobYOfRm5/iK
WDePviIjTc4kOnYGRw1vF//3jZRKG/MgiK1Xo0cLCxuVvCpL6eV49uPDSpTpzOcyLEnpQw6zsGD5
WSwTPhCe1WlPEprt4U4ZOGWdeLd/ikMhUGOFI9MBOQDZH7ZwXj68TgQzZF3ZR6oD6S8m64cHlZGY
v0ju/iGoVFkKZM/Y6RcJtKqw0t9aolWceYmzOOLjHI2H0y8MWJJvps4hvsl7vQyFksvcnVnKQx0I
QLXAAKpmFPMUweBcHIBd2HdJ2N2fpl2tjmZHjwobYcAICzUOr9NfzSevTqIrjeMpybP0XPU8LzMo
NQHQ6pjnzJJm6bxd76kLpeaBxEMyUM+Zh4LP7f5ChUR26TnxvDYD5BsytvO1XiWT699BchLu8mSY
/qJSlw430GdmbktF6O7Bz/995GyeHXuLA84wXf9zBNx6kaRuBIQBlGaM3BW505hD3YiagYj9a+VQ
KHvCgCeSUMpJWaOoTr9fuiA9osUZ92WsNeLo+UG4WaNOKjFJYaFiDdO/gUad+6dpR1PR6CddxpkB
8OVy56dNfVAgABUuYdK/X5kMaQjsHGKP7z37s7fE337OXploULFK4cVzU+jhFUFs6yHk5mYr+MOq
i3fo/O8rDhxcz3jaZC5/mS3h9PzPMN6GzdCC5Y2OP9uWCJFPl7ylv+ejsjSfhZ04U4K3NmnoM1wq
oJg1Igec0+SFWWoIQtu+oGR+Vcun/EbFffzf5AogkJVs7W++DR2S7LMTvTK00oLEprFo75Hs9KJp
yOTUwoeHrRdiCItftuREilOnUbRI+W6kzmg5T21KRrmQS4RDyygnHYoMOdvED5EhJaIaG77CIFjg
clld4R1eJyHpRxtdNz0tAK+oK9m0E84XhMpE12L7QlI89/1tQrzKg6ug1vumZs2yCGKeYaaH7alC
Nhk3tqPNrzYeT2sbeA0O5rpr16dWxWb9qrL9DCMz0Z80yZ8NOnG0A7S64nwQQWAvBr/8DJTWPAPN
bYo/pSYk8LWllrA6rdIxfh0BSMFIHJS+JrifkaaWj9DDdkjBYWTxKtZhuPSAQyM7m4VoEM4ASzZj
eb39ioeR+R71oXZCw3tBwuPHJpNTdTLIZqgFYv7CHkN6LH28IQlrXKyAI91wxZSP8hCmi8Kf9DUo
WByhJnpMXzsjWWbiGHJwe98WQGxG464nJaKMQi12VKVG8Robf+Q8VWFO1wGtBw3386CklKsFxvud
ewtzqRsTC9DaDcn7cSdeaV+4zElC9JRERwAOiOZaKxcnVQ3LHyHIfL5/naI+Je46vwLzFRfUJxW8
qCSw+k1lAYCfWRWvJFzir1dxx4m8Btb+ZOfBeb2c1npzR0HdiC0IzXAwFPmsdf399GZxbgR/vmYz
DLAJJ06Q+XVXlALXtc0vbXzUsEKByPFoGeY7mQMWRzb88gaFHBzZ5XECI5YFkxJXyuktuRXVrbU4
y1LTvLGOXlXJdSzgCFvOijHusplBbjaklDx/IywVoRUkZ+n4LN94rkcjuyPfYgvlaIr0DYr1/bIj
6X5B2yBiyLQD7bQAYfLAmZQYHDfycGulGzTlSbnmFTvbnZQq132htNsggIUljXUMk63R1D9mKFm7
/Gly9d1Xd0OrIY3B0NJ7GM0pZOcEy5AeMqeS7a8SjR62uFS9XqNXno80ilxZRxxYnWAPKm3oh8G4
+WClW3gSoVU3dpqCWxJUs1EfWegBnKkYWA+epssiIPQh1/IMc3N7jNXSudPA21UGbjLK6jzo47yF
yoiO2Oer+Wv16yFWdtRhR7yx5zw9Qatcs5MkoUqu4IQ60TXcSPy+4ULW7bcjdNiW9ijE5gpIKOv4
mLItwjquzAS3LHdL2SGp2Y0d4j0FJOH9pds/VZDyD8Soy+Wy9h0KrQmNWeIuugW3uORqCxWesAzT
9yy29eDhvW2Lsqq1wl2LEy3QBn/virATzzsLdBNibJ6HHsxCA6JUfkDPKoM4AR4JSXqEQYMVCMTI
MI/PhxX8iHXdcBF+9/urK4MLkSciGBRGpYwH792PYrHxIU+SVDwIz6auGcd9DpOtznzKsV2XGhRW
4lwxNwEHXRR3uhH687iJPH6IQEdou8PVyLgE9cUW1zHdiJyGbrWIC+urBs+B+EaRBfwrFOYgz9X2
tjS4C498TrDgAch49C4RzcRuyfSFuEPUApTdeqNDA+fMyyzUoTRWQCt7UkH2rLgD6pFdoz50+2lH
i6xct135f/wSHOAlOZsdpy0eK+75ndREP/MVKHzp6sJ2e7i6TcmGDngcV3w8HTKRMlR2BnjW7r2l
Sg7Y+e0unw7Z3UhIGExb23BbDdVRWjd+sA+gdGhqLrGt9TxrNLAUmPc8TNbgnC6cvnp7dDZtqCPY
5KFs7ghPjYwqgDKiWuFFgPCe5D/hQjPuFXcNooEiNXKvxb2+SCFB5XEudxGk1Eg5MyzeKC5y81ol
xXt0dBK+XUtznyVa9Byfsc+nhNnrWtACSzsinn1Zk+OjeAXGXzylLQVEY0s1XtPwzkiYTbknF3hj
5iN+K4gWTJs8Y3+i9Mun0DHtsCt6xD89wV6sz1qkl9YFKYXrnSOsYgeUrEmoD1PBfct+hj3PSc5+
+6f361KXHfjlUMbaf3j88/2myjx7GKQ9t4a+cfHAw5qwmPjYFRsYeNABU2bWApkzINHLTQG3Yv/T
i/5OZp+XFTaBvTEGsl8CzT85062kJHd37h+0kk87GKk+JoVFZv+zu6FYO5BFN7Q8inKhRX5dbE7a
Zhzujgvos1zEFXck+1CMQB71VTc47nFKHMK5WkqnONLNOJr1xlZg9inB68Ap74yv4qwoaZGYkGBl
59hiLSV6F2Xh1rlW+dLQLXKLopChjOUno2X68CVwrmnL9Ei8d+pglIs/rGXvNxrkSQc11wxGriZs
ijwjqt8c8O89Pj1iFHxCn/0X2/u6ZqsvoktzC89id0uk+vL83nYJWaP3ftHKhhbsm5LD0yCH3Tce
vYQl2OBY/p6MJDLQCsDRodTubA4sSbU8wsTVoypmJEYtmfjuKoCbXpy9dzjb0BG63mV17Pk1US7r
ecVCqXHAJaTIwp1v2n3nvnIF8SrXLCFxr+L+jhSy0fYvjacOtdWoqzCnbsWeOgUk20LcMxUUgpxF
1K1DI1/8lda6fHurpVdWc1nRUnyhuPffeQwEUq/Tk84iySNavj8OdUgpRUeUY8lAJU+3ADZLSYZj
KY4gdLiEgLTuqMmIERifGsnFSQGvdSklCI4uTvRMxVE0PxiNrGa85nHNro/Yr/TmjgtNQoHCteBq
Xlq0M3yvi4zaaAGxfPtMSAuzNsNJpkpAryELkKFBApNm/XkLF00Bgv6PZvk2/1Ndv6RFnog9240K
R82h0ooyubXqrV+heNWAqmck25OKGF/DbsLgwYfoyfKvLi9MXSKb90UiAT+lMC8Acl+41U8btLjU
i5qZG6LELJznxQeIJiE2xLdwUWg+SeCnYTn4JqR/V8a6Tu2qgt2wKYCqfp6JnGyKsLlUdk5IO9lU
4FT9IjA+nZK3MPrYMXkmXoLlP/IJJbvgkEJR9FA0aTNVZssIj+ksKVel+cTQtvuwtmaWjEQYOJut
9sZHc9AIqBDDO25txubTSx75Qwf7AaEx5iTGveCoP7F4VZY4iOqa/Vgbxb5em0IqHbpYtcOf1pzu
BESx66uKOp9fo6QRh2ju2vqSYgl7GB9IL/4LEi47IMJ3X9kYFUQdSwOu2InSENKXwsw8UCgSipuG
6NzdVBPpHJcyBFXA1/ezp2GisivZgyPwy3F0L+fYOt0thg/4wlug5DZ4z374nzksopLbinmWA8OV
KW+XicGXHq7D3OBBkRyBXG4bSY2Qlmrp4VqdU5dTVZHng7/XQ9K1RaZ3rtQ1MSVFTv0G50Ai9ul1
S3J/sjChT4NJT++268URb2yMXJlmd5hltlbbnyLytR4e4L30w07lH5yVhKH7nRa2WgRlcn/bhf/Q
kSw0idBBA+8PYeUAf4ZqRCSlS1eBaOxoHM8Q8Fzm9e6rqcYC0diXT6B2JRGhx2VOH6f9LItygmnG
+EamB8zKep27Apofd2ckPdWaGvx1R7BGLNy8iA/EeMNEoeNKTpRvxCzUOcZbVbfddEazO26WqG4g
206r7PlfcOyU+/s/im97Mtrx/IZWFJgEblRUjSXrltTjOYwEbGZRSNLAO8LBEgt8Ojz25lqUHwWZ
+yhu7Herb/gIM3SbsuqMYBBzp69tD1i5N0Xs36tXREakwZVQm/dQij11VfrUUofr2FE7eSAg5PNa
H/5M0KRvswsIRJxNXMMwFZ+940xHqH1ahcMs9Z6z3HsPQ1w6MBxW6WRnub1dgnCqjNaYWV6IltOi
hsJnT9n79p10p8daBbV0dTyBXGknXxDmWLTxClsdqKcxf5xZZ63Je5NOEuXN2CmYt5Bp2Ea4hpaw
i92+WIOnoGQOQK2p1doRJEtJ/JrFsQuV0HXd4GB8I8Wf+7Zdl5/60xhZAv/hqyrPC/608PMMKpVW
2KlKW7Exb/0W4icsgGD9Wl7t+tG3JkAqZXW4DbNyu6nD+qilFro5E33dG3zpjs8BtB81+KQk2Bsi
AxCf87p6UlbWVr/SXxjmE19ztfw6iVFtnpAhAWQH6tg2voQ2q4i99NEurOhz+6JfyJR5nzROWqAV
vioq6QgIEiNMG84FAPasLLTvISJ63MQh/fcPsS/VAJXSGzQMyZodE7tqXrDjf2LaJLySdV7yqSe0
dXrbqygzHTsz1lLGmEmUBwhAE/8sXu9BYyhBnCF0xMPPvRX11XrWQOILA3rOWNaxbkZtGTgJEqYV
Sr34U/C9YxOHjs8euBreXWheuyqYveaTNf9hCiz7Gvuad6R/luBkc7lSpLn5Qxtv9LhjhFuhQqZZ
+EYnMF7GhMyEvtTIWNR9QCy1qu+CjMdyw1DWhhTh20LDx6znFHUxGEu1ZpjxWubSurlGIO7Bt0EH
BNnHjNMfiKgvOwduRcuRMhp87DGORFL3swfSrlvmAM2YA2xWRlVAaCoCgzdkt1prnGseK09nQuy+
osdx26y4qwMpBaH3yh2Nzf3w4puQEqCnqYDbqWyhrCNuPqYbdaJ24HBjhg/acZJNhj+Nheddk7GW
gEM20JfgwQdYNUCGK+zLtP3ffl8+5xQNx7EhuultENyfkfT5jRzweW+wuJiy3Y+a5Uy5dANqwKEu
WL9U5gw7yld+UanDtihq7sxwNaQMpcOHVncQ6XPAtdiGZhP6gFb5Gs5S7Ob0q3l+qM9UIMxxu2lr
9Sd8q4NPGIY4IGQJhG4Y07V1rJGZUX8I3JsFQLq8Ipe7lStAYLzSPjptsVwBqJXvU0Q60ITUEHVC
Cwb/JnzHr4ct4dJ2eFXcxlhc+m+YahoTn+0nKLfPo9tn1Hi05vPllf1MOZ0rl6EmUSgWIxwyEQFw
LWRcYs7d6CKVuPMtZZ6swNTvKGJDPqsuBHXPb0GhzIDZ8Rk98UZIzqb8L5MPmlEDqieKRl2O6lF6
ivy4/XmL89xd+ESH3y6IwI6q11qVkkG4FlRaUB4s5eGMkmdlBRv3e4FlNNTOZmeJ+FruoPwC1uLg
jmueLHhFoXxt8uShvSQoLGveESXHr6k6x4az+LdVVg+25wYW5RZEfchBS1YQnn/gea7iJgXhlGys
+VavDUk3/XyE63S1hhSXKW5D/vTmwGzud75xg7n7ElJT8eTrxDX8p/tE0l3hNaom+TzNI36KW1vi
E45/0pqgZA4Qlop36jnLYNNj9OWnT4viZ9UY2R2NZqaLIXFMWtaXQtOMp4cha5VhBGw+E/WZt1PG
WjR4iL8kCtoHPZ7uSQPpFKyPWJRa2zyqCBci8nKk55d7FrJAH7D+IZmWFSBfdIh5n9lSGVguzUHi
XHovw13cVlQvP+35L41iGDuEKjwVCLTjDogLiCLroMZP1FIzjIwU9nFaPBXOwFxcJnciIDozbBtd
D/WU2qQashQn21zGdahn8QEeHNdbk42RtAUdY6YO2VfIh5YTk52T7JhhzhDob+CJaBKaeOneTuFW
KxhcBNPHMKzi4P5lZQWcIzpZQ7N35BlHzRsaKIKWxC/14WEZuBSfqTI5X09WM/uSCc0Feg9mJ83S
Lw574+LMkrWd3kX+2c4SMLoFPihmLdu+PXcGqgr2PPFSYCwPw7mmJ8AIf4cbnIqZFbKq4kVH+GKm
tHE5Qr6CU32vDoT2i0aCt3oA7Nl9/4H1IiXOqHeoU/+n6aFf4UEdR6XJJtX6/KnTq2uZCPCuvsor
sAb1A0DRSA5uaXpeFy61fqvV3id9szk0HRDHMxRMPZ7mkEtsFGeotKmXty8QQiBUAA0Bqydm2zmy
1EEXoGG2fhFuNrYO33sMYk9Hq3Z4/lJIgQ4jakLjXvTFvHKVoL19FXf1CRVIA1TkZFEIcYi8fESb
GVL4rYHJZK8jYjrGR7zEVmhqZXHU5bLGZTNQTcLUYUXblWoq0H2sd5mgtpBsmUaEaP3maqmDmOnc
9BrukcF33bANWphH8L2dw/MRsQxhC3MWNuXnz5HG/1eKRNlV5PGoObuB7b3/fvMKdz4xdR8Wr7bw
yGw0GYapPXmrn4XutixW3hXcGbcLEDU/1pjT8u2O1pk0ZwuYWP+cn3ZRd4Z2RfYPtwLGb3Q+blcd
ZFe9231yZgdOyNd/D0TjFZo12LuKKt8TRihEMW1uuXs0KKn4c0YUM/m150TyIU9Jf7GI+Q1QP9fu
vg+R/RPjzcVBl3dYr1cTRFVKjVuTq/zoWckKFoJUdIvJxJ851+yc1ytDP/TXAfWGDLscyW+Hlo1b
4a1g1XASNmD9ZtEc9B7ba69aJOCPDawF+XrBkx+vUiBnL1/mRZ23NSjb+0Sr9iWFlbf9YPvfmP0h
3AnFmGIS1adnukwxvzIJmEYAdbyVo/STVsOBe/FyXbHIxg0uxXovKTVSwtc0t2DjnsgAoys47tZ2
pwDSqkXPXmAq4JeesJlbufxHj/PrUI8LAGYet+FivMCcaPZmKKQOvjSyKbGC/VVltFIaPp9WJtJA
d7S028ZR2EBl7HiY/+9r2tvkHkLT0e4VgWSVM2ApE4ia6YsKsq7UJOXc4jinJIqaAJoPOgJ24SAH
UIkJai8DGr37YQfnUXkg+zsqwCgjTmPhOzn6+ppOdfCIbA/uYa5ZRNboz0PZSdi3UTaRglve69sP
MwaMvcVpu0eVu24mp4Bm/vbEXOOQ/LLd7b8ewiPq+LKRnnl0FYgwscoepqgvg8ATJ+xmqbqfgecM
A/OcNMk2tPDI5dfYA2oQEjckkMlphNvzdRXi6wvKSHq038YPsJPqO3Uoke7xZEYUbgDXPp2yI/gm
e5nY2BOejMFXwvctNED2gc3amLxL15VenjyvcA6sQ1qMQHESI/J7n2+SE+QrqF08JZ58DgAi8az7
Y8oVJwwfqMiLc/WbMW+/6wguU8CLXUWZmksoJpv9ITY0U9WfRx8x9pv+lmYbFnsw6Cp2o14EK43S
SelbvZhy+qzeji78EM90jxDVC1WUQLFVie1s3LM+egmBSfrgP1ybdAq6v37vM0C6gkTVY+rkqWZQ
c+w5aDgsiVZ8bQoGBI47Iic91LajXzybQAUIAHGmr0cnyM4PdWbw3Lhuff+NW11lG6n9KwBAEllP
7YconQnEm1cQAOjRQiHdilJOUb9qk1ewmBYlY1sqTdAfq+79QxZnkZam+Hnmpn1sOD/2G9sUgwAK
rwBIe84iysK85BSOCYtt9N9Z9+0VTC2IAxYVRXt8P5U65QeaoCLGj7sCdyaoPXO/jRTT8Sy2Sxhx
0Mu764zZd1QJTW2GiIVAOQiNQsWMZBKJZWRZD24RvKoyFZCbVQy49TZazHeznnn0EuCH/tQ9fu9w
9m2GYbDBwkmaEnw4U4w/fHKGsEPFu4luGWdJLjxWOiyvLqnJ+8Kl/VseSFWcGBgDJcpE+NZ/4imK
w0WzTFEGC1oEAWvE50TeS+Y6qA3ftxQiOpARaQlArMEg+1TLpSFTfeLo+g3eRWBfT9vMfYp+OuHx
iD9+GMDBvVgs0Rn57w6vbcNGPKRG1aODo2IswUHZPbkckvYzp4eLH2UohhUYzXsTG/g7g3IDX6Bk
EKvA2goTOp0NU9xhoufTCm29X+P0iD4tWS/J//Oh3hGJ2cQBZWsTIEuuuA7flC/K9WldvA5aq3JG
n1pDcb6i5VRAX3p9+VzQdA6nwfz0j4y2fR7cP5LF1Uu2ACAWpjV8O2k9MgA9gCbHbgxu0xTCx62c
RjMt25Yvt6J9W4dCzjpGXB7Oegkv3qFObclNjdOjM91+/MDb0OQPHvRmUPgipUYLr1L6/Q5DR9e9
DewRswB3e4hPmUa7hTgJ3YsnkxZ2Bb47wCg1ipgNSs/hIyyqezUINNTfgYxtgYXeDLc7HZmX/dug
MNXW8RlLeCOwKCpWkxv4ykGI/ypSCyW9IUfXVfSqzamQ6CjMkE7RBj6TFkxKdpC2pXgQ5Bf1zq05
GIJyrPBfKMJVhJnkuReCceXU7JrpZXso/VOP4o4/CjEw1GrTPydqH+OB/AF5rty7EIH4u7OM2bNz
0dAG5IcQm9hH92baRrc47yxj7e5G6AwDA+LOY4823hWHOOkmeam4EXi3/hf93sKcW74CGhWcNTw+
9Byepn/Jk4HKoFkUMMsVjmEYBTBnPY2XFDDu7D7lSpn1cYpEOM9ICdlDTj4sYHsndJwJgIpsx71S
jXobAYFJ9DGp81samQwlOjHGWTIZLRFo7CoLFV4vytJBlBBbsFP1vuuo5ve3mmh3Mk1BHvMQjL0G
8dmB/mlWOwRGFGol4PLW+1xUbo9godvHGFsnB5zg2GB3atQDIJBGVrOTTXPdlBOlDiwXPeFbCVDA
acwTjk0DxcGBuNt8+hn6fXhDOpkiK2Mu9TiePDQhrDMqFARn++7GoFgtHzCQtvmQ+AFlJqQW6oin
+hVeTgcAfipn0PGq4oiXmtYcJAetUv8rTaPk/HOtkImrI1jJKNzYbJrkzw2yqQT+RQkUofh0fXNj
yi6cM25wNghk5GmsyzRU8mbEX2RCJw4MPvqLkaB2FZrszDfA116Ov3U4yThqpXvPzzEJhumMYZ28
/F5NMf6y5H/FKdpPp/0q9M5awgzz1Y+IyHjLHSlGcF9yA9hIS41LhsYzcKCN2MszIicu/Xvn6zC+
NtfvRKttCOBrUNTlvR1OYiOqla0Z2mIee+BU7z7xsjFW7Q5RXEgX8P40PiJIWya8yODCitRJd60C
YIJwWZ+T/FRabBjYfKP+nY/MsftobdSmdl3ZHd66LJLlMKi7hkzmSLG5DzKVG1U6A9GECCaOqhkV
xTJnodIEn7v22/Uah3mnGWM88ePBQIxPH0NE+ljcPL5tV1TLlwp5gTEulJqhYrZiaPTQH/XM9H35
akEwy6NautPpRNDwkoWkCIy7G8juWc4CI0d3abiMEQQvA/DhzAt/DmniM93H/VwWWLrnGF0SqcMs
RBwMGEIbjFz194V36d5DSmOMFulTUp4SpmojSMD5MrjWuHl4YV/Bs8k1i778eO/vN2Qv7hTv6AIJ
RtJ7fC2oaugFe4uvhGGAhQd7Gih1I1mQRgg6ff7oWJdHbj89mkwHq5wVGRuYJH/y2lI/mtuM3rnI
lVDIjgYLQbd5ghhAobqNm6g2CJYhLpEo1iCLvpr8Fozy59FgTqWbz7eIoQvwq7yV7lu4MSaU0j2d
LDJhMNPI5PsDIOcZdVHeGPorBMmpyeMBk+Sz7wMVfIeDa/2jSwccbWvmgCwiNkApHAlKNLkQfbEV
3Ugm2OcL4QykisArBYDouArO9b+ZqKzEUOtYjp2KkWtVhoLT034xdqy2eP6Ch2ue/WMOwpgUak3H
ifdC47TCYdLP8AA0zc4BgXWBgZpvjwyps7EzPWC2ig97Evb9m/JcM/nyh1fwYc/mQT1e5uRKW81D
u6Z/c59X2zlXWiS5Z7qgaE8DBEDN0IKpkaryB7cGL8yOFwTVy7kg+od1qeLdGsLxMkM1rQ6RI59a
RQvlQ0nVgv5YRhRKMeY8fipbZNrlNiLKEcUX1851y7IutT/WV8DwA/J0xiOt1muLLCcbA0xgnxwq
xvcmKixkGWu5cyWWPal+Zfqct6LE7ocOBnwuVaKUu3FmdG7OhlPAAz/De+Rjudcr5obgZjZeYojJ
iUXULc1DKhKHPsJI/b1BAdngSxd/PL/NWFEwe2XmpIGdO0/tpGgrT1idxCGBsmSXAhWmzCrsSkkO
v487C6j5gmxkGvb9cpx+JSVRsAwjUwUVQ7gaeGyaZ0X1n2TBCYZJ7tDjdMiikqY/MLBDn0qnuhoU
L1tgHiNsNzL+T8VJIolDAzrXDkPKJUj9ZE4Kqs/HWY0bH7c6clJWj1mo26Hf+DJbpfAOECrHyn1L
6TEWDTMtA5Ovu35FHGR8SezVqO+foY436icp3eKCxzt2fdzHsGjnFPFOS3Gz8cfIfb+2ew26cdmd
ibZnmZ1L+uky9K8BTtSwXyi9v6SxRwtBLcf6Hxr8cIBGUBgFle9wSpDOi/gpIyaldieYpZbAyKJB
du3o3ynS+rWhGfRHgx7v7Gc3vAoUZEUzrjGQp0RFeIMxiwDtK8GSIjFl2X///ks0AB65X1U75uhA
B6VBB+ytiRcgXUl6FCP/FqDbWY0pUkIMWYHJo7LEN3eWHHFnTcJn9PBHOJAxXW+eCz8aIU8OrUvn
eLG5r/LpjEwedR7ke4qtqfwrfkIBe97Hiyxk4yTQf9wxvOWUaEEH311lEsbp+58Gp6rsXyI2O31x
uQ0XFilJ1LVhr39j4l+x7TBM0kccohy/zqCYrBlTAcW6QKw2ApeUl2FAbOuMBzMr9sfnIWEc54Hu
IGgH8hd8mqiEcJ/0/fR1w3c/0+5eF1w7ocOOo7zJupz1ML0QPANejRayxfRld/73Wp+ZAdbRV+NK
vUv7nN0jUmt1gg2POfSMB2yjndZxaoSDieyNLBk0EKll5y7yMG7Hr3UAFBT7fWCaLIpiPOw5Zw8g
7bjwSwsByD7EOFCNPIYp/vmbfLHZ1j8tgMSjDwhkPHD6mHHkANNu4gx6Re4q4xUguECV9puCqTGq
FQNgxOI0ZOoFpbLGRHOOTnLWBHP/yPLF3wJ7pA+zhItkG2T6ZItybFc9WrSbE95QQBLw/tE2iDZv
tgCZPatsc0dYnqYb8eAEpJ1nytV/VnqkRHuJXZIfXYbcMPH++IY1vLnlKJzVzn0G+293M9PsmwH7
3h7Yn5CEe/dnsdZcd0AZfEwBCARH4kMsIBR09nfvgWLVrDHuTy42Wge03lTvbbEUYraLSn5OwuNR
MUTZMUK91AxMZBUxRqQCouxhKnp3se7SPBkP5BIjNPFic2Spv4+4JbAREh2yMQLukIacnztynPCp
RH7CjWqC/O/XKhcDLE5uunR0hPBld9WnpaZnRT0AtbiJTd0FFANM0/kzoZZEQzsgWcUEt/Gkmxu4
awTQTAnLq+ivHlfRjMMV+8HBkG/Z47M7Y4+inwisMWzzL+hLwjJu6TWtq47HGrVYtaH14thyOSRZ
zV3PqVR9/kEJHQc5agvs/AajiHZyPsqYO9z/ts3hnQ3ZN8gZcHKZsXBwKEZbgFtdnRcvbxoxoD99
nSoJPAM3+cOJPcwV6zE9lBWtHOq2uvKXcbLPq3EM8etues1hBUA1cj2DQnHjFEAi2DPDiz9GWxti
3TyanUtWIYteHgJFfun/itDDKYAydT78C3jnr6xaTSqE2QDnQZgK5IlncYnhjk6lIgUd9Y1nlW4f
FgJFmX1uTUN2bXfvUReacUcff4Ktu7AM68jWfdoJol5tv1Pehr+Wm0/fxlmhbdiRQAuH9N99hF9g
XmX3pygcl4eEgVOEcVmDITgyGJhaZGnEaVwVGokoDb4EfQHSFR/7Jrws/YireJ5KODni3cfH6byX
Xqe1wlv7GR6rqi1smZTJQm95wo0aBv7W3QyIBbUxGH9o0k7yEx8Dr0I8MaRRtawXMBztufbZ4pXN
t/txWxAJMEyOe8P5XGYJq+9/ARo9c4kZZjWfor62Tj0PvtdLkLsBRrFwwmh3ZnCKQN2DHN9KI64g
MDe7jCWzNTKYmXaDuMNCFIqLShHMqXPP3cMfx3AyLyO6GwVwX9CtuaI4H3fPbpmkc7D7NPJnqXA2
LkP/v8F0kewneYRl2zCrT+A4T9C8pStMpMyqXKSb9mbwIIfk9f7SVIzNXZ7OROy/u84xKNVLhsMK
D8gqUTOLhV5H5bFXgHlxxbfm95puFNIGH8QBXY/Cl6ekkGlrqLfMaC+iPmx+pfs1rgmmxWnCFNua
xAIX6CBp/Cu9VpGoRiaS/zh6UQOVU3oSYha97cG8VrsCOFmjar5Si75ki4znCwVnWb/v2uyJrrf1
AzQr+vqyFqJwbL1tIGSMqevDCoAXBh62FGQa6wRQZE4GB1nvFgpDjejjSLYU4fAtfQlYonJi1qyF
huhGzt2Jw08QtQf7EDMB6+6XQh9YHmYCvvbvAVnwDJU2516TOj+nM+yMXB2lQFl+vPldtqkiAvXA
5Vx75OwaVxBliVGvUjCiSs5D14cfyMiFjIAwAcEv5dcIRG/bYg3SaWJuHmeVF1dwX1p+KmIqKo+b
DsOvoWHUjhcnNC5EzfUFk3lBk0uWiAeFnSTqHO5++vmZaGG7bnKk/qxwFsleBx8pWPV/1w9Ieonk
MQKm1rC7pXfuApJXM3x10Dm3P+E7H5dDBuXclWJxFS7+ijnz71+Y597Yhf0lMoSHWpnLSTwGhEpV
LouL9WDZsGbiNAz2F0xVfCGGaRiIeIZoCZ9O9JPUUA4HNkelDEpv5x2PcuDMosGZQRIS0r1kuMQI
Z98bdQU0rN6tckK1Sjd/2EaVCS1bUF5gJUotz6znZ52Nntd9HxorwNSTTUTrx3sk7qT9jYdnucZ0
u93juYYKVoEcB0jE1IbuKwVzeMri3dPKppRer8fJBZ4MYiv9y/ZQLyxhU1B4H6RtOKmC8U863qe4
7N+8hC1Hd1RWwW2S+lHYaSa7zP+gp32hBroxCRpF211BKD1SGKs/EFdXI1A3qIImqzvJFL/QVTPn
18iB0gAr3eaIQQz3TvzS/jTolANx2utIzZXUvFOfl19T2Mb3liRffdhr0zcxQLS7I1eiD2S+9HlR
ZG8ZUnNT2mJJzNas2A9+v1Z/QLMNM9/qsB7+N6HJpIPPZZElTLFFS4wf0paz4sixIzOw5jR2bfgF
TJpELtfrBugMXzSi0QK8wS9TCi6z5+f0wp8PceCzir6zLp/9TRodkvPy3q+kQ5rKak6IWtYoimeL
4kREvx5cSqzjhFvBLSyzBGDvGvhPyKhCCXfF3heqF1byajUdTKRUAzbmiNPPw93uZR3A3oLtQaVS
q+VKCEmJnQH0ShnXnDJ3vjRVFWnfhjlZx0cTHsszaGG8ITfnuTgLh9EfwX4OKSbg+U99qZLEtWgS
8IN3GwDkW3HrxPGgClgpuYTi/b33HovTBWyr1S28Bb3z2tzIcDSA8YH5ZyAxDy4Eea63NWebG+wr
xeos7DQeKwtTGM1+DXk+fNNqjPsxClBtrSRxNmpxI84/Z4RbuRIBY9bqS6UmRmyUZHscDg1zvTQo
Ifcfv8FfqgcFkdkkbmNyrt5euE2lSNdlooTVq5hC9cWiKGnfr+JHQSsDxsCttLWE6ANbFJVGp4rw
cy86NUDJMLdivuxh5dc/oUXJx7OnPk/SAUZFH11LQL67jhEbJX5BzchL1s/kwHT+p2vcAEt7bgrJ
h+B20OhXhc7R7ymcaYn6WrA/Cuc6rkdbSQMaQnsT+QBtgAZvm0XZYquB5vjw5h3Ot+i0oVF1akdS
ol2JYUWYGzixDR+7F9lmj72HYHn0a1J8rJmbnXBSoM58zpcqTJ3GbKhot0uIVY+NwOsIXNQ/qGeH
ghxukyVmxxjfdvvTN06YIdjhGuQIoTY2OvPrVG7DbWWC1yKLz7AZz1IPwBVUGCOk+oY2uWO5wlja
/F9Uo0M4YOLT5HOT2wnYhG+0WdUkkHr9alnzuU+trEiJr7AO8F573pFLXUWgPtvUqIuBVOOGNfBv
A99P1oLPFzaxVmAXGDY9l25eB+ltJXp5WJ3CkhTUKl4I/zKhcZRIcVFv7TD2JyUsmeHvRDkLwNAe
yyTaM9LExMBJeLiZy0Z4qbDLcMZ6OCg7RfUCWM46DN1NHNjt2YdXepTdT3qlHyfvlZ4pH5aBFa4e
FvOCZSxiTRAwualUqGO4yZf2u3gWwp119B9Q0TMZNQM4Cq8Q5lJktLX7qI0RqzCoX4pqB4SAlyQQ
vxPifwtHqQ3m1z1kYL7sVATFDLTWOLhcgS/LV2pj7AYOXOCjmq5q5yHIlh6L9hnzJlmCxqu93Vr/
HRDU9iN3TNT0JF+sQcs/j2xny42IdTACKUo7/Lzx6PG4/8wdm4KWQ3i9+0ft2rdOmT/bz8nFea6t
NKN+Lm4pQsjP9indi3iwCIVcS09E60lbZdQMoN+Hj9UQcY4JH++wUaH2VBGHwz1EVHPcuUbhNWAl
Zhj10NQDA/IEt2tc7q0s3J0Cpc4SJyrZUTrASr7ScIbaYsdM5cLboeRgZhgk1NhI0MPZrCNRuBVl
DZhuR+dXaBfo8mQVO+PTCIrYYgC/5gWU7E8gln6ZOuP2anLO9G29Dpw+N4/MlPc4Z4qs/o37/q6o
NXwVcL4oT7xT53HBi+HGLg/zoG3GhdP3qyuZOP8nvHCvZSUHGoYi+H5ye5+cVdPB1ke71dWZbXoI
86N13/nubXnACWnI+o+WGn1xrVPD9z0GY93F/81+FkgrQ3Ef2fTzKG/4LQEDeITl+X3Ic4eoGcuN
tWpu30g1DEpr/4pz997xLN1fJz+GWIvB21N5SYxkkiFOp6u1hFDCcgBR9yZMTDBStOq2jgad/Laf
GZqhgH/r6Cpv5XEXmq0jOceA4ZbLmJIWWnEudTdzjjNynE4paNwmQFFgFC3JyPvKh0OFMl2srxnv
RPOJpuNq9R+5aC7PvYxMom7uibUO87WiyfEW5OBgAevYc6nfE4X0zzTKzOFrRtLiZP/EYoKLlQaK
bULKYGQuX4c8cB3llC+Pot+5uTcZliNMNe40P8KrGpbiHeFX9H3iuTojqf3Ct+mtpAXVD7L3yJ9E
J7cT1HfvwN2hKP+eWLKAOTTHLFDd+PVYlXfhptfMhTS96NWG6BKB0aDjawiTlKM3EqWzZTO6Vgmm
Zvanj4c/P0pNUos4AL0L1jFSQ+EnHLnKmIIkuD9dzh0acu6DdbdLWd9nkHBJkke7Ml4mV+cR63ey
ZPR2tN50SAC2qb7bXxLMTD7SUfTsBG/JA+PCCFUfKx3vE4mqiWN/ZW6Drjmle1KXiMPPboDBWfBY
1hBbJrvn16aAHo8Xg9I8l3W3Dd3FefJPU/cWgC41DznueMb6OV4vZBDjERdfIlhMqjENO0hhLVlA
H+DK+4vF0HoWSHmvexlgQsTVlu1oubvv+7MxxjtCRswnMyNrrqqlIK7UxboYLcQj0U9R5lOs0uup
uHVibkcqJEhvUAi61W3pPAdGzfeY5Z5KV+tdy6X+eAcxH5fjBkeznNkV/ltPmMhIiyNuOQGLhKl3
ANsCgxgRmf6U/PabmYeukRsMXqT9Wt39xOT9yW0c/CpR3Dya6lf5DiNr7DxvwrcXXBN1q7F51iJz
PAzupuIEACdrI//YIbBT9YQ+lQtq5FgR5DcCwdC/aDJ9L30dT314Xce8AVnTqPQwgTulIvxmYHG1
pZoi6IJ9Y+VMU91x2qLyfQ9Oxw3WWCtTC58VDVZEhJtDej99Ea83rLUpSoM7iO7bRn5PZccwVFm1
vpM6qgULbdPOF30kkrQJfBOuibX8ADTScTlM+lV9HzyReuqYfATt/Gzwf5pT7fI+/dK+HJa+tnbQ
KDoPzPpfUxSjWSzUY12P25vZ3CXIEG2ZO1ZAPFsTUljWActnysaByR46YsXKaR8vwWGyHN/mRDzu
swfJvSpXiXttjhJpsMI9eG1x7oAZ5qRhkoYX4b/v08/eRTX4Ngqp6IGoZGAKY2XhyTgrpN8krERX
l7pkgt3Ys5DJNbovkwXUqIl0JuU4zU0/qhtCmi8Nu84u9/7oxIewpFkUEDNURmrmdBinf0e5noNf
3UCguNjpv6OJ+QA4A6j5VS6X5WHJXxFBvxcQ2SEa3HWi8VOHzAEoMequfvTGFwtd9MRjlOvPw13p
JUd0OjZtUoBt07ejOSxBERsrDo13UwTSnRs8bT82DxBCnGQcIf9J5oU6H3iApqJFgohvv0+wWQ6C
o8yoqb9pfVNEs6Yvyg/WeqEFKKWjOcgGb26/uxLXz0neK0zvt3Ux+klX4Yu6dZwmNFiKldCbw+67
gnHAfV3Zc1HOKPRlPZNPRvST2LmAFe/fBDffNON4DP3LZY1fKM2ulgdCJ4wd7sLzbRzTK3WIt8Kp
HjgA0LTZG8c7NRu7GSkrkow+p9TtiiBEPoOieWMQ2AEU0Ch1K7KFe58HuqqWg5D59bSppD5UGNFu
JQQsqM3zYwNpR/dge5e/CNouGVPqF6UvH0KwDYYvsYOTNzOUrOTxpF3AEWP2kiP4+Pw92PhGOhNa
S9Wjou08nwkNDmdBzL4FrW5HVKIci6hh4qpqLcuSw6Mo/ER27lz+ML/G6tyBlr6InpverdDuahbv
1qejOxv03lV+GTfCH1D0UGldnZowLMCuywEG2Zgtqav04QkZsy3NqGEN3pS0qZWrbu8Dydm7AQ0Y
XX/CvElnkcQvZnr0Mi4nB06z3uRspoqswKJlg0mOosfaZ3k3zz2++epn10mev0LIXsWJyvNHRqbF
GyU2yRGrS7op0kH1wF160/J9hcnNUXXPkD0uQGTPSbA0GFJ9vZFsYFhrqP3tGE2JMq0zrAMiblv1
5tYqwMflRuMX8anYbnKZ3sXsdhLjOZL3seScwicujhY6kQZTaYVQyGJ0Rlz1v8mLOeflYDvSZb0V
0HehtVXKtlNQEDzCz/AaLNVkocTKijUEuZ9xa4B9sNrVC+ye/uuo+DlhhHMlzbi21C3WM05Ad369
Pf+4eXirJLA/8U0KWxVN8EoFINUO3uZWjPPzquQh+6vRlgjcwQ73XJFUqy1wPrWxkscjR6nDxAFQ
OP5Ze2TxrkOuSDorzKEPKuOubQ504pCnfycdLGVyvvkfn27HHXv/gEZ8rjF4C1qCb3H3PexrlBjE
sxn97iLq9T8YxVWqgFrdppxpMWUFlKbdRNiGEWXgf/Bx/OoJLtOZvmRSKlSlGJK33MRZVXxW4HPw
r39G+ukZFog0lgGPg2Y0B0WNdf/WUNajWcbFPfwkVBjtQIboJooAuzET/8637q1rsLpovtdL7duE
d3x8yb4mVxMrN8X8gm6cN5jDGeHQ+DW18R5RtsAE8vJxaT+E9bRFSMnTh4fO0cWD3Xlti+fzC0nk
uC9/y0JH41Nn2nhA9M5LbBVzAtQ8Vr1Lhnp2UK6C7AN7ZcLK31ajKYnMXcoxw+YKoszI7UlZM1Dq
YNWuMTD7+jjWMkXmsLWy7OHBC56dQGpfRxGKKlcudCXyd3X6F1axu6duVLrzGkzBrkMf2oh+LDKJ
0JKnuaE6toQ6er2bX3wHXWwF56fAoQaEHfzoHfWhTwz1jK9IdyXvw6DFnPApnFs0h0okvUu5iIjy
Hl6et64ZaOnmZe8Vr78V+K4xzbGyZqv9VU9wy0/nWadHruRnL+IdOTF7zGtohAT9azDMVMtccNPA
c4ffXZFCKdLt1RKJH4Dn0CLwb9WA91nS3oThyJT1RR4b9i1NFMi/XC/NVJV0UGhjj55A/oZAeTMi
8NSwDiJhmEeJLIBetmOU6McxfS/kGuyILnPzb+TcL8phD3qLT9vJGdGq5j4hVuqhQB1FMdvHFf31
nW2PegEDrs67AqXZEId3kOY6wWouw+FhdendKsuhBmP1r3fXBSXbj1xazqUB+Tn8dkeyB+kB5wyD
0LMkfB4wr3hg/rgG3LVZXhKDG/lHZje61dC9MZ3ol3OpwM432f6G3PIDcCk1Q0JDnebP2iM69hh2
ndfxzXkBLeiat0ht3yjuiLpRS9eDut0wjDHjmotob3zVeP9GeNNzxi+HEiUDoC8YXRoolcZm4/AO
33Wn3PQof9yXn72jM24Ugl7Bt75/Lg9UeFENHTSzNg59PishXr/nhib9xdYrx1Aegk2S/PfUhh3T
VvoSzWME61KiHx7HB9mkC1q+NfdTQ16KQ+ySCxFw8GS36UisJ+7qOh7eRtJt9Ba+ul1+GIXmaKAe
nVEo4DlW6k3S28394liF5HXYFOJ8JDval4lfr2V7NtdcUuq+qnYJCmkTuCIXtp+8OilKjW2cn9L5
3v/iJ3kozM+NXMLeZhi3InazFMBvpC/yAlpsYxkXvMVRPaBqspRaG3sPI7FXzcdFROt7g7L3t9pb
dvvN3uN6zPnoLHCjd6Lw+eJ45fZMopTEcdPhS+xJSfY1U5Hl7QySi8gACSWPPk6QZPjBiCJ0EJXm
tlpy6868DdaA0gsuVQ/DdBP3NlYkSNRIDSXD2cmG/Hqe1SbMScarlT7pQTIrrQyyUnTXhR6h5WkO
V5azA67JE7bdIQ7BFRAP/8N1vBUtaeNBwhBaZVgMrRHj+4OlDFaCxMcqIwv2of4cEfg5DVhP0KwZ
SoHb+4pllKNrXrNuY4D+PUliCsrsliuIhnH7EIZOnBvZobP7svGqfmZqFiIAYsVhuLAkhkx6gpgw
qSHBoL3VbbcZ8n93nbAe03nE0/wrcwELrIzpX+LSs0cxjhxwx8+lF5qxIddEabjbVPslcV3OkVzR
OF2XzY9/iC7sJ2a96z0IW4flJbXTLfLrZ6upUTFCHlO1m1K6gZ+0qR2HLPZbsrJD8ZzjBFwVfIAc
oQnZSENPsoVzlrkgXIZvnlu8EC1923iZoGRW2zJwc2ohbRfKNN23Gu0MjB+WfF+zoVFuVI3JRVkF
40/kxmPSQzipdRh9orrXfhwqozpjvuYMj5095dy4VHAdRBO0luRUpD0vvfXivnn5yTJ+EtoqI4gy
qry06UeZm8Kc6n41yb35KSLVimaUtbMm6oKIuzzdQjJJ1LtEf2upubXFtJdD2Okjsu9/w17+4dCX
WGNRrxmdT4OP0Kf3uTKCxY6MFzgDFWbTROzr00HL+WVNcETZUmu/D3pmNX5/57L1FjQxd957uvzb
FtWz8GkbUkeZ9pz+Nu3MKp1taIaqjf3plf4E8BEyo/OaD6uPcvl6EEE9FErINT6zGMj1/92NS5Iv
LONEQW+w7vvT9kbW0vZgX+M7eSgxk+E/AZZMfUz6RhQFQmaPfqF2373f3d7l4MCQ9uw1jkZXqDLX
BBWIAeLHmgUXQvk4Q5gUobOIOvAxfKztRnP9Ez7QnzWyrMj0tPg8LFw78DA4creDvOrZK3Fxp9pi
TfOvTHnFm++2L4p6LuXsJteY7DokUT6iGlP8kcnbovDutOkENpzZ6P14f94CuDtN56u49K+yiNpT
mKxNUwA9WwQTO94ER0GXwgmgr8ccFKuljGe0UXF3LuxQ6C2HrexLeMjxxfMhaRdsmYMWVAmDjc+B
iF0Arysm5ZV6pdQ4Naed/5NC2qi623tCcD4ATDpkhGGFoRBzaIFKI7kBkB7VCPN94ZNzsUTwXc7W
eycIphEGK5yys01OeGeIEHDBGzKNPbZa3bBoA8XVdzrbXU0Cec127JckI0ZmHJ+cb9gv5kNJAbmf
nG60JsGRr5+kFjgSA/92v5soZLxJ8ay44qEC08K0UjxBdqHncezXnMU8yFX97mZ9sUR8e/+nz8hv
SB5aJrrM++BqeOWvtj0jr7GaH6XzkrFtTa+ojM0vzjlgKzx5qYVQA/zueG+fJCNw6DG+qk7hJQrf
ErsC5S4RUTds3meX6ThaOyGiGHNC16uuus89nRuzv85q7go98Kj0uBPlZYKXpNcGvtAa0B4toadc
k5BzGMWEvGOx16Mzw2MGIly1Zaed5U50BFvcpUv+TEeXU+XB/Ml/UjiH+b3UaWZMamS66nOWUyrY
4nTHB/a7g+Z5aJBDaK/DY94Th8mlRAIDpW70rYaWZ5I5WBIZHZXECertnYuAsLF52hZxJlLXveyW
tt9J0plKNGXbqvZKb/egSYEdc08DILxWyJ3M5VJqDU+TeEk2UaAdKM/LVYTqqBXWq+SdmKCXdIfn
JFDpgP0+TLCGn8aclnLXQe5jaGy7wlAs5W8TN8N8Olv8NRGtvfd+54BlDVtxcwhHEF9pP6H2eBeM
5eamuy7bguBi6La899pj0IcosCx1dDuroeKE07uuHbF1UmwZKFIEfKY0Yckd/VTk8R5uoGTL9d0V
9WsumHCbnWR478qa49Gayq2vCGeXt40bwQK6P+tCoc/HJLuxCQVm99iiQD4xv5Y+DxFISKH7O3Cj
zer5qEkEPaD0UzbWfJeUvSn0rFlQya8USX7t3bhXgsIfipxaewPAc1qZs3QqIoQ+epji4KfCwpsg
rl3bYpROThDdlOHvLC5Ou5Z/gvaPFVujiz2yhKmN/ru+IhtUM1pRALjhlDJb65AJAVSqnRyWQyGF
EmjfSjzJQUsjSYIZheqiu0W3iQWsoYHekGe4QvwNCyZaJ9MmogmPDR5mcw4ieRAtSz4DCzJ6J6ui
D7/qxkkvZfK6b8yVUakAi7CizdopEtjd8NnyKqVhLU1REoSrKoAdDeaTVkSXKa4wjTUT9sJSSmTr
Fv9iBHIdYNjXQTHlv9W4EdVzRCXw6AZ0UH8sYhMt0SG+dc8sFj0gO9MoWHx/Lvf4l/6AkH+1A4Eo
wg52CqYKnSv58dcT4dO9v1dy1MkXz8pgRNZBKQDBXLR+D4vJhfd8SibYhGQWnqDvJ/9k5Cfo4GeS
T8YOyQ/evG3hbJyHzbrLH3dHuGNUUdQCVSTi3hWmjJBpXL4Pb3yfPWqoHTMO946oksxymn08YDE0
Axjw42FMP8fglU9Uh0YjVZSqeYDftFKskj6N84d/g0+Bp5zOAE9MBpKYlVqTAfPOtE8bWBGr9Kjj
EqAsA5U53ZIszGPbxJabNK/f8Ih7OlToPh7aDprnpj+4BeSZc60kWIcJ2MxUlmpZ7uBzasj6X9Rn
5Qw9GBX0vW8z2ePYoAhCdm21vvgV84LqH+0/WHtuzR7oLmIZsgAWRMxdBAyV8wfzuwY87ja23Raq
te0mzzzWfrSxztYZo3s9xgdC/HkqdL6+VvWzmWcsSqJIcf5ai2kElDg/CAmutANOMaGRr8XuDk7Q
XMuA7W9PpzPZOMxcwU1AcK45/Kb2rlZ3dCQaiKbHuuHIQeElj35/YM4w0CwxFvPzA85iucPB197K
l2FFKpKGdOT93mqIIw3wbEmTHNij4AAZzWwpEqKOyniwFGGz1+9qRUOPjyhvIAnQoWKrjpPhxCTI
myOnr2XLPGdOj+n+JBsKbQRNrP+W82rgMLqEXvU0hLI2xW6NZozO/D3pItvyzNqXou5jP4r1ZP0y
93n0mIYcpl/FVeoWrxKKWFG1nMxM3drNg6/2LwbEbAK9+s+TKGOqFM31h8g0tCTs1jN93T5NX6cM
/Rj2ybfgXaxPKdmRoGV79TkT+Lp73Vs1mzbFOMe8SZc5jQ3J9mJ5U8/psZaZ2pQe4WqZk1XVSCyC
LmFDdQUAYWQNPj7+3M4I4OxXHbUcA+v2X6LySAPs365VvAektugOWDepeoQqMT5WVDI5/pFZM5yq
LUcobHxDWeMaz01BvbuMRzDNAYGX8jERvFlPKYqHg1cLcZKdSWg4XkFLGqPXYN9sF0udSo7DO8b5
GMk3/DrwMu8nDnLT2TcA1zm26VMjKg/Wzl7UXTOgzXC6YSxSlw43vpew7obWvarlEEmpMWHK6PTQ
DUm1DILTBZbncOyvrVqgRzEjSzvbK4h7rhjOw3B2cqy25koHCmhvp0WiekWMLzN6GhyumalXKnq+
/1AqYqoQAL7EVBIr7naBWV7TYJikvtDyvstitEkN1LcslDiu78c0JrMo2SdR6i/UrE39DHG5WxNh
DxJ6+TxKwIdRHF10Myy08mj3N6e/Y8Htn5SZwtYEglkQsXv4r/adrMoOxfILm6fyOBUFoHizbCie
AfgKadiabDGLllhlGHZ6NjxviXzpSjgrsWvGtL2g/uBn+Yx5R0AViRqFDtqdF0MWwXfOr35FRYAy
kPOKZpkDwBLTUbeOL8W09gyC+zdTvU/RjPFPr9W6YVOYKzJZSNmrpArGVYD0YiEuCDH5xOu90ZmY
HPBoWmgHNejT55P28LF+6SigaBiFKt0RaMMz5Yj1vNyaqLEzCGO5buf6QAfBVRjypak7IwzAMbbb
j32Qcc1RxdSB5YJ64HG5AoDilHyinBsuLeU4qENlW8YUjdCUyLqr8IQChcBk2XCkudrJTDji0nkT
EKCYz0I3DCQD5YZwk6VWFBeyEEAL2pPzlZ8dk8SFJJLtaCcehvOrxTpV5c7etdHXckavMW/RdHY6
Vp5ntCunz8S4ms0p1PztVgN7sJxO9AAbSEbAS7MVFtVqiSmP3gZG8vFWBLvSJzL7FimNyNKXMY5v
0qWUKaMzezAJb55ZGM5hKMjWN8yhw5E0JkCoWRMMVihehWrwdQTblwxr30HfI4SS0JKjQ7V7jVJW
LdfAoREPoWUVuo3hdezxyvDjlG19AFKQ10FHlCOsdSOc+nHCMJOHV1498u5xWorvZCojNLgRPjfU
oaZYhu3xJ/IhL4mhPOndvEE+c5izQh8TXF1AyKyRA8u2OPWQugpq5Dh2wnAjppwZ7l7xD49bihK2
tmtO0sjQgzNFf4dWMLaSL+uai4CvnXN6m0r3nV0MGUsVz9+zfYkghi3A+ufAkOaO+SNou309Ce0c
60ovhxCkZUekhdhqAGIktC+vwdGl+ww11asvV8HnI6oBfum7S4hBu5M5YZ/B+GdxAYhRXsL0mu6A
86gWrnPXswBSXNo3zJ2881qENO7Upd5B3DnqqwEnwU4R2jJQxJdvEl6ruIXiLKUKmB5v94c0kt5u
4C8D7AwGG0Qk0/b+h+2WdrHutV7dp7UoW42Uox3Zn0L/FYNe2SGqwzyNvLQO6x4G2LFyLu7umGye
x1jfDxm13OPxfnrXfGlEWpC16yeVSoknAEtVLw84l38fuYsV7IiBz7nteu/jtRn73WxiOcoMlrU4
gziZ9+c1+E4RZ27JdQRkuypzDQBJ7lCkRFbSA8oejbgwKnInwQbXnjQsfdNP/vUzkzNFAwxBwJRV
6E3Y1ZxueYec26zt5AcfnLC+cte9I6ZFJDMQF51zRkqP1BKHfojZ3nsoLBbu+H1gEY/hCPt1tbyw
XPPGQ6UKqiQxJC+Ztj1YIgs2NvGWPds5HAjZ3I6s+3vrtd8Zq+uuB5+w7QIu6qZCcGYzXqtXAEbo
ttdQqHY2shOO4MOywFerDudTNUkyur9KOhY8kkzADd7P5EVfDl6p0fBXcBguzOT6Eg0YcC5VGwcr
iF3moQgZ+12Z7PKz8GbzNUQGkLPQugj4fD5IMdxUNHkzoAzPVW+yIVWRIOLwAfQSx4AdiNLtriGT
r4Z59s8iDDh6ODM+GZO8wIZgsftDunkq48+TQq3L5xGa5QNmXlZTrlfPoW3K8rdU8CnxN/bhgXA7
hqarWWZ3ieKiOGhl3C6nEKMxM94+yvb6hcNNa0SqcncjZoY/nPgznahlQ3UXLwPkx9Zw+pMNJvo6
Nodif7F4zAbpEe3Gqwd6POSfkDj16BOyCHvJy6JTDHJCnZhIWsRFu8dBtnEa/1JMfHiz2hrXK7yi
kc2LWGm4/lIMJ1KbAP8fCSb6ByxH9f+ewG10vIHzsLv4wAHXjZghsnWQyq+IWSo5dnYXEcWPvdz0
R34uozoyO1gdDO1911sMW2DDdTi5OkMn4TGZ+OwSj5sC5CxmSzoyB3xdzpi9wNfwp5SpJzxPlec4
RecH/MjCgdh8lQG9zYHZbAd/eeut+SGK6jTONWo5vEl/4ByUF2t+vJjthfRguSIOsSIO9cI7vCTD
X/DYyWuFZRFAIE7Fsz2yMvH7F4FBmJU1Ld/U9slJHz7B11KRs6Fz9ZfhbJX6yuI/BdMliabclsff
hSWP9hWiKBk62ccJIFOKMlrPjanJWtXdDC+hzDvhNpIdbOe6Rws2pHpjHLPi08SiYc46Bs8p3IOI
kVfIRMagpRjpIxU0h3W95bQX21INGuJ5SMiN67vjvL+qa/Ri6WNLVifD6dn6brPet8SO4oWCgSUa
UtjXcZMUv5QByuHmMGgU0WKQeyk6eceUgdhkwSPYPaEjWmeFQ3q48sd+B/3tbnA/I4EB600neOCx
dr9NOJzEm0EftX0M1M9/p33NrMSb/OpbqnfADDQwSAhASbd1qndcM8im5iXD11t//HIVhVxU2dXZ
SuuJcxPLcZTE0FvrGveo563yuMh0A5IOncbSTLSHzIjhXP7jBFI5M7pmj6nfGejECISeEm6IJqLb
IlLL6bdqz+inHne4kxJekuGndBMPVPLAs3Ihk6+ddeSyC7c59dGER//Go5ij1VCxQ7vbbfcuCRsv
3lm4SrJJpLH2AZNRmeubxYTmk1tiPkRqhpLcRqcoTCanFutU4PtX11lYinGx3I+pPakHNhd4Rt85
r2cChwTqc9DoQ8SorLVxGczVA5hi+UzfDrghWzz12snaxWbN1C+bxhWlH/ag2ZMYAEnFkd9nXFUM
ieuZGAqEt4VJJg77o0kE753vPpLM8gc1s0KPaeSfhZZzUzb/VvlAJVdDRDOjZ2/ZfmdADoJtzQLg
HqsSW+whGZwcHVt0+8Fw8bozncZ5OXjszTf+LDa0JBtlr04iioRF+UhHAPF33lIe+PYNw/UVrcsE
SStUlNwTST2oEHWrDYSMMLwvw1D5BqHK5l0NUbCOtV3uCIBJD1WBaRXG14nS7J03QAClMEAhg74N
P7bK6Qvm8aXjmOOlfgHSxG+kA4pWA+I7erAB7VQTLAnUXI/5GauPbqmfERn8cojb05/b8N91x0+4
hN6hh71xkhwSrcSucnm49zKV/J1eqEIcwkYVPiJVl/uHfKU7cHNUKKO5M61dP+butGClYKvk58IF
7KoXT8JUJxBPFg6JWIrvl7LUVTXBuIFUfQfC7eYni06CJcGe9YQS6KUj7kL6+QDJuYyyyGYGc6Io
VQs5xHXMsQybH4SSn2Iud/9da+JdEP28gu5Kfr9Q1gbNDS6w9lHFQdsl8vxl3gChJx77xlEnuf0t
UjMh675ckIqFAG3geQz77YauSfuMjZKTZtn1Kkvf06OfbIeVTOtdOzH7Ixv5WCN50NnP+PxtEt7U
DzePIyvucGYu698pCVs+ao9TBm62rwOLNqcd7Qd/eutjhGDWtVu/xR9BaX0LsK8USx1y3FGjNg7q
TsU2fdfMBvFxLSYltyGTR3B8RTpVPGQ4AltXG+8ns10H+7tadNsKpnMcNJc4tscH2kV4vFVV/rev
zyHDceL2F+EPd8kyIRGb6jJMdkoJZ4TMCqhwWIHIo72H2Rej2piwR2uHrwIwlVKtSYrQeM6SKxxV
/PmTEoIlBEzRPxsEgqI3ChKsjspVPlWiuNaZjHoRuRxasC4hBpeAYBiuXavITAM/ey46A9G/IcA/
WP4V2gkvB8UQCjjcggSKvHWj+U1hIgGOrDlTpGpg0kjr4N7MJ8SrFmnMhewxq9mNca+jqMLYjQXi
P92YLcAUF36ehJ0IriadVGVK0RnLSbHVJZVfwrRSclxZNwbWPp7sD0VJ9u/BxKvDciUdSudi8e9r
CbYh9TszSnXSX8YQQE1m0nvomI8MRlRnBFoRTL+59F7b+enNM2jdCE1kRKQnnnbbg/r5D7yurWnO
dfL1w9d/pHm76lMIXWWaGqzINO90HJNwZTETPLQk7Ry7GCTBYVShp2/OjcB7p+iT4QF2/v2d6dxY
VJoHARPaaaxPYgiWoYktL7aWHhi6mZqP2A6ggcIHb1Wiu8tohifmrwCAakE6UD9UOePYJzhLMste
cPoSAdGztw5oeIovGMfdxHtVKWqUrjpVdDpd8CWVGQCvIiwgVqJQCIIhgwVq8Nv4cEr1C5E0F+zO
otlAbbe7yF5+EI85iHjkIffPUzrQbGFK3wQowZIdvIuPOXhSuV946VeQdp1Gzl+XobCRQZ7T9bsQ
Xll2vXSjK+7q1/shxTathZN7XXgYBs/ua8bJNSdZMfzh4Y86H+auWIDqH2DdEKsX16Tq6keUfMrO
3tZDzGiVe3pEYfYVRlR59mMdFP7gMPIHtRD9yDgu0/N2VEshTJcbNXQ4+4tcKqi1uAZGSuUEy9e3
4nicjKJfPU+4pFsHhsDOBav4Ab4WzjKrrnnC6FoFdoX3xwgcpZqflalo0DVt722hbOkly0ybfLwW
y1VQBfyOKG6C/BiASBnk6u7PTYsdmPC+PcPs0tAvWHEAupjtQdb78XWZk8U7zUZo6sDhaxNfSU0O
mL6S2C2rE6Es63TTXoRsMJdaC0ExAx3/iRwa+MdsEw0jE7JbNBfbEwnWS7LZdzxbE+R6nw921FPJ
A6VSC8jnw4T7ZoN0gE7SApdeohyA0vqFRh0NXS6QRlqPn4SpeFRuCW+a9hnoeXOsPhuAAwpWv5Uy
5tn3krj/RaqY//ev3rR9hJ9H3S3A4GSwSj14wOjOwYPsGI73v3H9Yv/Osg1fckXxmtRyfBcpEi4o
br1mN3hd/z1ZZUKCV7gmblJkWT0KikFxNDPAQ0jcWN7Jf/u6KWAkJ7jldEA5kfB188SmYD+3ZaTT
so3LMFTPlAX4mr7yAvbCjoy6gQ0OiBWsyineChxvO4wjaOYYsiNLx1kyOMe8wCeBY445fLEOFK7c
ATdxjMHHDIetH9Nx1wkEDHiPDSImaWLI2bV8nG+3mHI4c0BsxjimhPttalTNdvJPH5ZzpvQCBX+X
UFzg9ym4u+GhRz4zifs0tw4FgCi5O9Roz7/23RWmtyXyVgolifah2nUwifrBed/JDjfqHcXFUpj6
YaFq7QNkwftPzyO8k+U34sPGFSGR3nyBWDbA/Adja1s8001EkTUb47IMuPD9eo2r/v15RQ5sqqz7
Hrf3WdBeq63oZ6tQfIV2zvuxLH59BguVU9Hv9YR6Jykh1Ta4/xEk8iCbpTJzJioznUySMUnFs73P
z1334BspLMhZ6Dju/qyIKtdLQoUtXqlRhVBOJOEm4LMcIYNG0uljNgdruzoTFBEv1Xn+SXQOBVrK
UDSAzLe+hc0Cumwv+bnLq0OSBmSuH2UMQMN1+UobmyKGCoUNscj7442IukA7qIRxA3y3Wmu0wfq8
GeYU75S2NsZJYCuXNxWS3YItSmyyDxBUeRlFcSZTO/Av+449srFflnVSCEyWFSzrS1qlnUSpOVRx
Fxgc8QoUcAFlILfYNM5utFiNm8qn9uC5wtZY1B79dj6sTiRCsdci/2dkIA9Po6U2SlDiBe4fSU1k
eh41YieyxSddYJVo1R18LEfBd+0hoeKzBoeUjkLkMQifU7Ip3zVim5NN2heEoDyxxDIjraxFGmyZ
rWiSIioG4wqwJhKASMVK51V93h3eaI0AcxjinFrQYDR/X6VKqJDgg5bAToSNTEGdKoRvtxJOYCyJ
zQ1LQTAHUMzmvXLGdHoX42Vv48hLyq60FhJcJVFWf0BsiviSrY8V4/EIXZ8ZgQny3qR39L/gUpPL
fKwH/ns8x8svPYSs0Gm90y8pnWlwWr0zVpsVVjBZLsVmUCGZAYSLc4nEnctXt3/rBrpOk6Vy4XHA
3iUsb9HGhtrVgOornO1QUTq8NRdcWsNJpOXoo6SheV2R3Vtq0sFSZTuOuUxM2a3izfFtONvF28tn
Nn4zAIWPA22RYn1HqFi3EJXF7Q+VhEyL7IDMgycTe+9dU4p9jYmI29OJ8eeFBGwdV2aHy0VTFeYJ
eLfk0vyiduW0o4Nd5WePCK0xhPgftX0t/G5rADHw31iuyG9Cl0E7fIaYRz2p2nl0U293ImIlUSJf
ANpdUqgIuXoKJmY1kcUR1eqX9snz6p7Kz+/jgfQIEKHokic8iW0lu7dRp/u7MQpThR/CVzstcRxw
byrNLl2mapD90fYX92h183YWkgeinG6jZgukW0f2SOVMn6LAjMpj9sv7RPhDSGbVbHqCgoxTOklJ
F2u724punzTTRmBLPw6wEeLGeJdaaiEbDdp7VsSxvIsMkBiT6DM+6M9Rx+0Qp3kcMb2yyGMr6Syw
VTEtsnLsxdnRGGIhwCKZWz/5T96eTTciYQI0IyoNTxfxzb2U+VURtTtEAnEIpRfmA8FTiK4BCEtQ
WRa2/HAEh2lK5LU7JfIV1uCKqUzNyn5J8z7O/JMJy30h9z+VRQorUjys13KdCRIvq95C6DqFfPHG
khKPQv0ldOd2G3QIBCWYSvaeAOQhQjasGrYdHuZOAk+h48HlOR0iXujP8cvTPQHCItJi3+1T9dt7
Uq1nt6bw+ZpIc+YLsItNXOnpCpt+XjazloyK+9dTzEP/WOhKCeNG5s+5L6Q/UuyWOPvhFe7guRdI
Jdfq/mSMNWmHE780etTewdzj4BuhMBqufXJseIKW2xrd/sNwzQPhoSbR4WHX191GSMzDtyrDw77F
73VGYuTmKIUYmQMtn6A68wypTRD+BzQRbDfw/EN43mm7STLKb97OUyJbAxRCUiGM3tDd4Z6Ix/H4
5MSxoHbDMfNSmpS8fjS+5kacf3VXRnb5KwH7mBvV3dKOmz7hg8POAb2XAdVpQbyUJ1u6wE3OceCS
jvNp+/vgImmee9rsIFMr4rc/scZLweQzYI4b8YYPVAgs0wHWq/vqRR5lo0Uija6oWauDgZ1UroeA
DpnIk+bgwN9l608eV+p9Kgp4gnsy0yRci/Vf5eGtvt8+Rg7ybrqiW0pZMa7JOK6QlUNg+JYMfIPF
34ICtZuvMjy/B/IyecFbDL6xpEvfm7zqtVtgymVBGPMmTCBx8JAWMMZHXL8LC85wV2k7WecbdJRy
48AlUymgnr8lFhvcs2+wUsx5sL7p6f71LZz13bCYVcqyWDk6TBkE14Sqvm7Z8usvZx6vX63s0QRz
21SEqSZAFjwpNffMuMy8bujGG77BZIhVA42RIkXBB9Y/EP/Q2zEeRTUgTIxwJ205chUWNPzkQ2NP
RAM/D7T8EVvbAvhEbipeKTpJuW7lXQRnxXf16kUEQcpCPCDP/l6WYgpdDMxEHyiFdqQyzdeRg9A/
G7fOQo19ORJrPeZbBznlbSxlvpAYhQYVf5CvZ06DCKZebYn7v1/+0X8AOAAcDHcHvsRiSEGbllts
ZQFjFLN+xtywH3OiyABUsEqLyH1N3R/x4Ri0Y5tascpAnmsniTwY8kwDxyBgaVHqDw5bG85YqOK8
9dpvjnRxQ0jgX+aunnmml7K1MVouYUmCvK+qireqeISLpbmDiSv8kn309niW2tLp4jmrwa9KlH8o
237Ab3PwrXFWrD0ajXEhMWroKvKGID0KH0zkqoQXD7AnBWo96QVG6R6GGBEyn2DskCQU8eCiE4EZ
ARKUprdjQuHXcMbs0mUGby+6vF24k9SqWumUGJeYWRSgE6O7yCAUL1SsZAs6sQolxEmq/09rRsuR
1O/mw6UIWb4nJncaVI5lCEuquI9+A0Jm7kpIjdPTRN4tYXq7lbCGWqraldvIzBckugGZjh87/R/8
FLRNCsd5/MeBqGO/OPKA2ax9O1AmVJsU0LcIPrAZ3Ni29Z5gqg6tqeLGcAvJBGfOnvtpK0owyTuy
1pTeDeaiEL7Y7cYBcnj6aJ0B53TaUWzKMnZM77Jb3AxsJhjwqg/6vlT5WK20EJ2/lTuOK020PIup
znFm29P00zKygAy251BbVXtxQkdTQLUanno62doI7pOfFcE4rtpOHqW1O3CeB3DfFRDiuZqi5MhW
lg9b2ALbkUoHDAfrx944pmZqoVMe6D4Mn/goFuZj7W+H+F3uM5yRV00EZYn3FH83ZT+doEZ3gqKU
2IECXABHVZBADxPU5SuRXg+mnkpyW62wuMVrCqbzW7vV1DyXX/pjpbemB6oABzNxM84mormMSKLv
cLzVin1NTLlUTLJObK3XDS2BlJ9fAtP1m2mVSeZ58I2hbcF6e+OHGnQj371RwJjasyP41eccuh1Q
qSM2UY50A/8iE2EWj7jAcSu9/mPzyucS2fx49EVVKrxwL3qyD0QFTTRLjOU6gMSfCs9JbDzhA+iO
ItfHlUqz3nfm25LcCvRnIm4pa9Y0XBW4mwTEDwOfo7h7t/gWl8RWVPFjWP2HRa/nvjLkm9P649yu
RUHwQwKRpIpB4WSfM3b/yIQ2uHv1ZI16G0TE4fdjbWgfZV+243INSwQxAukm9W/kNhzRX9BK2rvJ
hwwC1dm6RJ7zx/P/+YyU3nkiiX+7Hj5VKXp7q9xeFkI7hkf0AUbQoaVLJO1K23qvUfvhDEqmigO9
S+3manZx/Q0O6kUMyKeCmnxN6X3tpBr4EcbYB7uQFUn47oq/9uWdrGlSvZQVmiHvD5tBdZ7hCYsH
w1FqSgfMHQVt0XErlApyOFmld2gplIOaooAU90bkzjPGuloe8gtEmRLK3NsxNy5EZH7omngFtjo+
BC5Fqo4wecNPwsWO18XhLG0rTYOXeVIMJavDzWezYppa3QsJoLAZOo7AW6XRxLqw16z9gTgPQ5oY
jR2p8R9yWUeIhmjELPoUQN2QZY5N6NY5YhdyA5iLglm2qOAOhTtCqH7cHFK+7Ime1cLTnBYraihf
Ayw9xPa4Ub8DAXcrPXAQ9y2OwfqxOcNQaaAPZNrwjfAT2OskflwJpsrsGYqFxm5enm483PYGLJP8
J1cK7h6KKGzDEtAHTbT4PI6LP/EJNclcsf/njDJsy6653d6VYXiXvrFuJwp9jVbqz6nwicwPTYJm
g8+c21EzpNkwF7A9MFHCo9arE2laWCxJtNJQkD2kfA7OXe6p/pAIG0Rsj/+65LlaR//taXwgn4Ma
US/3OJgVGBqdxvpwx+g/cW6OG08BB0Jz6XO/uxuRUBMCdsq/RF8FMx4lnQbYvbwqwGpZ3vOzxL6b
ihqftshjt+6hqis6TJYYYh/UKgKbP/Lw/Sp2SMZYNpNyVN5DSf+MPz9CkPSyHtqWXd6g8GWU0OT7
ZtN01Q46DNHM1CnxMuHvVDJkloGpnPcm4qcO6T2iEtXFrSZQ1j8bNA/TMWdrrrK4pL6mvvWosoMH
Qm+yEtYNhoGWKUkxCVsqT3laI1PDgo06B1vl5KQDocv8L4mytUl42StumEIV3sgS3eCu7BlgzdHe
6h1+qVmMOTceMPqJ4r5VSHi/L6ven3KDjI6o0lfWGwupRwMSaY34vk86vPE8R/dfKy3dzxoBvGIU
dfMFu6sFsk8t8idMhSEBQCJbAZSOyXNBMyx88JUleDpDK5+uQAO3cT8zuEMKyyCfMtlOqbgMknIl
+bQMIif+WbNq/UOniY8l/u5IDiFXN2tEMiqsDMfTqb1oni5NeBUMoJYArQazMG5CG7eqjb+GL+BB
u5xk8tNHa5TBAHqvJ8eY8vn934XeoqRv3p7GKxg1f5UpPMzRocgJgEXqajIhiH7j+6E3jVmZjoXF
uQcjrS3W8EthrL09yE03FECpWknFs5/bo/DMJm5ifnywboUncevVPr+LVzIAO20/2DXE1cXAMzPE
Lb+LoHAoztW6GGmhsTaxmGUZfzTKyPKqrZBHvA2VAW3SDKDp+fLBLnlZDejQ/c7yNboJmz/pmfQC
2SULnpayTBL2wDAYdOCnzytjUWsBRwPjHAbMfa0BSShdnMQXKKL3pKI/AphIJAj7D+NjO0nWjPJV
gAD2kJ6SIBJm1q7abUvuycWyGYL9/UB5gat0Qt+Txq+DLAcokRNoY4lsFnKJGjm+T0AgI2Ftk0mi
aV5n74S9525JI4/J0yS5Mx2gwVqNZhWkHs1iqk5mZPxKTIxMy6uAHK9+BrvNXdTBx4Ajy3Q2FIAn
w1z8ha+Ine50xtcHDAds4wiDukD8ZTN83Qr7QC0EQTRBXVmfxJb8uSMK9jJ6pHnapM7AtCVCCJbv
yc1jq15E/nEZPpo95UNGLbtpqQ8NsdI/ZTayulIpZlD538oL5wlgHgYGjBoX6X9tDQI6178jV9BU
WQe8JaBu9+ptqD8+fkWu/nvf41HI2XqwWcPPzau8XVebz9pmYFbeMmy+5mKlBcYJe1e82WX801Cz
koyf9hlTnGLmLYgWjQRSoXwUq7XKVVO/sCPPtUiDkNMlqNW6XV7YGzlhXs7i2AwSyiYCqWdOUBgG
o0/pmZAsqvCq9JL2E0rf/yoWhky2pohpIJHvfwv6FJJsH6WTOGYFAxlZ8NUYcDAafXA4eD8lMoJJ
aZhiV0ZfhOYZZ3O77XzceN4i84wuHZ8fg/P/wqRU2OQLQMO3CGRL5yIOxuZyVp4qYbg7bypdFVDf
t4/xZLkW7ZpUkQjzD2zHRZsHZAWBbf5X9CHWh3w441EPE5jiN+4Q1hZDFO5dIJn+zT6QPgqaLtpA
0Jn7mGsqVjt60Pm8iJtfMUVlh7FA52PBU5w7EXNH9W3mVYXyQPAePDVKxpSocBVThk7eTbbt+hp1
rkg04GKze+Ah5B4ftAOgpJa1in1fxeHWaVwkhNFwaYGlyPblTYenl8VG2KqCbkKrheYIk2edJCUJ
o7Rtw2Jd/Vp/N5J/0RJHGjtVwDYVTdFS1HfcTR5meLG2J/gkV9ufTEPX66D0r94c0REg/h89jUDG
2gEwvXL+exy3IGCtftdDRd++3lve3pCp18ct8AWeJNy28uhMPMabU/UaxGB0mbRO9rXivrhrZVk6
Rui8MC7zWsFR6uO2/+0nsikaTRvgsb6n9kYdcd1fTOJYO4BoCntXGoP1E+Q53SrE2w7oc3322Nlk
WahBpnHEUgXXLMvvYRpTLfrrEKML12uwVwh7wSSNCHuxtOKRP0zXwpEdBK7ZlsIvgah1sniQAUYJ
05fgzfMqMhAW6QonUaacaW7kinfxm1huVpAfScT/5CzPKJDfdCEBaynsQv2sY727K/19QWnLDzJk
o+CCE85YbNYTVqwv3pRfpugzUKa+oOmsLbBloWPE8zPtVJqPnUC1RJ5JAuECCiwy7mMXs09g8oIM
2wWiUDOOZx+hvdbow4E04Sb6PBLDYiUqztpDczSRMk1XENV2qGXcm+yxwv+z5fzIyqmLGrNR6eNd
L+WUGwjmeBB0Hkd/iAFGa0uOK+kJTC94FFY0k9pLtGXUphqdHEuH1O+UQo+hH54OTpD4B/aefwc9
ehquFFkpOnLjc8DelXQTrE99/4CLLxCua28hlsJLyoQQp9h5mBe78M3Ti9cyaRXpI7MM/2GQOVYs
wo4lYza/El6nC28dwCir5r2PsMDhgcp6cpRt5W8j9CqDMwhSg93CGguxQSF0ZshpvPFLJCfAqpgF
zkE50dOG1ae/B8XQ8ptcI7AepYfeu7Vu8zkiV42Hqv6aTCTp5CBp6kfN12AJkHarMijHJGoN/MM8
PGHGB1St/Fcq2akqF+ej1O8k4ycL6L02gbbYr6odLpFabIidPKifTn7kx1kK24UwHJONh0Yrys4p
4gUpyxS+Sm9xuLQGnznjTCRMvVbJw0BAHVgQowOxYXew6yC9hg8+1DDpbphMQPYKHXQJpeqBF2V/
qMI39z9/hrJd7zx8wziQ1OBpjV3CqJOzh8cEa+z6FKp5SQnzpskKfSDBArylWOvZLj9BVjwyS4E+
oMaE6pKJ1Q6KldNyaW26hT/cqNWZG8KCfq5S3SUYNZ3ug3r9L4I3h1MaGL3PETpu2B1GBjFRR6fR
HxISv2ayF6WsobU3PVlMUCojw/8FQB+4SP924PSrz9SVQ0yk2mdWTs0fj/zKvrBXVkS2/vP3ONWy
a6laeGtrnvXgSIFrtgGkbhFpGWTfIuUOEPfwIvEsKetGv/0p8c0DZahlJJGmA0rNvUfPRDnhMpCZ
yJaswua5hzMQ9/bE7HKN5oCkJm7PayXegUEaNO83hhS/yAIvScThZFaNee+CVkOH/d9ayv/X5v+d
nQDP4LR2oNOBn/BL6eJ/zgTE6+IUNctyfyvKhRp432OrV01Czz2amCOkezNDqeMDaAO9/ylWKAwP
80rQIVkzwBjnyk3iasCys52EI7FvQ3RElCHQLmjGSXFEiTBUBIWf4egUu7Or18/+M0RAI4emNvTf
rF6E4HfwjsD5GKo4YoP2XoxxKWqUX/hhozPBjKaqAqFaSPciW76HDpn4T56JEzzf5rTQ/0U9Hxhq
uF/FLmLzDAiXIUhAHP0Q6kJSQRL+fEZuKV3BEYsyG9xa7prTjwnJ+y/V3qhNYPNlMFLEk6OQAOET
r2EuJhYCuVKRkp19is+UdLyS4oUGyK68DKNZaHQeSwDnj1nM28NAhiqUwHNN1SLj7KFSEjqoCqJo
FKhJ6XpLQHtrPV4LzEK3FbvfSmMP1H+blIowRN+8Mmc+2t4xzybezqtLdj+lSbcFtGk9SciZpoJJ
RUCVipg2ZG2BnHN5/J9PL0X8WM5KHGH/2Pq0SjxXvDDkE8ueKWaR0N5pAqfa7L22Q0ZuSbWl9Ycw
aRKuk8HKz+BSzOYKgLoiVi2IOYMno0uwcfZw97MXrfgtCMr5rP8NrMhs2HWNfXyA1E/GcZ1UufHy
KrxakX2MgubZlKhIMgE0mwuI9iRsdZeRvhv0z1XY0AAhf/06RT1uo1iOkkUb3er9bo+zkCb/C3cv
si5YpjUx722N1oRknZ7apOfDY8+XlUucXa/aXTwekwxhjIsJGqaUdWBDbg3kk2K06Mzv772Y061A
CPGsNEmhoVSVA5DBIg/XW6grrnHe2gExM9s2ryDYI3k/Kb6eL6lb30K/C6tYgwpvE1SwVDeEo8A5
XTDnm92Y5iz60Df0u1N/IXIln6t3pa/yt7m27UqiXUl7Whz2LBc2CQp9GtYKvmUL81oL/Ekgswfi
hVsaFxzK95286AOY7C9kFrjNQ6isYjJamF2HopEaw+3Q/iJxVpYi1RpBjYljddBqMYOAqMMfYvuC
LY8GUhXir+p0HU6zfdzR0+bnCEu6P+QwKvTff79wqanNodh5l1TAVwd5U0oVU72VmvE3JVUdzl+q
SqlT7Gg7WgS+yhOgOlWyxcP8ZjgVOfVnuJNQ1MUHCn+7Vdx4v6Uzw3t2AGQDsFPlKwhVreOz6kp0
iJbMq/V/4qhAFIkrTghQ1mOw6nAa4RwQy8puvUz4fXBP+DvtKULDD22q7q5jGOqMB2ZG2hj79bOu
inf613yQ7dZin0PZFlduMOS56s7jTPd7svKfcTOPppTkeauI1wBbKAbfTbW/CC9KRs3NRiLcTLz9
4xqQrOmWzpHIVpb/c0ziIjWZJcIwxIK33XfZOWv/W9VsUlH27CZBoDdIQWyMl/LoZ8YvJtRIlGqY
8h9qu30zc2EksKTBvi3f4j3RYYpeO10uZPSi7wLzFAdvkShg+QsFfQf1AXgkl5lW2z6HxApCVv9F
uMr3HD4cO9AXDThOJ4NSqGjU22Jfq2daIKfEOV+J1C1ggYwHFDF4tgCG6fGxQaV+RLfZp0qGxla9
9hNRoBLYGdu3eUBX8R7+1P2VP71kJElRaFMai+kLw5tr5PMH3EJawubZHFhAieXgzJfyRYPAeZNb
5PilqSxtCPqUkFXH6Bi4nmbJqSsHgbaCYW50mGwipFLebGL/Necc5oiGiis4M+f27ziYmJYo9rjQ
0mpa+5Iy7uNb6am6r1HAnhk+n7awSLHGV1P57lbB7DtmQhZD+QWGKNk3rpoRP395wqle0E0aWjan
R38YmcIS3pVteifxgIehDRwwmXo1q64qMLtRvTTE9MP88v5jP/DOlh41yxVOEf4EfPFxdtAqBnwF
c9chlr13acmbAUxwcxNPllrrSv2JPygyRo4T7FNxvDZz3Joa4jeU1T8q9YQwd4ePwPliQlagHdx+
GdS1dbcSJfEWnadjGyu1DqzrXgX3xpnQWAsZCdSizBilSdSlEaZZdmH088nfyJ95QzBjtIwDoJHr
V7e+Lij4prRpynbIagSd8CguA9CtFyY3P6u/fJcAyx6X9LTqXv06AdNu29vYmQyyrTC5S1zFfe+n
oy+45CXcqQQUZzrM4skoOnQ8SwPeArB/V47tIA1MrMCp3+TmiE5EwYZx5Eg6yeUK4gLZatlOIsnx
pLpmXG8Q5jfzmjsYOEuwg+4Z+/pj8A+hFNVidqZUHFXdXFLhQXkjbXwWw2gQ/qjYUNLRjrBtfVZW
+wUoGk+LyGYXUCcIBa7HwRSu2z3uZMLP6BC0r2TCW4o+g59DQs/sVRQnQhddPDGBrvk9SOXDrXKD
hlXXHuQsJ37RS/xQXKgnosSWKdHsC+Xc1H7lfpXkrALKVg9fPrWbSx58gdrmAy9iNNjl+Nb4MZMt
9VgwLWHALK6+w2boizoFkMFTNvOPAADVuqzqsJE2VTaEjuhpgTgDrxbvKgTZjSkP7CQ8lDTn4BMi
NUfkT5nPkV9maRGHxD8jlloW1svYGknqA7A1jI73Xs2bKCF9ChHqE0urzi0qgD4IVUeCPbyXW4aZ
7wBXJEGypr83bM9xz+ymR51cA54cTVZtJSjQF4FnqXtjwL0lsjYGy0oGf/bMAES8CTMWUH8K5f7s
AquqjlCsKAjp1Vr014TdnDMbti8J8lS3qvB1L5KCAFZuRMNaPBriR6pHEa5Vde13uUL6z5/LgUBc
URjlnm7D4Eibf40Ml/Wz2Ew9Ch8vSSl744venuszxcTjVKF3/5/MqxSHdhtzj85c9GTmh4UddG+s
lTr1fqFWwvUccLZEPFLm0TDcSONwbPDV96ya3dMhgUvdcfBf0YXTA+f9uJo+xkGD+DJ9R18m6XrU
mRAoj26RrSWTOIf4MU0a6VYzvf1FX0OtR9k7qlwH5JxZ5IJZhg9HNBQqiQakWz52Dp8TLh+K/FNJ
MgNF5s/72q9d8PjZjcp7cDrg6w0Thwfr3JyMgYQMy5JLEs+HSkQrYZTusnpiPMy52n09JPx7yUgP
R3PDS1jbmQrMF9VWm1ERQRpaejct6T2bNOYKwcSRTHbCGpUPkQxouDXV62EDwT0NL8yFyJgI9zA5
1k2rqzej093tI6Q+1G674cjBPcxXWOraTubQN+7yx1e25SXyKToBf9ZRz7T2RP8WtciDaGOL6WRE
06xADJqjFDsAbjaaWnk1dQ4+Oy2Z/D/bmiy808DZ1/2hYpHrUI6/Y//mw0uFfBACsxztYmN8kU5H
ozIDrKXdI3/08QmkmEdEm3HOr12KgFCVrGQipF5feln2u0+nReCX3UEG5HLP0mUna96Z9kaLgB8n
9W3U1UPTR3419sDN8JemWwawgIWTh4pAKisjRlfkIEvPGgviOAKu2PbnSJGFwDhiehmsaMhXOA4a
MUJwW9e3F+kzm+DSIbjS4mJx10cm8qOR/OkmbOifOjUUeWaagsqrzqhu7/d6xMqbE7lKO2QwFHHw
OfDNly9L12TTcfhUyX62GJ+MY6Hi6NfyvAMBMjIhu+TjauOVrzRp4SX0VLCws6Edvq/DWJuE6czM
KZlTmlbF0sTjQZ7qSY9zq7gL1xFmkPx8Wp/AZW3OI81P6PY4BbuMUY9VmcZwhrBDJ2rEhBMnCYU6
PvUXTK8sOsyR0DdEB0DYQdteJPc8yaGmyzEEZdRdGEeBVfzbWGtCLhx+tLA4myYrs1RLliTD3cnK
n1P1OvKIYGRcl505vk1hi/Hlymn3ihK0HlhjYbllD7u6Vkqnn3YL9rBsodxsO3lksf+5x5m2sJpY
SmsBQJtxGsykW4NUc56vzRsBWrbhst06QhW7tTIRaHOjY8O0fP9Htf52VwDYWjO3yGqvEdPJmB4J
yTTEsHDpA+y2/BQHBtai51MW+Aij6IhuB++kdEmGguEowBPy75fJrAfMaodxqqyd9onWOr9dZmQf
KLqTqM6tap9Mqi2Rm7F2j8luSPSX9DMq/0RTNRViWBwhHb+CZqLHjCD1Do+0xerwnBqPv1sBRNH7
zQa3fNqk8KCM9iIbw3rL8EfVF6NoclLPjt/ZzJ8zkjnY474pz2GgJ+OxQ9Xx6WepB7bsWoxQCx/h
x1oTUS2XvetfpzGFt1vwnNre8YUxSiOM609Xq2QGUTsERxw7OwYriDgft9Yh1BsWeEfaYLg/hz0C
0sPA0TYAfoPNJNElXRGEHsoUC7N8rinwyIuIQTjHzgqdlXERe4EJ43btkfDRkX2hnDBVKgMaEHe8
cH8EN3+6EcFsxsie5t0OrkeVzD+Szf0CkCbTeiYVBRD3YufWPn50r1ZF5TbH11uwFJhonrn0KRql
CroU5pRWUvq0zIL0i5rL0X2/vxKdvZO+yicFq/kVLKb3hU+Ue7Rq3Nfj+KQR7s2kb/6lO2pmqVbD
dBtzRrLMHdJ8ltRFt1esOS9KLcQvcMjRGXMbouJ7oipAI1zcyRcjhIlccTDYIk1p3A8RNMgbKn3F
7yRuQ7u8O6XS9RTT5MnXDHCQe2trjPnaF4QdHb4RQPsIsO+seZYN+P9iuhoURHHLa/Ac6xsC/s0G
hltr/64qfiFJX0xuLHxAQpe6KARVmFhOoEr6nH4jHXr9oT5UnfCBlzbv/ZjgMs21D+hjCBBKMaMa
5c8iLhPSa1/sQRFbFCwmSb7mUvsCgCjVSpcaQxQs8EEi/78m7E7C/DYfYJKalyUhlAQ/Kd/+NqgA
nPZGwyLFypcVzu3iBe7QqRbOQtTl5GHDLxnnNTl6dEgocdZp5kFhi9omAZKKv6HgIpFeXde544na
rnBeRkiHR+U6QEpCIr6TK1J/T8500UAYk20e3tp95bYl47mjjxI4OpS14YxgvPSbHEjCki60FOGk
tLLgVzo6UJTlxBpUZbYOVsw8jjpm89oyZlc8Veqq/IA977hIsBQG0M3GbQ5nAAQ9P1v+kDpKuuH9
nghVvT7O9+2GscjbqLe+VgUqKXPhTgUK4VXEnfw10GW9ha0Y1PSXj2/rBjSCRnFElQ0g/BzD47l5
nPR63seqti1ea/PgnZUHr6kRTCTw8RdifHvsNEwrvjuzILliJ1XSkYQhV0OvqWNi4Q5uLVNEsQUV
5DU/u6eFDGRK+z7DnCZl7TP9AT9tNBttIWk66FpqoXNTkes4Pii5PozO0ZVLSdbUwJpwU4+JSjnQ
f+nmKiRk2WLw2HfARMN6F+CzD5YEemUTGYfryMxcwqkF6JxwJLLNOt5fb31ngFnaQRcfI3lMcFUI
87jh+u4N+K3wgQ9noEZESOG96aY9PLmHzDQc5R1KnE29Ql7bK6Iw+fdHdutnRCzaNgzTaf8Ptppg
3m0EuVA1NhUffsGD8CpkrnQJKQvfqZHlukGcjQnoOA4VWI36nARz56suhKh2gPP2vLKngFJqU55T
Wf4pA6LxTHjgSCAm9o28Ea84hZw1aIkLRcZTyVOfFC4GLeD0FQajOk0elNt7ISdDHTtIQkncLHlw
fnkfm0s2ZWPTqKpNoecGLQoM5B67sihyVQBm0vwuzphBKcTzwTuDTyBEhnaJA6WsH6h4l0Zv4XV+
HdvAwmC6fYjpBcVj83K8mOqzyhON0qV+OmL1yRrn9PFxJF/zFmZH4Em6xwD5ygkDrZEJbhRaDfaD
RDnVgIwzwfvbFsLl7PktlUzd1TST/Spy+wWz7XVwO+qwIeIBzzZDgZn3iPJBPexOKPTCPtOUaD0P
Q8M4jqp+2nd51V3HCXqhMA7CsWcRP+ehwWo/0k7EsdaUmNlNqfZpVylXyv/XhPjojFJa1jQ8DmDz
/kTP4+H5l1Xqep4J0+p7z+37VvjA6wIFoSBjj4aG4JV5FO5lhg4c+sbAYBwHkKJchuOlSDkWG3Ps
L5i23Jg85Ij8barI6n1aeNhGCXz04foJU8PJlnw8frKa2MkY/AJox9SUVbiSi7L7ml7g7MYG6zxx
TsmQYOxIrWihJuEr29J/9FKV08z0/Su/nsI3g6wid7J4P1aRaRESy+XnfEAZTsvU2ZMDODDIf6k1
C/I9aBV7WO198qsf7fLCqMmXqShES0ag1KrGwQGo0m6oKfPwJfdbaTNyJuD//L4EHstdx/VTjzUV
WC3dNtrVXByY7A2uRp4uckDzsx+oHWx1+ClNy/E881AfcywqPxhtJYT8/GX/qyBxBHBG1lR+/rrg
gI4Dnx/SSPu1X7C8iapeZVBojFbOYzt8nuj2d5yDaIaD7GbmKimsj1eiWbYofKFpi7xzlTFMFurB
88D6HkrjFjRfBOFiS0OONr75ynhfLL7GzOr/0n9P/P+ZMiR/q8nSX6WUgG7nIIqgT/zQxGVYoJoU
Cw27N/L5/GKqROFVux+Ld5eHZfMlCSB9j7zzMIfErYOgSW28XYB5PWcEzGcSJeQTxCMpuQQkHtUM
O+yUqxJLyxfDmHO0OnOYx61Vv/LPRi6fYRhk2OeXItQ2t80zt9IjU/Ia31gM6R0gWjIAAftOVFN1
H0ghtorU5f5XDQnQwB9gJlgtGY9/T2w3uRHrMGtWiwostyHoUqf8AC2veaUlCM3ow9kTU09Foo4n
wI4J5r7Ig9jF8MGZuJwaKEjs53StVCzvYnK5scZlcModRomWbHNcyAzoJAbq1i/ogUnrMuvTb7O8
zOquuDT6O4eQobLsmdd1kGSGU5rr8lFmMihnOuhQY1eoRj0X8lBNXlpcxEOlRVm0hTVn7Q2XDi5R
C2/MT6Zz8Ts0Qy1xbcM53OngD8mRMD7Pvi7/strAkAcZ+Tv7xRAHuD1FY7g5AYwcAUb05DACjFMt
W6MVH4nyHOaeq5zD2QcQevmLw3T+sbW+SGx1waiu6WDP9yNqPtIK8zAv/rSCSU1iM9Em7HNamIGx
SamDyuS/kAgOpOOpkH4fbUzk1+X3+ja8u+YQX2mpfpU/tNv6BuBPtzS4XiStbHQL3cdeHU9qIN7i
3lNLd8FsCBO04DaFqZ6Q7ArGIFCgpdjXiiPdwGEYPSpp5GDo3sEyY1WcPC1sToPtcJ55P0FTDYjL
a/dB8zP5YVnXPIXS50ezUmepGYUjKfUx62panNfK1w9chabWJl5IvpAFtO9ALY5pTF/b4q2paGeH
aURg03mj+GuhpguHvvPxZ6T2m7lrPC0uhQ9XMs+q8vjL1sfgI7vrp+Vxq4xJcha5R9rMvUXwpXaA
MhC38CiDUdPlbRMYCDttZO730P7V0mPVbBG0ONGwcDEjM0CkKxZrLXRLoZrwseTDK3+y5VZYgOFR
yvDMuyDHV80res5AsaDIh+KfoewJW7pBaP14sUmrRitBmMrVmPUHyrmlNGpIkB6SDzabTxzNDX46
5t7Z5J51/dllkA8rAXdfMUD/H3DPeKgSYEbzEkwt/50Mix+oOPf4hP1UH1MDXf4EGRYeUI15H9TM
YCvfzsoy5LIT8Ljj/dFaSXF2aIg90lS3uffLZs6PrG6GZxSGHwE0sCxbA9rvphk21pgYOk/egZ0C
KeE1fw0MOhYB0iJjo1ldVK8qgheLZswFvPaTXg9/VVvGYdvmkwbZAGdROFK8+4/+apar+BXkT1bS
lyCq2H0sR14w5mJvf5WEWah2fo2BglwYqArmCdn5NEKrovoNup3ugZn2kS/1REqiJXE1j7DGNL/s
okzydRh6cARo4hUaZG489/X5jrjLfWpeWj9J+kLLMxeoCi+0z5anMzvZ9T8TItrY4QNglOJrmESi
b5AAf7IGxzeCmCWoHx9E2yZg0hRpAv65YeKaG4p2AVscNIUPwbjGoICYbe7aOTJeQepIOweq/GQe
cgnlbbL6+j2CDMkqXRXWQj2EUDABrJ+S7ooCRJRWzotphMOrnrWTJzc0nokZysvGfeig4PhTJ4gM
nx0PThlV8qc8hgueyfjakxMWZKRUCk3k1xk4qrxR7s3dsaWotKCQMol1pn7CWlE5jbH4L9OnRuOC
hAxcuV+tqRPYHv1eIs+LMKrmbAJqB+HxOhyT5Q9sXF7I8W6xAGLPMDiX7ye4zq0NkIxCkJ683WhA
zOicGwXcSEcK9it9CH1gBfJF5mdaSdDJPdMRnXnE+SgkVLWO0CWS8K9cheiOHODUYGqRFxWLar15
9qrsJa83x9AjQWqWRcOLv2Jwb27w607oGHfbs1KaktD7EpZxNz115BL7vAlTMloIvlgfUvKbvabr
445LKG+HpT5/4fXx5mUIxFdpUmCt4dl9AcrXMYahZYCbNGClaZtetBOafrLbspi1NsY+6kTcAcRq
VPkO70Juz2EKPC0drpUBPk4xxozJKmOVxH2yeNzcZY8gbeGPLsK1iWFfC70BTZBfi8F3ZFGegqoG
U80uyrMVfW8ZI68UiNm1Gha9OjGKHf3V7hUx5Y0+ZQWNY0mz5O6oWUt9clKQFP+iiZV/OK+dVewn
rz9Klm32KLwV8q4F9VDcLuzKQ6+L7JoXfg+qquqhbNdmvInDXYraj0NLcJ0ZPQMV4qkSwdZ5PolE
dZOBymTAmr8ko+Jvpvg2aYJY674h4gMnPL0LD7nkuENeYKt+JFlJYPybfnXrS2xAOqSeWdkGmtBS
ziy4XBdpnEEh9yiaUJLUzZhmvYxUz9LylG8whgsrLLWGrhRdtRwnUe1LEKT65n+0FQCyzdZmvSZB
Y2jt8leRGkOrVnEI/sz/wPQLlQt78U0I2/wut570UNT9LFG3wJ+3Jk23nzLXGqE6dAj+YdNTJO0B
sSgylEQpU91bWGcx5rlePeMj32CKdqiwKLdCO1vJpf5nyegsc4CLsrsHpJjpEbq/01lFZ83RP993
vwtJY/XYSP+ZHewzxz+QkzY5Yi1SCtvJQexSHbT2bQdmZUYbfPNcCvF6i8NqS1+PW7QAaSZxghjk
dA6xwuQooPmNa6kMDrKPWyY86Bm7XOaT7YZYbOj8fZ+Qq0SGHkXR8C2zDgdA+eP4w5Skhwng5RNL
MNRD3n/vsqWcWEEp6kdYl2RGnBSou15IsBBnoi2XuHc1HdmV14IDcoZ25lsbRS7JI8VDkpiQjmyg
Rps9Ykoa5xrFcYuGycvm9nKWqxerpDW27GVLbN4dmj0Pm4hAsFgn8JyBfkg0KGSzJZ/665pez+UK
XpQGuzBgy4VdA81Yvq/TrSMOJrY7iz9dkVRzroGpHs+8xupEVerL1Gwi5Ywp5MHiseUiuyJgz5eB
pTiaYTuk/g4eW7RXs3Q2MjWqw4HHzopR9dHzteCJZarG6N5Oxsjc91SYSRaF8Fy2EDvy/5o4bxCA
z/DI4dilUMRbx4U+fUE+CQULRFTVMERhW4ouTIsFGa7/vDiOkUcdRtb/rG7hZP4QZNHfbNWl+uK6
EQtHC9eAZvs3ew/kCKtcHwLXsRBvYPjlN8gsCvZG+ghn8Mmy3ETMIMeNz0a1F1FOZNABBNCsOipd
AgVuSLTv8dad3aneDeVcRI1S2U7rIg1QlFOwduotxBFhF3ofja6V0LLsnSkEzZakVSxMUslbuDk+
Ov7T3xHF8Y13SQ6hurs/2ReLPumMU3VJe6031cYl/v/m10+IDHsUl+x7QZGP1RWTcQDEehlxpv7A
KYmPEcOlr5qeFViuJWzn9ASAr73UCyF/MRNeaE9YoCDwYYyupucfPVGNAcikH8mxVEkI9abwX7lg
iH/fpNR6xu1MuoKS5BqMNz2jVAsxYPf/BOwL5ea+H+7qhGNRKYf4wfaMY9rD6HWVBtWxRgbL6kdR
ORj+CI6Mvlpm4XDqz7EDtqbAL+MdKknLSATGWjbZwjC0x5ODX5E47tDx7B5gVUZNfCbdDASJSxjb
K7dPhIB+ayLbooC5cO+ixB2/RMEmwS//7X290jSG839DzARQh+uLDbAUokJO9pjBvH306uJM3mLF
iqPqLftMthZK5DK8blOyCZcdgpSLWj8E9JonDJxjp2h890sUbtBBmn16zV2lesj76dPezi/rXJc6
r3rSuVka2qOi1o5xBRYzDT0fLdU0AiVjGlL4tJmsJPeVOVtd28hUG7nsEUOyumHNOQMjd1EnQSOc
tMn8oVkHpnrIRkFE6QxCXcAizJeTjgt5G3qL32uEFXAD93NM9KPgjrJf+uB1sUdQlGVYS5H6hmRr
pUZn5TuGVAMb1sM5iDnPKXhW3Lzhv2kY3G00jkRRGY5q0tU4gKG5N58YxVBLA3YSTDfZavU7zDLT
mlyQqYMKLiZnSwSSmiMeG3070Z/G3wE5+RmdxawPtyE9I4mvXCxDwt2bC8ppIBKeud64GAeQD7vq
9TOk/FoxX9ABt8xBue2BmJK6kco5QQlALkPi40Ec/tWjVhuVA01cIp7uBW+qgVZBpL3KTgVAA6YP
36Gf0ejzkd0zMmGp5yQxK0tM46KRaq+ABn1FDzMU7Mt8+11pgi4xpu5asrQOLHJgX6rZIrnEYnFC
pIp5qKPBCpoIgAa4+/iI2pcFH9iFfKqjIib+Jav6TvxS3BlfeE+c2RbiJwpyVY6LWwaaPVCOSZ1j
8t6KNluF/AQVFl/KzIJRC39HaCbCYAYx1mr9PIlSD916e7RH2T+2LShFGVqAMZyvDOizj6MZIYRM
KZYMpnaL9ekF8fPkm7Ms8Dm4GgB0YJFnJ8ml1mtiYY6CiygO+6epPN1VkeCnaLkOVwg5G8Tf1f5b
BtjbFNVjay+Z+FcDXA8CDt0n2vv7Qu8sSajCSlvRGEblfNalUItgjNd7wER9MM44lBavDJGP05cr
kLVEE2SrtUBB3juV1G9MKdSPGLy2LKchuPdySJXL1UzFlMyprMLWEnlgenSA+wSiIH47/bduQnU5
0ZVrisn+pOtFFfKgPXLW77mPRptya6TLXvI1cHuBp6IoxpjzRLzyODl4jEq8nMPu6deygdMORfmy
1qyNipCaefnSvNoC3i3uFwUbdiyAXUGuhwJRZSR9/CPgEkitIrJLz74en2bOXd4sNMoWNz4Ewa3T
WbKGsA7J8GdRVFjuY9QDE7OXC+/ZWWuxVXgsMdLlTwantk+Opp1lld8Bb+2KF9ylh13quev3wTTP
YcOnfQbk1ReOJrQVRiVUdUdIvWMMNCPZTQzOYjwra93m8wVniCfmX+kZX1LWlLU1Hrzcx98kxWpa
j7Zw8Tq5ISUMbUbY7StOvxLUdz/n9Up2W5N1L6hLLenJTaR4y+KCWReWmoZgQwH4gvvYnjxeToV4
TFY2LsSSQuaXBbVsVxWJeWNUz2JgFHGQGNeJx6DpItgUU7PsJK00UCpkSL45meB6JdvUUzvO+uiR
uCgqoXbGcyR4aMvzFY/rn525ZGcqvjn7V7+zXGPcHZrxR3051+Qfb4e7UEFJM3HZqC1uWI/v4ciU
jPDH2GhYTbLx8t5mxeCnYvQDhdIlmbtBxsI8klErfXLHwADLt1+F6f1px/sIKi1+lF4CYg+fpFW+
ZqdYswSHOgPV1nI/Ox3tF3sgpiIU78ga+FRJ8CYXARQhctbPoee0B5zybY6Q4T4guKIdvDs1sQCL
3XGQXq6vbH29SlCnAG0XQWncCtq9slP9kzJVjDvCB2wNqdMTSwNmDt3bbyTth8PQKcIf3KmmZwJT
zhbWFk5KVCZX6hcSHKSzgZtIAoLq/wKPlcSkqxyU0q45XkvTdqBRNROdvifAJlYpfbxzyvk2jpMj
KLBzSsYzaXqLX3Glraa2/+JfNdpWJFFXjFPnIBvCdNFe2S05ybBfYhkqvEsuwMUFv+Hf7P6Vt7nx
EeslALDg0WHb7wcktWKNru9OHRVbzVp/8aZ4jT9ESt98MKr7GPWpmwkjPHgA3LV/7CD0kyO1ftQj
CiChTliga3banUKL6Bm+slNwm0srAJP1M5ugN5K25seA2+vrj6jv6Bn7mCbZttwHXTHxNkNDeOXT
q4MG+QId6XVMU5uUPgKHWddT+Wus4SGRBf53Dx0h5PGA2QiSiBEkfHviJlAmwOxqsfZQPqp5LrwI
4YX9yc5SPYPtz2H2UsvyCL51KO+d3r2vzHQvktjCXijehGW73nuTb6ndH4J4yMI8Gwyc41E0nLYx
UPQf3OmlGsgfJCXa1Lk19DLqqmiDnTmsOkDIhLnxaZrgDPlQ9QgiBIdg4LLp/X+cI7cp9u6U661Y
daZ5t8aolTPkZ5vVpb9p//jG2H7eqKd5NcbEIdslSGZcfIzbKp7Nuy8DgF5A4qBPpj+mNfoQ+Qx+
bn4xzx2AkeS0+9T/qyxNnzEHR9VWgL+NwV+NBOVXLsdEcH92Mh7Zw5DAtZcpZ8n8bG2FZ/A/9j/7
1eysNpilMPsNjBgRMaAE7ZdaPQWuDqWR8lSvSdexLkHQiZxBDU4puMhohBIOKNgGqjGCn0EtiwDm
OEwEHFqEPdOCyEbIoSqxW3oZHeJYHX8xsuzPQ5FKt5niYLpYaROKRHiTJIVmzRjCZsXVG4uagl6P
SOj5GZhqsCAP6OwvGU6kBVquxOCjidZGWYt2+PJeNMIOG7Lt4ZkLEJsUb6fmxT27httGMifU05fx
cmof9MlB2IOe8bzxN26iGX+e0/IdclYtb3+xpD1IFmRaM/ky7Puy2LYpgBnXwrQqeoHbAvkU1Zwz
k6e9DaYuVfb5zTJUlm3n29eesCdJomSutIO2A63I/UWqpTn2nAgrrMkmzw3iLJRTgaF9q/DJqdmM
07Goc1uUsqrfcAEFkzj13fFaaeBluuAmBasiR71uGpYz2Urpon1oYJfSz2OFbLnEAOmER+GJGfhz
CAY8WXBVBdylF6UzjaG+HfMTpNhaGLX/1atqg3fdwg18ubPX1U04kdNbw1Z/0YmC4n/W+Ai8OjJ2
kBHhD9htdd/A+w8v6rKD2Ev5pAgeqf9g5/nmdiNDAPcOOz9yDBJsy0ixt6FYMhPi7fRmvwVNDufF
RiZfmn7QznGNa2wXZ18DgN7FmrZWga3h139CiI7JfyyHMfNbMDlUFyQBmUX3+NFL6LKDm69bWZi7
JAsloHXZ4N+DDAIwGEEfkHB04ddCS3GvWtqJ5PkRhGHwkW/v1kt36U2vHytiFy4Lsp+oz8vRQ02R
N8BeiZbt5JY+1tdFAyW4Sbnwvqnbuip/J6+b7ISmuy8yWzpRn0qwmOwOw7e1/TPK0FfrFxaMgW9u
+4acMf8LU9ZD5z2WaUwhFOzQHIXbswU7/8dY/ODlIqknpSc+yWJNsgfe3ypq/tI2CMfKuOiUyD+q
v2i04PRCuTpWcKwhHxRIa0qgmUaiXPFPKHymf9fjY33RvQe5WLm2LwpvUOjNaekBFgSJSpdLEVA1
QbjZKWGJU2rTDXy+Z27MgOQCvbuir77/ONyoE/Rz/f/onZX1ksUL0NdbrCd2cQpI8CQQrp+B0d/Z
qkj/fDaZtYIdROFMGxqbpb2oG4ZkOf774V6N4IUmynrOPxdigMTPZpjtVePv1Z+g0s++MFGEfbTT
hBFAiNw7994yvOH4b6nPhOkzPAbQQtj7cBMnWxBKQ5PPAr8JRiCVeSf3OE0uYC+OmXRzThIeLjpS
ZETBpyt9rOx4xJiJh4nNp2Fp3aTU3zkKufabTj5F/2/cJWLTbUIqrKOuDBLsXbVrTcevVZVfyI8G
fqLnNqelith0AH1rtFKIwXsWGeej/3EGoMXKuf2uV86vXb5Xqd3mMNwVZzQVBM7KbA8Fv9NTFfoe
i46VNTFVdXoc2IyHlRZAv11k4pbfWhRUPZrjb/+RlkHDniTR1pTyX6ZiPhN25vOC67FK4uWdMgqC
cmnP+GtSKPzXYhwJO5/QE81eJ3PyP1axpHje6mBwvnGPVRVIXuyfJBXFKMQZBrmqNwJo9oM+vLKc
CNQsGgp1nfHuAlFxtU+VyOoJh89l+mMW35gCoOHcNpedjYxlhgzMnINzlIuoBG45c7wnI9De4cbw
xYk8PugmLZ3JPqIieVl0izzK/RNPVDiPgI24fyqVbMCRF8MZWh2qlB1AuHfid8WLO0qkIN24b/99
COe1RLTrE6qoKr3TmIN6Ic5+rdLIK7lEgELCcndmRn/sWNq5Q12JAVkiAkR8E9kz5n8f4C1nvrGW
PI0x1GR+3Eq3GhGebqGbahxK5/2nulRnFHizpel9K2mPkj5uCHkkK5mfarFsrp2wfX/QgueB81FR
uBiBbjAQEAxEbl6a6VnnEBA7qV4ZGYKk3bZvtG2bp6QLNew80ykFkJTlGsPGnaZrg+hw7L3E5rAm
hnHtaasqhn3wjdecHxz6kBrs+0/29s3gnnc8OfkxHrp4vSf6afKoiQSZ1Qu/XPfCHANd6YOHYjbl
MtciVquymlHq7Y4qYLXaL6BPgqVUZRGqIRsR8U3a+7KLM3Gr700s7EK0t1vLMsSFv06gxfJ8JeEo
OKDKS5ZLVGv/dseKPIFSOE1CFrt1EY+4Fub0s29I6HbdPQ+v7UP07NvkPs++TWTps3PDnT6Kb/2y
MDNVRO6/7aYYvxUQgoGQIxa95f/ntAXLVAWmAYc46dabI3da1NGq0HY9TqIwEqkaN59n7XSuyXOt
JrCYhUfBq0jdGCaT7lqvzmiJSZUxidAA8RDauB7alYByGvnHn7UZTJVVBxPdd3D7Ib4KlvnemE2D
6J5lNO9ic0qD4yCmwM2z1h91iFo/xpU7gOR37TckkcfIf4esBM7kBoSWR9hlojC/RwAr61vH1RQG
js2loBHEG7Gsjs0n7OK7ncEwZWYFLtJOrJZnMb+zybMczm1YzzEynDJRzlwEZPSjZkNOoxQtQ32V
Z9CKQLpzAkLnZdfZMlUt87BHMyqcVfyiI+Qgx3zzyEJ7XIbciKRV0ROnrfmgjoNk5C0kxvRdSGUU
zaw3j291GIb0ULf1kapuGtL3YnTs0ivaBBlv3Z6ghMZHdfooyy+y6GGLlHJVBNk7kSbPha7dpvwi
Vae3SBwoMrABuyxleSjFG28l0N9I9kb2m7pQOZl1BBpq4l+9BRT/9Na+lVdVa+kpdPhF1MzZ7MyY
ygrZrHaOYEubm7klTIJVST1KWHlN1x0tHbWOL0bDa4iAmtjCqwrN8enoKKW9vEPwnxHqc5cOPbnc
phEtt7ut3OjuNIhVHZvZnbMDHLnRzjCorLuJN+r+Z3D/H9zZLwFSuF2rrw7EUnS9XNRUNR59wSUI
suYckf9Ww2tJYRaBONKOh50ydQTDs4qeJAh7cG7Oiep18MZM58srCgzSWaDxtKpGXGwFh8V8trf0
QNXJ4MHeAiHy2VhV0TD8fH8Bnv4P7agiY7QrQVMV6GVYE4KwBcvB1U1xJ3Y57sjnHg65zgAgWEk9
xyxNPGsLNk5aJkiAwWhEJWK0nFxP48v84euDPwrh+lPscvP8No3qKrac82p9iaGhUKwvrFSEPsj1
w6fukJ8/e0inUSiDismugqnVQgHOugm7rQChqdY2e6EGAVNfJcyvTzOVdh54gJnoQUfJJhq5ef5X
/aAtRvcmrhgjZbSh4+tChM9yPLx6sfbHHC7ZkhZZWAP4rhOBXdjLej6znPK4LP3HAccbOzvm6se6
ptR6HCSU3bj1yLxadc/s+YbRBAED1IfCAdVgWjno4ZdWRlkzqHKEpwYA3srqcK2lEGmjZcPTPn2U
Lz8KF5fVNFaDECc8qYfTjRP6FTxO2GM2PDTQLevnxuhNgl0SoBYeVkbUmdUhzvprXJyJaQsfTh1t
rP/Fk5Fsp9+l0Yd6canCqzBLjl6wyPh/M+1eE0saK49BgH/ZTRqkUSaQco6t4NZIWY0bT3QQhisn
GeqbBjXG1/3Jsx6pWTUhv/fuwohRAYN+8Z3aYlKn1+pZKKxGGLX0v8jRoYFc253ztQKN+MqYZWNR
qUS4+OWWPiW5PV3+WYV2IBrU1u+XTPSN3V3SqH+dyTxF9GODWrNYx/pE1X35Ul83COWbNqLF5pB8
IE3WVSKUOOnZtOhoIWjPEHYMYCrwdFbPHNoxTO473wtFinTCGhtvxnEQipTzwNUAIaNzzYfnxWRT
0cxwYfnvLOgzKoV3YBBdTdgEz2qNpwkZMfxY4JBj3+LAhVE2/UM14cQ8H+yMwjESH8Wv5YdsnK/V
X9ZWIkrO6HX5bsGx6M1+/kWmEv4cEd6TBAQq1QmJ6Q2z8cB+axpNgqA1xGKiuzB5k4yoOEhZvTld
46B6uIiXxI+4zWEHV+BFQiXzVxgLP/r2x7RUwW2jS/UAGCeShSBF8zXHffcKIuSjhczTmVF5xIpX
hE7Oxh+PXZlFQRJ/5JeXmbLDqs1oVGEqn5QssUufIL5UPwPEdAonHwOy4yW7AI/pM9qwbZYtCvLV
xDx2NrkC4sNx+3x/01qAHoEBlyPWlCeJpJchYkt2kab8/tLNGcS37ZiVqN6hJXg+3M4lNeBrCMos
2cCKPmW6KOZEd8gM2Ojl7U8GZffHqwghzrJXFXiS9hVj5JYviLQE7j5EYDG8llKPfKFzCYvhL5ey
wLC4MHa2fHwEU/XsET8FBH/+d80Mw/3k54JF0aixwI66BsXynu/alr472Ns/iUAoDs2ryAcmOHZ4
mgq+lL4PbTb7jSX1J3qdmvPTZdcSoOe0/TS0WbgLUP7qXiR3KlBPvJDOom3dHoeQ7+uHQuTNpJ0T
OdQeDNjRSAMtDWBN33OWdzFf+xMd/XWZChuAD+LdqYtSaYNNKHrpLvj4yw5VWfs8vNSweOVLOWVT
eK/+HLg6iSliPajvhPEty7v+pgwS84rE+xNxOM9JavsSMFy6V/eMH8E20AjLzBywV7bRhwK3ZdC0
bKsqjOpZpF4n9eMtr7vaqJRTqW669S63UMEWa+UZqAJih3kGtohigr1bqIN16nP+T+oREItbf8HQ
wmvmmlpg4zDsa+w63mNUU8poetJIZtwOtdPOJbG5qPTxkK8rwNA8TTlK2VzWKunmkS/SJlxRgbp6
3cSLLnp2h93MHejB+S/tADC8AcQYi80fSSVjxm28CBUcsCbW0lVA+xCBf5jRlTfcjSU7isir5Km9
Npl7Y+As1EpRqwE2mAIN8P9TTrKy4sES5aHlha48Xc36y2v2ByGXbv+7uWE06MuSxCHsreEu7n5i
InERUE5u5dfCKitfDWT0YFIlMmzTV7uvuo85emEHALFD3yoYLXt5PGEY8Nkg00bdlRjlEV+M6H56
o/IFstm4WZ3hzxicmG/Z9mT2fP3dFZLXXMUobYsgm68cpLpvfUTp4td0hFq24/zgD5iQEqtVZ+6Q
UHUyEm4XTnDjQEilR9e+Pte9d/4NXVU/bA9RYfYgG22kKLQrLY6mG/mZXOShHxER0pVQImcLL8wA
LWC/Gqi0QTvThsmd3YmgFANVvrkePq7l+d0gihLKzTwUIiAgaP6Ql3pkgUSayul95iv+m5erRd5H
qkqCmTSRFpHN8pMSQtLa7QjTVTPG8ae5kSbT8l/80f2U27cOCdb7CwhWtQkeWr66VSz0Bu1nm3h4
xoa13Hj4Wp0thG8OrrdmTHvvc4xRCwxkoHHaXsL7TMW+FuShVMDr1RntYMY1LRKXahqIZStcKI0t
VFiLLUJLCecfUe0nEsxyeZQxbitNe3jR4iCD2oOHvE9VnMzvX9s8xK/cSZvBXp3MXor3rX9MZ/Xr
XGOu+ecnTGqaV6DMkCTrrmM9HSPqbKXJ0o5RsiHy3Q2DWcHPm5T57he8kZB743iYcRWkU/wa/0TK
bHrWdj/LWJO3PwmWdFDjc7i8cb2gAudC9gGDdencnYDhRt7jkrEjl0ewVzXJoK12c11S7zV3KLiq
YMGGYFFsLM6RWKa2PLcg1Wh4C4I+y0YyoKaZqHnLTLt1UqeDK3KXJHUhAJYTvJP2K3MUCCYHM0pU
dpYvonzfsJyPfrU+W5Abt9uMZXfs9aFk0qBiCXoVwABmYTJxsuAiiVwryzomzBPyEvLWLpeJQdMj
IGq9El6rdy6p1769uBsMuBwdjHZzuxzEcINKhmPPIXZDZ7nwV7ymEKjJ9MLQQfpXmXdbs2YuO1on
74YqP42g77gdgLepXWkFU+VKvPgS/Lh9ZDoTY+F46t1RHiR9gHVduHQqnsW5Nr3J1huRKxY+poc9
rWR53Yf/Ux+avIunqpQOZHfT5qddSKerMSiVok+RxqtUZUAF0EXJTj39C+s/71vo41w9gArL5Det
r4HeEedbQFtTyVjAah3tcRfaRL21gqg5OpOmHH/FbUXY0YVR/4EDHFPyRsDdnggRwhkq+Tvuisuu
v65PJfVf6xmVlz7+5LHTqtF2uBWqYZ1VswqJDhbYhNMnc3RvmvQ+92Uq+YyTKWjRDF509K9IG6Nd
j10/1vU6vv/T8uyyjE3Xms521TE0D0qafUP8+PqzFO6pMA9RYOVtILVQH9u0zXZrwe+DmzaLt8V8
Hhvru+ou+zVhiVyOOT4uLhscDQb/6ci+qiloGhrEbSJ8usKAwMfLd2wfUEJRO72KAsThi3OOfWY+
N9mPFFvfHOYYBwVQsILx4jErIMgmI+MI6UXaBsSeVJWxDbKONyfx9dKdSaISzBeXfjzh/dBqKC2F
Fs38Tf+yX8FMSRPVBnN/giAeDYGsVj6lzNe6X4OAWVy4QLheZORYVolROi2Ng7uYGv1kofSE0pKh
OjJ67aXHA8w3IfoS1nFnTJGzW2JbBXDyj7dZa3M1FYayPnVrUCdoQXqxdcrxfSOVgf/55CbAPdK4
fOSQ6E72ilfGHjfaJr0box2PajPQloTZamNbKW/gpp5RoOZ4hEv2JDdQ6TH00QarXpbL/U/2RHNw
ujV+JRrJenYxBbUeWGHLrEeJrx7WM7/lngSbSaHsrGOJs4KJ3R/QQgO9Vp1L9ZPZ56NLHJxk6Phv
2Ju51iqN0MidyERqu4QM1EUyNRhvtyRm8wUizgvIZ73ogfAlNVeGLMumix/GPnR2tunjwbn9SA4z
55eR1TxuK0GS5xk6jygMXc0gG1i7Lh9VyTQ8CM2by/9tJhMnS7t7bmmbaer9K81MpLeegZFqJqTU
vglXnGPBK98fCHTWPhq5Am88lZ11EelYIlOKYtA+gfbu0JvBcZqXt+1LzLRfhEWrVuz6HSzdQOSG
ZpJ/ayjZ4f8f98Tb8wLnLS8MYJgBhSg1hfOoi2cFdn6SObXb13AFkQ+UJrLaF57RuY8Xdye9KeiP
f4ehdt+27ztFgW93ktER2Skq9U/MMPUQ8nkuviLYOr++yThVRSG2XqOBr8NGYcOidYZvNfD4TbTz
e/o7+n8alV+Kv7PC7cjcRNNeUYCcTDSvDUARnW0jfyJzeS58iRtNA30g+NIwSAMBQoyaBeE7n5Yr
tEWigj+AhxBH7B5wTNX8e788wTK9wvR4bef6FcO/4siSlbUGcu6DdYkjKyblTKoLgtP7yHIMv3f2
dmgFtW6SMjPadJ3q9PgjC1AKIxxCCW71eaKfiWO2YuDA3p7QjxZFqnohh39RhsW7dbJw1bpLZKz8
eKZlweoyrYBBEEPfGc22WsJjwiDMXSVbwMryzNLMvwXEVdwrBPxLqG20K19q8MB6gJiiv+LTLPB2
aTJfLoydSn8CtZpfxmDyMGkv8AqTiXNFfO6u1r38MDsXTTh+9PBCYxAsAA5C4R4Pah7+7e3BK+Du
Yuiow4ncei3ySUcNC9xn5jAkxP4SdriYFbOlUgkoUZpSMKh+Af9Yjo1VIZXmM59dsVNTkxQNr/og
kITU6DLa8tcmzc981PJthKuH2A827lZCBS8gDR7JMY7TW+KsAhaNW5dc8KmrEW1T6JBe6YCVfmyp
2Xh+v14xhCToc0X5Wy1MufQOL5Z0U1YpaGkOFkWX2aTfmYqk6xqTQ9FgMDRTRWaHDH/cBYcm3M9w
07mbgqE192XwayqRW51us691EeS3Ph6Rpde4+R6ttFO2knRJQ5U80CQ8uTMBZ7DHdJbKVO+WWQLQ
Ez+Ci+abG7QVgrRQYuyOSzuIkEVxqUfiA+hJVLYOuxS06CogJj5wSy1vXbD4l6oBobSdN6WBiQs6
8amahhjDtcY23b3HIjXfkNO8LPRJpKZWfk3+EWa4yVFQhdjZ/7sCRiLINlPh+/GIAqP+gySAzH5m
J2OCDB963jMvELIqXKq3XK8jFi/KyhwVcuzRW85H2LCI4E3soQUO3EaT4MBDt8FFsscaWI3Y/fws
e2sQeOoKuQ1cAGPFIiUF+6PDdvAIw4EmP9yw1MjqQh3tj6YEYd2ry8yik4C48+Z90XrCT2a2tZuI
A43p6JhICNd+h2TajSTd+FZgIn0+Fgd0iNqNdPv+icyxPKrmW6UX17rTZxpr4e83Rhlvx46LXbxF
IHELCL5YioTO7d3H5lllbf9NOmbyQBXv0DPoH5aNdgLUqp/mC6g6FJ7NODWaSC8dc0WETAEc6lsK
sVwbnbL+CQ9tC3RliQoiLdN0H8kSZS/47watWtdvitDextIFXKJZbM1mJjYADYx133l6ICYnjgXe
AUByiUzWToOFS1/wK+eAc22jRXZLQo5FAldv51dAgolt/KXn3YbvRaQT18v/ZL5qpiCM0HA23ODb
cdwlQ4izz2uUdNJTEWMcQALr8YHnrJQXPRkiC4x4k3GiEbjri+FC8Nkst2TkQ6I0P857yeCwwWH/
UW0rs0MUKXoZqitD4eqsLLS7IWiqoW0c1zom8e9XMylYKMbB4n9pFWY5rtDEZemKR8PhcEN+js9q
q05/jurNZzNzCybrFsbC/G/XXgQJx3bTeykCdp9MlHYXGofMy7J/wRDH+W4TxLCB+epqLqkG9O1T
oKNpMAd6tgrQbZO7ZwpRau0cf6bjhi3zSm162i9SOf2La/F+WENVpAC1OP5Rgf/2NCPjCZrXs1dj
QWdpGGh5XgSZVz0vNszpncoGJAJwUSNDq1SmtrJAsTriauAWVISnPmb6HTEuwYd/2prOgmC8oQYf
4y+fcP8zZmnXP2F8Tn7MlAUhBEp01epdPXQNlDQomb2zsNxGfwDm+iZgAQ83r24h1K3fHL4CuWzc
g+jxuDcSNxxs/jqf62YNBceCwY115ASERQRkwR1iqtPU2JPfm+vkHnwSv3jC9pFdZVUrkRpXhRvi
SX761NRmetHi9n08Pamq/fCIvGxM+E0cOKifLJkQEr9pPyCayiPsxoPa1c7jn30tB/B+NvAfDaMn
1dEfuuiJzbHiSZ3tyRTg1XCzWfJ4ble61krHZv5oUZplqIsi3R9JImDM64JghZBHwvYOD+sEuD4e
bU1dXSeSTJa1IRbIjnCRlIAg/UPWwWoNzRC310uCkAK0L0U63rTRC0mVuB/7a1AFnSepUwQk++xu
Tau0rwBBPzUF9oy/XeIHyMMtOM02ipmfKYiEHJs/X3hjOj8BvyE+hGzdwgoBnhfSZAzq1ded3JFL
ufkCvPe0/P0/e0VDa1ToCRb/JUeJux3LCSeDZDo2XvINKDHvFQr1PdAy10zoKlpBPnPC9zXzMdVl
kZ3MyrfQrSaIENThClqoUklumdkqGb39fpOhpGpqrvJL3tXzKONwVb8euIGX3zqSivP1PBWZK47Q
6O5w3hBfOWJ4TkVtOQK7ZQFFoe9IfrDsPNMD1xpi9lvqTh3i8mbe42hCg5sTE+vnEaKAkYCQ/j/H
gsqErklTba5jBX2kqGG7RPqIs194KqKAdnVn8Kl13Ot9JpambRRuxPN3oXErL5Vg5pm0JHGAc3jK
T1y+EvF9XqKnUrMdY9rrzAWCEZ2yeXPW2TkqRKMxmjd3DW8W/w3tjtGl0iFDx404qgyPq6IHMMOK
RD2tfFMtABz9HwoeYjyCiaDt87MSFOE3fJ34IV+Nj+37qVdWyCFIi17J1frVJJRd34hyBK64yu0R
pt5ZoXf8vaL/ne+QVTPAk9k5A0qiWvimwvgqDTmZzQ5cSPsmL/FeDG8lqC3ZrsrpTzObSIOtuPqx
WvDiCjv25sHD5gfLyyQFbdS24uZKt+d3M/veEK9HamYp5Ea8e0RgfMxss9jeFnXYkW9vLRD1Txva
Otacevt0Bz4hNPyGUa85wGatfBiFIbrMNauaa29uR/qqNB9gXIoWtH8KObm7b5kC2QeaZWBmlz/6
9KhG31uVwkC8NtdkzEw5QaqCLhmUDXOb/tOUUF/W00ihJ37rNB53CXr5MCQmW605K+FW9D+9ziZB
ZAJA0jLCO0bXKqUv1kCAQRKE3lz+s5Eh5gOZ4CZ6EKcV803neTjcU22/6nEN4q2wCi69WBQHBUfk
3AsJsOy6Zo80bO7/r1eCzFGagf08HtgbNOJQq/Rx7kzNATDpHLL/R2kx46LzebTT3NZiVJXRC/Us
Peb5/XjVlRKVirYLYkgQ1M90bxxK2hDIbde2itX6ZlaXrxm5Ov8KI5v6ZqzNA40qmrCrfWBOuI82
BRg9Fp0E3zX5bB7Kenu6C0tekUpaBbSx/jk3+tO4ar0H1iieObT8XldlAyN3hR1iHvRb4WlqNGHY
8/hjBmUvtR5XOv43OaQfVBSE8gJB/9TIzMyb6c5m+6Eg4JWPgPvU7rliVwp067/BAb0fObbLpMpk
2pYGnFJFFkkwKvnHDxAEMZtBDf7Y0B0GFzCX7NJFWs9BifIEMXZ9P7cO7jmOi+wQHjdzrDhoskNN
ltvKlnB3Vose9i/8gpoMxC9NcM9izRMqE5Q1LPtN6ulWIGU7WEfgv4hf5WbEJhnPxA812DyMlcds
611Ev8sHwcvGQNSwSRfkDVpCbXyCldAG7hENykzb55Zh7liLAV9dRQM57zWrB9JpFTiQN708ziwB
6CsSMcFdHpwqA4i5lfzjMaaj3f+t7G5olCHgmcWTSAzeenx7xXiCXdB7WC3mYxsoJdVgpYzQWIqf
l6vcJVEoJ5B8u8QYfPBJ7pksBQmaJhUZyc8OmoEcs8//ONXTpmapyvPNaHlN4mABj4sB5c9XQEf3
jAxz5LjAC+T1AqGmyuaE7FE571MfjlGjcw9QWftASxCWOE7i9GYl1oUT4fK3a+zqYLzt233+tEHi
PUGV017W9rjrTsUZbwFHXnsO8KAnAhDbGWyj1i6IkfMXpC2uH1CGt/+Lo/1xycpKEIhRrErkB/A9
CP78LyFiJS7goY/cKdcksw4YF28dwe9jCkAMdZxA6fNJkDybBFXXQTxaM78OExKEqcEij9hPMA0t
6/mVkMSgmO9y3IDX6MzLhCD4kXPzwTm8izlOss63fAOUlOyxyf0MIxxNGLrK/noBf+T+L2kSWqvb
O0UtN6ZKrke482W8OAwPk8n6vmTbxlZaLYP4A/VfSzaJogoXRMI33WlTSqDYT8pR1XCMcRsUWRj2
f+pY6POvCrStGlmwAwJTPXqbUBsiIxLFpXpaGKs+K16ZO7KbJOa21mdB3Uo6ooz1MMLOSu7W7EPg
jfxpEkgIiAlECTNX4xMnFWTik7MvG/kCq14+iBTL18CkC4ZMEvvbl5fkH0Lon20AZRWyANs3BWpr
i7OO4MOdgoO9CcofgAUC1gZs7opZhUqSxeKP5D+XI9+WYfm7OPfyvGr0n54yprqSvWS2eZY3RU74
ilPAQC5GgVTdxC42zbLV32ILXkJs9ZNv3AB1ms+a5k+2plVewa8T31TsPsKqRW6BZp0qvfxlHDt7
0GpX7voAru4CUxzeWuKgeSVwnDdEoGWmWi8Br0fT41KxPo+oZ2Y09YTXm/JPASENVdMyr8fFWBEW
dekxSVWyHcZ5vHrcxhOWjj61XntZnKJ5yB9WUAZfjNTwJu1KQIesGuw3WGO1YQJ6jge9x26LXnBR
333g3uK6XJV7/D9iqxI/k7DiSZ/ZzZyzD3Wd0vywxTv4Ol/ScL59KeTPtOC+GV3la+KHwN61Fh32
/wBYV6L8Rl3/tpI9PUXueygsNCPb62ldvGRNJ3aqC8ipSFgxH+Z5UTqmwJI18OfkmMeBmvWXt3tM
b2UUqcvZG+WtULJRaIxEwdbuOJJiZFxEjhqQQf6HlDokCrH1JExe8ynRaBrq1LAdozhZ3UG8wJEL
uC5boWIesi8vO3lDccWPexnkLMhoIKcTvh5mw2bo/+ZXdo24mNrQVzyYgt/Qu9C9VOx0GxGQ1oAh
wn2PEjEOSXm8iePdPtpL5Wp8fEobrlooK/T7meIyMiYCQznlDSDEsoJN/fs369vHjiF8Iv/L6MMq
sjufjJYF13r+b/6OIruGWgz1HgsNeRrCjp/2QQpORmG8w5t6xtNjYj+3sZCECGcOk/rOeUPd46cT
KWONuPAIytmhVdYl3n/w+955h/QU0M/HYEoui2yZ5pJJqDOEeCM6b3heObJ38u0YlD4SvcKQVf1K
njuJTSlv8zyLgbzlF+GO8aWBSCNmbFwKnM4DXJrg3qrCFSwWpgefko5q39PPvprex5YOesLtmc7y
dYu/bjTrzTxaWq7cLUs1KAlusQAU0IOwEuN0ufCXC+4sn9oZWTbQf2IWSrQfAQFWpPgFeMZa8qlp
4ak1zc8JodRNH+VXwFPbhLB4Yc4rf7UzYrN5yRShfiNMNWUXFAy4+A4RZa0to/40Id1Hs3wdMiRf
UITth0xtTV68dkQQWdeqiN+4fjMdkqD7WofX/btGUPuOGT1ZeXlRjro4TvlMJysqoS3KZE8005wP
P6raAWacVZP7Npe9+64T9qkzR7kgyL1m7r/0yzrd0FUK23xZh4O0g9semectgJFfxVQisAALa/KB
ze9Jww66ZU3IbLaPs9TjD9NFRjPYWbR3tCHQGhyKszXAp5OKLNQfhsN24PEYqqbw7un6frRBtq+U
NrItIlm2CwBnC/NlYgjA4jFJRowWJxV2HHJbZfu8SFy8a9PBbm5cOtUQ+pbR6MvVBh/rzBhUFBuX
hkBBPpyYKgEPgSvyrdW6k6saS9uDgkqN+XSDo53BW82M2NWu5OHtGsHIU3hkEhADdhjwlSUmblHV
lMLgsGY50Loi+KwGGBXCU8uX1hUF1zIN2PjsJNvfd7D+WJ9z80/yLnWVnY3FYIHgRz7vA5WWMujH
7SzbTO5yaopdhdSN32s7B7dA4LsosiIuQMNC7n3IRdTmNokNDfOUAazI2caaThsjxoPdroPV4B4z
w6eKBjpK1QTdV1VjMEcMl4QVhQCEFJV5cWeTy/Y+AZZjckJbRHL9amUQ5OLWkyjCCvtvxxT1lZQE
vP71v7JqQNXJVKDk/Ifh6FDAJ4ipa1aaTD4C8XdGoKdJ0Hno0ya6PrAWHbB6wFu71d6JhPy7Mq/W
U/wmUAvc2XmY9GL+HYHaHwEgKdnN3dRO4sZu12zQdBrBkbUVMvfZ2QQNsLV4JGFfj5Pd3c7jsCRY
cxS9DHDg9j0OADaensioEL+p0F2HUjyFxXpeOGmLnlA+bKFMopMgkb6d5RHk2HEvmFcrWlyvecqO
j17IE41nFm81Zm79wqj0wYLr9WVA8r2BAZ5wkUIvUz0bjvEuAuRAgYC60bIgUDQfSn1QL1PNij1M
7JV8eNjgz3Wculenks/1hW4YjqKq5AQrEzoexoSDuB57nSvuavsttMxHiAm5TuOkmjz5w882ILrX
H5Ti+d3IfP58h2+n8IPvCKqYjrpNc2v/brp+P6FcifLov+HbHXS5RFnQ13jcXw+SIUekRLD0WCMl
FksXkWybRbwQWXdD7Q9Ty+gy94VyhFEsc/sNE3j7BqfhEVrxKx1agizIdlUlbEGurdqYAIFkv6cy
wVN/TojcpYbeydO6h5/Ao3Ip2ciEaimak0dxujCVdoIxxEdXXM8LMRDuT1Zikt0YFQtFy4LEYKeq
6i4Z2fpCpvKJHbWve1asbCcZqS2Q9DrioXj0AwvTjSX1AFcy/DuimdlnpGkdyvqML5/bphEJE3K5
TYmZNhcXKtjAIGzpZakWfga/4xTyKzU92fIvLaVFeY1pFYj/02gp3vM047MEvwcrCQnrRR4XM+ZW
dyHPQh1SmQ3bo75R8QZyIJchnaYm1kwvlV4UqPq6/CA+H3PSi1KmjdSt7Yif2YRLaEKTosl0mQpf
AiCN8NS+HJw2FRLHtZnXcvf1lXgUBb5kzlt7qQARnjc1oJ3qVKIg6GuvypWDfOnBW3JaSU4lbkys
46XgaR9hdwzRGUI8VRUTmZo5/reCjGtff2J/K3n+cdDRUtnSOTEudXrkMVYm+nUJ8ksqazbSI+M/
C0LnHpackHKPm0xE2NWaG9UgUztzStl9gvXpbXaK5Ahi+AIWYF9lb49MxdSPBYkWHozC8QN4eMOx
KjCJOBSB9G5PleXEZYRFzSO5tK7yZc8b1g18sSKN7VM3HhpezwdYQELeFuz4jNih66cxfEqcSzru
HA2fhyZG+LBgnRP4FWuvVr4NcjwRryQUoF0EjHD43uhKyT0+UKaZogASSWUvSbFV4UeNrD4mvdEt
ZdOf8UnI2lE8SJ1OIb5wE5hyh8jYfMOwk9NExdMG6s7Y3o/6Yg4kGMXhQvIdie2lrHRkTr4hmfQJ
MuTHMuhjQYUEk/ME9ZWw65tEM94mxyzJl9MOaddNsJriDmqLGkXiX4t7rOEOCvtghssgvz17jrZX
kGAp8wIYdEX0AwunNCWzlrHbxRJZCeN2+r6PNXyIW+yTe054VjZmyulp0alV8+7Vur3qEzIFAH96
ttj+NtN9X6slxT/wHlrDbSwgtKcTmTk/gr1kB5FbzRzsLo+Ano374QURygZHkFxHpOh2wDjkiZC/
ZlCdIkovig3pJNyF70Nq8+ckrQIaIUpKXHFoWLxLH1lGDQDqyd9z46oOSusHSGC8tAvu2Y3tO4dc
c95wygHZBcW3Fv5I/9Ukg3gFEIGjVCWuZzKSvoLuytS3OoAPvk0h318vYQeQ47ZyubQKM2UIHL5K
xX7pmr9C69xaXNhofoTCo135QhUqiCqq6/FFsoskqkEXDjviiZY8l2257A6d9Lpmlp9F1xUWPfG8
+lLmXKKrm17cmDVYQIAkyRbWcPs0IwAtJ3MhJD+Rm/vqffsvoQCV+0ZPwAa0GsxXPfBMf2NrZrNJ
GKbBlzyjj4E7PRfqWObWLmvsjfIAnPq4C2e95+CHuWNt2bqF+3nFNWRAU/srfTsB0j4P8UAX5Dwe
DXCzjk6gL+yiMUO+hZPEvCwuxnkDWwDKt/dVPbid+wNOFWT4pQQBe4yCtbysQDeHxdWitljKAjT6
J/0dSBcs3nU/RLpk5TQu+4O/Nl38q9AYwu3PE8EkrX0i0SHdAf22myeiBYUDUpV0Tu0+0p8c871p
nc6XClk0MRqpqPIS6+05dWCaoF2n2nK11qo/6IN2lTtB5prDHhrYe8gyZO3gKV4kl8ita0q2RUz1
czkOtI07rAqZFH5v0WtZ7q+TAq7pRA4j9ttUQ85VtGIg6wIYRJ9qvFdikxnctGmFlyQXv9rcN6IT
0FRPTv/noyjbES/zi1opLkU2ywUzR5uVRYkC2Qib+1yvs6Tk2l7pNchyIzjk/4ibv5xfQWeQh6fL
0/rdPzjcRNDN9xkqtOPgQ+Rx7xGy3dcl2OX5cSNZKomdciSgnWr1udeGtiRcSjLHC1OVf3pRWFVZ
uXpUQcWpqxt8wc0S8wAZq7vVn2C4Bwjb2JHZiKsA7IXqf7f2035NErtcG4WMk1fIYYJkDwEUHbCS
VpppGlqQo7B9XZpWavpBIyMy1dPoZ4V+TvhIAKHmp0qdhl/HaskkKV2975ZNP8a0JbZkZKknclNz
SQthYaWqnP1aKnq2siu+rfPwZMqp4k4IcqXi9lj66nU0jMiS++nPFf7V3Nr8m9esanGM80920r2S
d8T4qCc0G9tGHEjHKZr1PZmj4q4uWA7RnLYPm+6cQmSQah6c4//j6gEkHXklZnxw+FtmFoQWyiJ6
LGMj1rVCKtRzdWMotCCAYBa6kWlArvbz8CBbcVHGMc6N4LMtu+Z34+a1+EG/BFJrl1Hv8BFIJH/B
WfTIaF7pgwnCfU5J/bCGQkw0EqWjNGAV5tmCrYkB5moMM6DW6oeAp0rJKxBPvNDf/UiZlPBo5jCr
Wa2+5e0TcjOn74A4+lZJLP0+YHKFi1sTLbVqYqD7MG6QPep81QCgG5BLghPmRi1mlk0hUeXpB9ot
e7nNuEBel3paik9lf+ywRpMeQAHuw5PKTGV4cRU+iOP20sUnYgJHO9aJJQagDNS8HYMuZa5t4orM
4HPETw46mnkKKTTclzWdecZqkatD1vt69yEfs9fLyo+YKbGObV2NR2v4A09a69zP2eXJwf7NcEia
EwAymuCvVaHx7WSsX6FDIIgr2sdno1+sP3C93wrKbRVsqFwWZeW0dvW/4wx3XzM6VEMn+CGzdQlx
4gI+588yHrpMMUoUtNZZ+5kbvFZox9myHuw8ENX0+L6JSd1wLVysKwKXRNGL6kGn5xyJRV7mb76n
K6eLHA9iUpyt1WAMfzE5ueUHi1Ya175xkMvYgyiVM/mTvet7ryPgWxdnKFLiMcYSgfJYJHKjj2Dd
OdIYYWtGzUe40CAnZBEKaERF1Wz9CuLJanlMgnT3oJYFcHuzka+oGmD1VfHSEfeJ5W78jSTb1cu6
rQv+7VnmWsuY9m1OEYb1tayxo2rWifbp/OJYOpoLGVRR1s9xU0QESXPlagwL1imy0lcGtUwnhyID
B3FYH/voUP+Pv7gupvntGoJF0AlnGrs+p3AUUvR/kGK/gEs+7skIkYe+0SFVj2GPGXOceIDdgfqK
Q12jrbfAQjXVDcAkfYqXPaRKrJ4rHNLe07lCb1irNjRUCiYdewAtP79APBIJHD7+bnWmZ1FJ00hs
jMILPFsGFsaMFoGjurzdsGYtcEMWNgg8ozMNngQD1ZjIXwW6Gk2P8xoLCxVMnAcyvcZIvJVs0ZDt
RVDaq8QN/JqGqUp+NIwx3yQ8yekiid3Ehq2uvC81ncdn3f25EXAvPHTFdTobcKiXxYt6Af1l1C/S
Pm2qKIrdM7N2JCRPBeS5pOLMLT5hsq8d4OQ0nkoTZukBHy84didUwK1lCMqyu0BFsi//azOxw//6
nYsBYj1QI66ptKhv50kCcjBwQOOdTFw4LdujGzaNogmQTfxvFLaanA2NKAJzqjUeoDrIRcPmiop8
HQ4k197oDo37Jwh6KMEaIYJvaBULcxgu/xZRl1t6O8lIArZUf6zdt2xzDPuJO7OS5SubgR4J6ka2
SrbilS7lROBRryYV4iEvKdoyRJw9guJtOfqhV4VB6dMLLiMttgoo291tHpzn4hjEPg4Ubmn9JvRc
fyrIDpg1UP1mvjkDjmMzokUfu3BQqGBHSzdxLUzWrYtipvadWRbd3Z+uhTFNPFk7qnclFzaIM6hV
RmVtLOqqNNRH6BZ5beUCMMsGG4IBE9AZUT9NDFudPi3GLg7A1dpOCN/kh+q3JFkl6eUPtNXJd56r
2KUzsxvilCjA3lvhXAlTyf4bt40unF/38BcZKaETBaO0Kf/NpxGIGbtOjGxIq7DZ7l0FLRFVFtdH
8Z2mY8Pveeho4PmCB19xCt9u7JKOtOgEMSttqUB4vXj75vGmftbILUuVhbH9/T1cJbqNqFty7+FT
cFhW1JKcWV1Qghzaibc7cgo25uf8LSnymHB9Tippobvbk09kFF5avUZu5APgJ5L8xF+C7gaG53V/
Bk+z2NQmP8Xe3tATmOJr55YMOC+Woepnz/WC/R/VJODT1BDktW+Yve2pF1Z+nwMRvP+A8dz8QHGJ
WetlUwhE/YX9CGY+F58BucLmJKouvoGX+FnHIOQLF0ITzzCE6Q6xaR5q3g4Eae3eFQSqKKi6JuGC
K7hZQIoGwfk8bqEZAtL4ZtbeabhNyfT2BQ0xJh8gfZnHtNxlYsKkeBC992i4voZ0RVPVblDuRBoD
RzlKo9MYtdvciM6WK4A3OYbAymOJl/eLmQpRgeHVVuONC0aQioKpAkwP5hKlKhxOiDY7joyp1G9Q
vK20ofyaGY2uvfW1C2c/7RPCjEjKzJzMOPFTFEz3Yn1mITdrzQcCoQFhUsPAaim4KnkkmAfflXGP
i7QVpTRNo46+uvkQZHYIqV2QHIa5kJUXZUTgLwbRuhbfZuKNeLtcXN0/4t/msuPnh1ekofzLsF/N
LJ4U3zrT++H+t3nZ+uuHCHAye6Z9n2kRYNUgH2hytvom/KzvNlWahQhRfl1EasG84SzAqHyJTy9I
iQLibSI7nrl8gPeZIgbiANhiB4XBgsWDL4kblluSIgjfbVdKkgtInnkva38TrVNy42y3uGqcDUlQ
RTRvWCB9U/BkS4bSm5vSp/WraIhHJtyGzGSaz1WG/K8iOL4VcWrKWFCBnjQbTcH3lRx2PX3Hw0t0
yXxd0UadPFWEwlwo+z0FWcGs1X8Ivi6JvQ6VOwwJ7hzydthQfcf6QUsAGWvymj/G+6vxM15nTEgi
WiSdA/bQRhFi9+3f73qASQ2+Z8E2pomJsqKf8dWPqYEhbfIowQb1hmrSbohJrScld58nF3cGm0dn
P7hHEy+IRg+ZcuedJ3dAubB+f0rLfSPVuRNqJKH9M4IdSN+HWP4dB0eLCKZQinbB11Om2HXPhAg0
O1eTNtZkGGNCJiucKVVhkqU2EYw2gRXCaONXB41DGoh58QoqHWkPmIdbRaxk9dvlL9y2KA35+jUW
spzH3YKpymaoRrPfAB+MTyHKtUaLsEuSqdD6rZujI/89cNk8D6yI27UoNBO2tywq69jZ9MRyDn2u
RhHN9SZtMDWEtyICvh+ple7sjYTFsZak8CIXo/79/Ia+Jo1CqYfTJT5szHHkQcdo3/4DRkJTzTOr
ROVs/sa/SCKJDVIM6ZQkdRDmIkGPJn/Opyc/jwG4pUF4VMLq8CeqfsyuX2SQQkprAal9urAIQv9l
2wmXdKNxdo0n1oWdXtYElhaYlHXbt9ZDKhTzuiCuHjYmAMEHOTwqnSltwRWFnKLDbmUEM9sg+UCs
Uy64hNmhBwrmf1W+gPkjtKvfMmC4gg8+1G7TM7fO4R4tOFJG3qt4UGGnPzx3HtXBzzdjX6grqMgU
GQkfisMKYIJlBixC2QrNA+Ehh73PIcAX3ZrrXOYKp/uzImdx9T3sHXc0aBXYpRe71DwV0QEsqMft
iuSZ42IT4Xp+IfEzS85g/6M6hsOBto2WaHJ5oCWp2cxgQIFGL2Z0VJrunVXqwpOvwxAm6Jqt+QFT
olCqmcVlIDxeNAYfVH4NYtveeNX217uYucD6qpmKlkXdI4IB4QoFSN+rIOKksCo/quxgfrLt+NSk
F6ZumvgQXNTfa/SIEMKq96kHvHqEb5VfCSbWkzmcsHRksmc7p1Ir38GB+3ykbzcfrKLkCsonH8n2
YdI6x3urfGvb36xy/l6zxaE48tfKLOdjKtyZSjJmyRjC24AufZfCudY0jFPxJH6+CKlTkiMr/gsE
HKfQHlRiRxe2XLmQiKctE3s6CY/CooBamg8og92G9WUGOaAKzFcWScrdw6MxM0EGO37s28TngRJ8
PNPcwHvsfaUrvx3P3GQ937nOsvTzQ9U15bFgQgAX1yFTxiraFEk/egkcWwWiUDilZz7TZ6BmRGC8
yxCmUE4lsmp5EpCtWtjwg1GMozM3TJKC/TrqBxUnzTTlntJOpTwCm2C5iq9qRa9F5aWpURJp48zd
mPGFlx6uVn76wAjenVxM54WnNb5PmGKfw7lfZpXzkHvnewB80gqGPxOlS/Nx2mKIInCsdLYFuzjz
RqzU8grOgOYdzn1zhAGI2htUuYNzcOlqmby7Dtu7zr4BlvHkluJ3TE2USLlMyvHpIYEwmwqfDLKd
cFXRjfQm60FDj3+eeu/AOuWCUuOXcmrpLMawLE9ejxHKQkm2kfKxNjvP9H/FOPrOLhZ9l0n659VA
orNfz2pyizGaRABLem9HJ5XpkWqh0rMs2ONwGi8tXIL/7oqq4ThjUDqYeg/y2DKQ0a9jzrMNZ3TH
4xrmspItaWFDwd5tZg2NLqDzy1rWqNw4SwvN/swJUOBtVvUz5eyr7Le7D3/E32CNFpUTwOjiolQc
R3bNyeDSRZpZlw+CK/I/Jbtba8RUsMu5adteaRqgrlovgztSA54N2y7Ns+wHBfzP0R7PJeGMyukO
tbPpdK0SUqylmoFa2KhBqHjy8wO6EwdOBwFJ0L9PfPe/BmwwmkRkJEb5mnSj3DJrUWjck/QGiWF5
vr05R/6QMI0fl90nzHq5xCISw4KU0/KUam1DInf75SehEpec8049c13ju3CSMikwGGBRGVp6Hiyi
r3nrPA+eL8hs/qebdxHJ56CMFKRHlJ39zKA+8TUuXFu06DdQYx3pa4De3NGXrgdP/Ci7XYb9DzIF
6V0zNsoqbKhayK65vE1mNYaeDzVqp5QYEE4MP15DTxs5jQZrGskYvFgKC4nFVix8qzV0XN5dBC37
yYaKdlYWUAdqpljJgnwqEPH4DqRXJ0yn9d1nEI8ZrJy41wx2Ai5Lfzj6JIVZgFa6WqY95OhO798o
sgFI4G8zWlaDHSa2nSqQhXJoi2PIE0VRk1p75efZT2oVQXc3TwnEVxIAYOmxxaQmoiHpih7vOzSa
KG1bG3WtTMepqe9yzYmtT04tDnSl28/3nmH5SzpHEFEAUQIRRIZnv6iaPgqzDeNKgddKmcBuB84l
x3UQF3NXSr9HaHxUYpow453aThdAOLCNPyAkGqjHOqUiSaIr5TPZ2a4ZJI4iZzhcMVvAlA43kxVR
tpxsaDnUlkGEBAS2PH9R9EET1MJ3PjMJ93Se7XtsLlAiUFNryFJfKOeeZZ9O+nRUzrlZUf9dHEy6
Ihx4jTnt5rJbranN6UFlPV5o+pYcKIGC5RzjOw1lLD+82UPIgo6F8munH+IdrCC7UeMAVspgCBMG
6858Y1KMx3O+Br21iMrU9PV0oC3CXTGNZ+zx+fYRxYa+h7rJJsqyAm1yEPfQhRMo5JUtsOqLylRL
5mi3x+UxALTCaFfxsFWEdqxeVmdYbUxAV3GFPdicc+Yoc5ZE7JRTs807H6KTinlqhQB/QksZR3Ub
GT9ZiAj6VNQ3bu/L46KrEJeyz1vOonc7kVpAcF2hkC05AslWFCCA0tKJrJ0X1L+o7QJbd05IiR3A
tJd311UpY5lTrQRp6Y2Ai7/R51Wg30G7SMwBSi7ajtyZ4hInSsesLr9sHuXDhKpjiMqs1nsjZJ2T
CVAg45LcqDfNErgpj78IvSsZ4W/wfOIsAMhETt5eh2apr2YtahG14lS1V72Kltsi7nx+4Uwlta5z
kt01ywMdUWzt3jbLgZb6tRSjgXAmHYC9k2Tc45m9MW9/BLMPXO113aO3bG9Ex7UgOFUvAhX6rdAm
RDvTX5jGs1VANKiMSKa1+WlJ3+biKTqMMPydookd9jSjEr4Uu60OxRkU53yLcq9+yjQIp78n+Ksr
oDhur35Y/0MOOjAduAAg7LiagpRUzI4ULHrScXHWZRKgx3EAZIdLZql9W0At+5gmw2Nn/7cIaZLr
ya/iYD7HhP6Jd4H1fC7wBiKdQv8UD9rxPGiZCZrLgX0lGeEw8Efuhb0noojmpQI0AsHA4aSmrfxI
GAUT46ve0eQHQh15sdGvUzV2xd6bkHgAuwv/fkxcwpp9+32s7iFBVVadCjm3ADRUTJcIHxWxDKdc
DNOOTAowmF1nvRWYWJubh9jJGZnscXr5PHLVPRX4CCi0qZksEeyjs0bWrMm2bOEt8877aB9ZFUF5
D0MW0790DEt10JMnMzQoCmHAkwtE7V2PxTgHSs7wqNkD+c58nhyEsNMdvzw9sR31b2S3FnRH5x4K
+vcBbe8wBkyUtnKbi1CIZK2l0aQnFzeGXQeM5tfZz4lvwAUjPtfsXBzqxEknrPA/ATDzIxtI4orW
hAin4Pok63aYLEkYJP629QflVxHrm8g+LFtpM0b/kTNfqYHA5yFdCUppsi7OtDnYFBeej+Q+Hk58
S26c1Lq36qC0vUdcZYUswX8SUyO1ydMoLCzLd9Eg5b7Ga3QppbcnQnCRz1ErJPdqg1Ll0bF2JzGj
b6Av2TnBXJl9teriGk1pKwZxDR2UZXLWFy1ohqQaBQrtknOX3RvuAXG1MthWHs77kkRt51+DaYNV
EQH5ZsVsjgWwKQ9ymWkD91JDY6qRGG32CoiZawi7VexOSBC1GKKyP1KXgYQFhfY6/e7G49FIgHwi
nkM2cAMeNLZGfnKMSBcgdlrDbyxREowNYWautGSFWDiecVZ+sVdE/okIFEDWjXBzZWe/j1E3Zmpv
kq4mnYDlldM7kGw/IGEq+WxOyNBUBfgM768syZhf4Vzuub8okGiKzOQr07hqzyE9hxcPBU2HMnqI
9lPntjAjc7nbQBCudADFbw+1qzfEhaCK1JzCoilNnmC1nQ6cIvK9qOaAm3PXYiDeFvxWODrBy1nE
LALBKt2CzHK23KNKm7vEOnxl96eYr25xurtHr08YoPZfSUXaZF/ZJGwsR3X5tOG4/oC4ZBV9ms93
+JZY+SRBcPiOExkzHC/WMxAV/19lXyU/ysERKc9yCmngLdBTzUqAnmc82Q4G32z0ezXElu75yt0A
sz0C4JAYluu4dZDQx2imxUtLSdcoP2mZBpV8QVYoqfGY9dg1RktcLkQ9NBQH+WAYKIoHuQ6KQWTI
4Eal/ACB1bK8z3MEFjhcRx3l8zi3FYc0lyajyRB4yaSTH2rTf0PSY+pBvD6vCn0H5/jo1anhHPLR
McuI0LKo1LGCrbCK/h7u52qa0xhPkyJu6ZB6RS/zQuObDFcwslATu6EVtFkzcSU09fTlmMKV9cK7
Pb+AYinb6/qkzc8QBH1aoo1SKv2rcfE3COjaXZcPwXrZMGuEakQEyZ6QLP7+HvdptvGfVmF7a/MZ
TrdKwWtaiCKhCcLDkBKNA55YQlmOlqT4F7ivuc//y+gvNd7wjKDGkGUrbjw1cntbf93kSwTlYsdT
diE4AYIr7O8kz+kxTx0YkS958XLIZtEK8oDtXqNtVVbRBjGnrvTv0SW0iOTkUUV5SK+jNi67g94R
AJcBeo3P0cYmlpQMUmMVr48fNz1mFNF5AyzbuYawMMJKPacKX/5QDGLEDCGf/pOalg7N30cSxegS
2Jo+siOnMB+oiuNH/sbTi8aEACNZn1wERYGEyzTUbrQNMiNX30ehdrVCmhRA/XIWqHMeggQy6Ah3
uYjBCzedvSikzQs8uB3JT9uwKSUt/z+ROwEnLlOEp+KFXvBh2uj41qkH7A71KvJOAi4UbYWURNJC
JbOR8rJXk2+97J5JbM3mPSThZl3B91he0pRZASfB/c9dgZrZhCkBcXpOcrrV371NNixifB5ZrL3m
gASBWeW2DheyV7iyo9/RaVLOJp61MIcqK4JCLq4mpYP2GPaif7H9ReEMpdC0CxLTBz5K+zu2IDRJ
Tp9/o8TBdcoYqg2qF7wI6iZSqSzk01fVRmy5bKEsQyx7uZRy8H6aTH5jtoUZ+t7Te6qpzG2SexZu
tEQ42FlWvxTfIdDfxd9OAgfEDdk76/bBG0TreljHJmCEiWZ7G0snDQOrWbVtVjuXGICHPRqjNe5G
3LU2UNAZGa3+DDMF0CTx4YKhnwh1qU2VS9FVvtEK81fXsV2Z/3zJuaKp0th21LjCrk21VWhY3Ejb
0NX/Bs09CSOU3Y85KbooRLrKBc3aW5ZSzXnPKlRPi6Me8GeZQs2vuvs2+IqSt4GHwvUPbzqU7FHt
mrOh7EoN+N8AUsxaAiWZeSgurcCap97Sd3eoyQUkfv9M803tE2xCWrFVVwSaPlR8/0rzMcVdDASZ
ts4C9J9O4FEnFH3SVEggg0fNbHYz79jj2GNV1arqc6nvWeQ52fCNQTJg7EYBzefn7J2lkhVGSYzX
RCAOKgivYCTpHfZPuNtv0ZF5iSDfuyuG8CjDiCg3rB6dCbTtpTUMmLlTQ01NNW+deFKTbsJGwC7y
lUsjaSyhsji3ShPjJsnJ+q3n3suD9fT3/nsadTJYbMoj7uaisjiBOM5FXNcvHIfxour8avkyFy73
F5HjW80BwfzrkU0pY93XzCKPvzC1y3NAiYksoU5L/MCFPsDkoto6pkngi7CuspsV6G92uCYLNQFU
d5YSdiVgUZ6WnkgDDimq4brXecqf15MKnnPagrVB26ZEEppcEkqmQna5Q7/iDEjp9J3pF+qLT2+O
NYFdqBQem3UaYl6bcugdThExWMFis8yi+gvM6TI4UWy2DPE/b1x6z3m7s2HIKHbFfnGuSojEhAi6
cqEXTAKMyRfhRXa+Ua1dtnDNroNT7PV/e9Zam9PZZfFo0vYwPQXvO4IzHwlwJlfposb+dnAPLb7s
OD/GLrWUQiD+6xrerCo0q7f50wACQfmkDfVmXb0VUFyzFfcsja5YOsEp6mR9oKu6wQBd3QmeA6jP
km+fuH34ISqDXeU8a402eqBaKIP+EA0D4D4oCwQWeKx504CPOoCXsRc6NGpUilHm5fpGh0iZ816b
gP/JdF/Z34Wxi+05oEta3XyoPnimMSgeBzMvDV2RX0EgpM3ynqCsSqT/mgx3lLFyaCk3iDtOJ7VC
TSfwHPKqsRyWQ7UHeKet3FGJJTorb2K8mkarx6LDN/+zeX/KJyC7VMR+FIlherwuYG8+He2b6Ihh
nMc6k3WpU341Y0WCFgQdz1hj7TawK36oti0216Fy0WFUnpKmeDqW9/LP384Gpss/Ko5DVQ2TPLca
dJSGiDskJ6xanezuyQCMhB6tVVBHnrSmkK7lwLOsdGvndgA1SzWHwZ+rTl4JfGBrGFgjyasqu2Mk
boSEk6nRHqpvRSOtdnNlqjdLIhU2J5v2CBkZ+e8+00nlMfu7Q+E01BDZja9jI7I5AQfD+oInfSjd
eKYXdkVLDAjp8UrIn7IM7Rk3iQDo8585Y8K3wA5vfZk9cM9oNRdlY7qLsqmC0O2THUO1nEFv8pm0
sDnefEXILMquybgc06IOZSPN0DGDtzfKwsz/Cp34niL5ERWd9JIcjd17Ai1L/TJJBGU+FiJzZIq3
vVKxP9MNlFSUVrZEci+UiysIZk9fDvVZ0zR3w1SP1zclauLMhToYOVbCYDi773DeEVUVR+s1uMr7
2BRdtrTiC+74fFqtkridEjSdbBmQeAq8Zcl5Rp9jxoZb/7cwa+CQvzOL69iN/rdaghAEL7zoZNMO
HqFWWgQnyEgfWil6uNkCgaq6HcpO375e63J0F+pwADGYwtO12l9AlR/9PtB8vaBfM0DFI/iCm+lm
0NJJinonRr336ilafbtoLvzh1W+B+s1LE2cbbdZkVe/GvMHEKwCfX/uJ99sqiI+LXoPEODe731tp
bSkTwAvee1mA8Z2GdLjkMgOYOtROU9EftMxzCabMVP+twFXe1Xjt8fucuiEPNf4FUfDsVb5y6Lcs
A5wooRLT48+Kxz9DvEvi2O7H4um8UIJ0aBvxKRWfWB7K2rkmJroVIx8t8NND8iqVrmNRrw2CkXLF
V0emdZGc91SvYlRf99EWyPxhUNLEak8FLW99k3qnULbxbMbCxn7orZWFYm3LufHZ0p8U+xtDZIIa
UQ2wLodwzx/fulmyYobDjcWQub1RYelM7j+LXbPSxs0I3coAGzwupBzaanobSaV23JAFh2VeTFNw
1J/8DorJMtCkPJ991IL+BdAEQc27fNhY5mPuEd1VSzjrKizOs6+RTsGyr7VAxOuGKG66ZIK4+1cQ
SjNAAliAP+ZvWdB1fnxOGsFyfM/5JwSEnL8XfiV2KWf9jyFhLXNopDqcBrfACYr0XAyOiWLwUutb
DJ+TXFqDi5Bgtue78ruUOXlE5qLUON3lszHEhVlbN2tkyxPOJb/CQLPr5robsHoZa8gHM4gFRZwN
W893hGJuYgCiERkcgJRuhxWp8QrA6d4OQ1USZRBRwe3t5bKqI1HnEbKMF7xPOcRnmxq/TST+6LOJ
s88i+MtbSo0J0ODue2CUbR3EbddBB+HmP83DqLyc9tBs9UzyKcHD5GTvg242oeowQoJ9n9Vhb1Yp
tiD8frsLP8E4CQF9Wt0bPVNO5/EJlbeWZkbNopvaunbdIA+Gqpv8I8uDoaGlB+o+EGIDLdk8WW8C
Auyox/+LJJ2+9hQjuLJs3j/Fdq52EbUPURaP8dcpfds0wZKMebI8odcKtyHXyVTi4teHXK6MWb8k
yhnl1Wwk4Qx7PdnYHf5c66w9eFjSdJGQ+U2yJIu4jiyCGBXcBF7H49rcvCuJyvJTJSbkIRhyDxh8
450wXgCNcYCuWWEtAUEouiurqWy3UnRoo0EMgWsZClCuYQ/vrUwxAe4I1ffV+ugia3lh9Gaw5mSl
DmFZDZCTBHEFYOHSTk+/nVP2Ib5luiym4V4xd7IJLgYaZNf6GBQIAsrM7icBTtOB6zJ2sCAQI36s
WIaCveHts7+KIEes+4BcF+hxV4TkZk00TCfJBgCu7fd0PRnXv/55XlV5NOqh44DatoKOVI4QBfKQ
IndbERIVH/loJZeeOet3jasSORbCvpTtJ6HtnrzWDZEZ3/87bh7P0MdIVg9umvg/uy0l2fRLDNqi
Z8LYIRXk06KrI3xhlq8Fl9esoKzFanpIAdw7H/iLyQudtmcN9plDheBBeZxOGimThVydLyDtZMqk
af2StzS3xg6XGR7Q6d/p4rcOb2n5XZSYaZAMTUk8NZu84oROzrLRBiyDODrJTLGqTFt3yTjcKAuM
XAiIrCnS/y8tZ9oQWvbQJSN0zbvDe4IDOaM/NIVzAuMq2+t3yGiDgHK5xpJRj7fG4nfioOWwJpam
InHJFw0qTNzCNSjfM5/VDseQWk9mGJnFsIaMIidavKrse4EWQazINvhP7UoJ3U3Oqv5qy+vIK9dD
ES8KalGH36m+vyC4s7K2cKjDfpWwJB9qT0zABX8COjXpNnQ9GVLq9ja7ykkAKDWrTze+OWQc+Iq3
imqzI9shGCelYzK7CgHpkih1gYAtUKDi9Ao/0tfmW+IAvseGL2y9cP7fBGQpezQgZl3MGjv3k8Ky
IviW8h1twb/IB/pWkU1Nnib1zc6TnLw5SM3F0nsL9fD9mZOt0PaOPPBOlptB9Cpc2BhQOF1PRyJs
XCAm2hrQQgHU0mKWuqvi7qtCixMiB3wzznwjeP2LODxdnG6Q7iUebtGxYsg1ezDj5wrzqmR4z+/1
jrwHEJ+XpYvAgT4FQoEHF6LdcM6/RSdSQ6Ah5+zgrLLJ77QT8eCB8XOiunt4gVja7BsVBhwS3v+7
4izxr4ogOmTOo9xmQvLMrbNRGVm/LJlo2CiMm3w5DH+UFTVluZUen2jknltgDMRYgYKf7Nolizxn
303MqhwpIFMqAdtSFKK88Nhq+rhdR1AYucg3RH+zhm8QOwgVXUeqJnVJbAuvmaRT+T4Rbj1p9OD1
EEaLx64jTH3dHSJGWUBKRNvdLa3QCgilXHiHgvSzlcx1Z88PxBQ+prZDOd0hMZGKT7KBaubuS3Ps
Y5HnZUnY7XcTebh1rRRRqpdunyw06X9d9eIDGRXLyHY7rtueiYCewEviWbSz/Q5e8JbfhL1YK56h
6tfAez1i/7Zs0sg8flHaqvihqatFUA2TUBKe/oHSygYt/Rb5fa98PlK8XLP9QWsn5tfbjgdAItQb
WqFV1FszGflPBJLPnSTV64G3VEUe6uP0RsMijTFrFr+ZVB1j/LaNXFYwiFdQmMer66+bkxsxKVyG
8whLGcgQLXxUcAy8PXPCQXSXSEbhLQqtMNL1d9C6V40ugdrCO2mK0mp8JvdWKPTBjZAON2WUBnae
5PduSvRILBPyqEOf8btCtAVdV8NEwTmikLVp7w8HCCRawVHgUuOcOtEi9a0RQeheSNG4qOcCLLL+
KthJeflDX1HpnPgn5AK7S+U9ORLoQst0xZK88KvCMNjq4qQofQml9E+wgOjwk0AHSaQtVLSxFqSx
fFw0G/7eCnpel2KbowjgE5/GwRldAPn+trOiEUJX9CpbPkUaaywHUabRDwSMJUazqH5m9t0JBpU2
E6xVp78X4rDWlZOn+g5myebxEhALWN8xG+Q2dEkajLNDijFye/SMkmBBZ3IPz5Y3ZzFRw3FhfEgb
+HKgva0P7Nn9rvxhCTzXm3XA8/45ZW491z4ghrjWDz0w2EtVZy0yBnpkub2mXxrypHSiojGw3Wah
vSrX3Xu5C9ND7f7O0QJdAk1hXhhDzqirZbeY7I2/X+0L/TL8K3aRrJnQ5RX8xntEMFH3/dVxpnDZ
7tk60pjyloK2PKzNZV+lL0ZHDYx31DvTtxJNM6EDZO+6rt29ONle2fLAUiu3I09IWpPb4dT0E2XZ
5ReT8gzjTvR0uXgW7EN3RrO+lR4oGjPMGsBVOPhYgLzKpDFoWhIYvOc7IvjWifpqj8JaQelybp8n
KPbfXphwXdZeyqyozAGE1R996vkgtZ3zGW84BZYIxyMiaDo6oyBafhVjAsBtIhqBWmmE+qCHscPK
CIfMX/ytXxo+wumKh1gxkerI/ZY8k6ZdjlPnx+RhjE38mdmhFxrTuA3aHooGi/p95Jj8AKtyDKom
nUUtv/H5kHglyGID/HiMYi4BZT6Pzy8v7+wjO4dGyeZCW6sL4/PodO64lyE7bOsuA/N45HVROd6T
p13H0gT8JrbWo8eV0rZEFfKKNTA5/eAgNZIuX0cLXJdNSe8Bg1T1eLlwlli8VLFajRUIHefeoYDO
sjuzZ4cnVBZOklNjG6nR2XCPUnl2/Mgw1d76wQUmDcNONvImoXi7Uxv971Pa/nHdaqYWCynZKkge
PQy1JoX0VeumiNDBHV4gYT/yEwX5sspUDKw0Ah7tlvEaDT8GIPTBbea4ZAdQ5wM1ixbU1oHq4bwQ
eej6lUb3eIbkiMFFIrq2RrK9YGw2Toh6+8HuUFK7sBhyZDbj8m6rY+1ri5dQKgQOmYw9xcJbmCH2
ttGiW1eDGpzudtz00ZXXKIU8k0VpXFTgS/AM+QYrecZP35S9NHze6dKLDlQ1ugWndQo9MofXl6K/
yHvhg00ZTdDNr9jtKhVK4LX64U8XjS/KSdBIKbY8HOLxfvT5YXQ3x1cuwsbAoheBfCd2TOAE2pss
Iz+Bc3I7rz9Su/LYZ5uBah+gcOwqpRmmSFsAkRbJ0OZpTyM0dciUisafQV/fbtV+Zk8ATY7RHw8L
WgV6S8/jS6vKesjpYZZOWJVOuWO8J7srAweQ4SWQyLPAmpYn0bBzz+Iu6hxLio7b6WswrsJOpLaW
2Tp6Xvb3xHQlIBSdOM720sQfsjYS94gB3UNYLTtKS+xmQYFnPiZZXR1YXwlP0cYefZUvbkQtzVg4
G/GvZ6EBrMfeT6oWav2AITezhfj7ANKZlU26Sz3s7GF0MIkDrNBs19h5jUnv3Hfeo6Hnz2Vvc94p
82BXm/9YHRgDYrxNze1GWQyWx8V8iFxPSXufF0M+tR8uZHf11nkXlgbQv1XtyFpfoWpXZHFqSHdm
ZxHmZ3oJKVEk4IwDeZlGcXmkweT0M0fjmS5GNvcaaxpYoGDNvWkTacPJq7tEsHZ6vkcmOpgeeD7b
v4cITGndXxMymos5aF2qgTsKZUfBWbToVMccVM2W2iz51bcEeSVH5vIhtPGClx/NeNE0D/ZoKDxO
RquTtIqux/6MiOxVcsemJD9pr8LdAtwvZmQUyLSNGyYxKExyWq7mdM7aB3xUdg7OQi7bQsq53/wb
UdBgUe7xIkM6evqimEHF3xl6wmVu9zB2tsI7DnqJ9G+eO8V/UoSLxYYRbJtrHc3NDvjcs3LbGVZl
GgC3vdhUMXYBlBGRXyVTgDvVrF8FMcQlRPtVp4phKJC98VcAYmZ+ympTfzVlXY6dj6CGYzY5L9Nj
1CePSqmO4z8uQKicyYI4RAjB9FzWLR9xfnv2nXHUAwIsB1oERgo2Krra+U80Qxv9DWmQKvTPC203
WKgr+Jf06GM83lxwKpRGEomdvYT8a6czPKmtaFEA9YhL2hLPxG1or4zD/aEIaON88RcqAVUPtnE1
gNp2O2xeCk4sEXyN/DAnkpT8PZv59GVByZygXnsCUN4IzWrUSoHTGI6b4OCl9muR9wmRm2svKJta
PPyZHMzYm4Ncmosz44TaVrPLdVgwbJceD2SaRyJ4uiQ9JJNrSYMcBLncC6/rl9rDn/K0Y9kCmmd4
iaJazQWgrW24WpLX/kp0zD/4BNdDQdSZ+rt4VdGHh4aSEL0Mg51s7Il+dr6DT8kfh+djy8oX/QLr
0+wT0brbDW3OompO/BfAH3lG1ikkQ3QJubJ9Gd+6mNETtCN9kBSGYV+6VfVzqzRUnzdro1EL78K8
nNbcVgplhZdZPwbzZHl/8hY07qcV6k/kMZsZn0nfx2sHwOeOapZMCOfVK8CxO/mo6TV6h+DMBUt+
HhtegbQvWXJd2givKLKjMwCkeDs6PjoOhuoZvfTXMXyGWxNov61ovtod9IhkMF+KNGgChIZR5zKQ
F0hh7otICXnyIu02Ukx48VX2PoqY11wd1GIgqrjBNMd9MmKvmUSScI4IDfJvzonL+4TIfcKNuKmJ
g6Mmg/cV8KvpKP2k/lKd8/oC1pVP2ba1mDl5s0vmbtX0Bycbhr2Z+cAIzw1gyvsb0IU/VIfa/+zf
yGb8q07yPh9wpYrQPlrM829HWj6j9teq9zPya1JKVMAl9oxjItrnYZcJfFl4FynN4RUWq6HppA7r
X69GRJKRVtEV6sJRGYcvqnHpDDA/PKOUCoqmAkJGcTgTp/MlUu848j621e/f2+/Fhji7Lb6btHel
Alb/B0JNERxLwALpuHGToiFlc8s2WoNkMpZk4kVIOrh+kokMpjfdWGQWgC38WZY7PsrRpuLPgbwI
04Du+kYqh/d96r2NzTrNQmARkvo3UPpnge3VrFGvp4j6bzkcJmV76VExpV5ZhBBUx6sZ1ehQILDx
qTmXzwa52PJxTYIw+uL4jT2OQ/MNP+QqlEP+dDv3Y+pHCYOZKGQaYOiHPbbtVhVy2bKEoSGnGRNp
xUpAh4SkZXW+cCiAGX05bCRDBdEw0d/5dvsHmfSuTgq4LWBC1jRLGxaDsfayP4i0HDs5CZA/qwsO
69o/+AxiILxbE+C3TjdK32tPcdrO1waN9Wyx4KNbaZxqQUfNJHo6BGyhnB27Rk7rmwz8L2CpRMpy
VblZ9HpKbrxkIYTFbaRRqkIPqaKN6nZGIn0S/OUrJr3va3r/zQVBORhoklHkq1GKFv48A7E81Azh
cV1cVAbcf3brJ6gNjuN6WEsPt6HEkJmjp2aiPJfyrySdH05zcttfdjYr0qbwfQAvCMKRMdvu5x09
MP7o8BYNeaobT85TvSVbpY/9WZY1WKmwvVaUIHEzplk75FdsEkzKdN+ygnMpZm26EeuBWLzCgp/J
zIK4aYO9/XoADBBRf08oFaj/yPXFqCDuUhTDUyish5tCl5cCiXjr53IUfsmk9wu65mN502RT6BSD
qFGwE8f+Bvdep0wr/QvKB6L0xEUYDxsDdVER64QkcTH4P7yo5kgBaUYHQdpb1av1IhH9aO9Qv0zn
I028rMIWvy2j/M5V8JG3/JunivZkjmCPkKIwW9VR5sTtQKgi6I7M4sNF0FVR98/JhNSCCme9JqKp
m5WOXeKs0ElVhZvrOZCCRBIWuiHRdbHUsvf5eBynxCzBX/chWZWsm3mymQKxcIj2Kl1ZIrshH2OP
cbwRO5ZrQeSrOZK4fw2t3R92yBGhSnzIhZrOGAyMlcXPNZRYaAkPX/0kudMs/EK4F5kERhTq8UH6
TCIPfmw53Aqs2/Z4Y/YP64qzuzHbOwpnKKthOx9qfxql8W10sl03UxPulUm/5xQcGHhkxvVRBsK/
x3K6IRoK2hFVIMqwB2iDE9XKTksVdNr41roL/tAd1Xd8bofubQvEMfoAat+92a4ZHMTqqcynrqzG
YPQ9D56x2gGSfh33NjWR0ZxAPfps7z4TqayrZXL7G60i4mohfOjwwLjRw/XkEraX7wfmrtALVVYV
FO0cvSY6GiQPTgw3CB/wL9oq79o96pcTdjsU/rzfMbRDuViFEIqi0OrfwvpGrQnyOIks6oF22zx9
sniKDy9Oalz0CHXMcnzpvkCYuPAr+hR7pyiqBWEN6w1Rbbnw4IAHaeZWcPW/GecZXai00JGwMQUZ
rdjB9FI12aC72J6cIxNQcetV0EVLZL8XgpV37ViFxgEfIh4WnKA4yOR/YFQoUDn2bfPGQRBohCoi
OKmFpqAzGBJHH9xtD+qbXWUuqXoq1aEMK5HPP3Csve7cZ97+1fjo/QB35rx+orwWppSfKQQ4aHYV
upCM8DPPP5LNRMMLSrm3JtjkhlpnNIIl2e6mZdGhPhML6nMf4BPa9aexDbWNPrMRFAVqDKqXw3ON
9Gj0u6QTPzURHu/cC/1T0WUh8OdOXjhw7F+Vjzf4q7X+BqAEFxg+S+/FRhJ/S/yOv5gTPMTyvc+i
xkSMujglQpcxEyqiUkowzNGWWBxmcEvplJCY6HIhmMTo1TQtR71ihAUrPSULialuYCfacag3bJ51
sbud/M0vP2t2/3uvSnwm9sqBjzP7taDhJXYOSl1FWCxYouCHF2WRWEW89il7x4pCZr2Pu7SSmn0i
S9sTP20cvYsFDYXOOF1EUGDvv1k8FMV5AFKm6gRuiygvBiIyoqGFZ26PjXToaGncFoj+i0EKBmHv
YUu2/SHB+kATIMXaGN+EvzlVYvRFZc3MG55KtAipkJDw6jh/t1HdNA0cLHMaXgcRZ2vBmIoDCExy
eAyfLJN009B3cV9EVPKBoPexkdzuqlzIyLcT4EIPrBlslTyJFSf0yj2UlSLHFtbTxvDtwqQ+UcEZ
BYtPVBkapIRhqrF4OzCxMgku1URTM8mEVjh5v1rflKsBylzJpkFMRvkpZcjyCTVAP2/TyX4iKOd2
BRlXRBLLutBhxReMBDsYQ9U2lUflgGbwKJeuShLCeg37avIvydIXRLmK+wWgnzNwJa4pVgj6nV/B
7BPebmWa2ldTrBqgqBR3jdMX1/o6xxLt4rT9hLs86FsbrGBgVg0wZMgA+AbbFyPyrs5UTa3vPGbS
CHcoLzw+V674BAfo9ZrqnqKRttNQHJKxteqPfbvc1BiL9PFIzNW8U68Q74GarKFVqU3JSvJkEz2c
+wH1wc79jyIpvILKoFt5qFpPHn2AFKXa4Vw73JjfOmkUZG3WEnY2Q8BeGN8DJOsed5K6P4X78MQL
RhOz9IhZj2uK+lPi2eHoabkE/ixM5NYmOCobzCvyXkZBH+eRB6nkCMRomnhXlp+eDAN96zKbzUFh
C8C4gUIsm+cgdTmVM80oU2f48U74/ZvKuCbuyyCfPe2iA8skhlrKhLo3W3f+yQSqDlIp0RhU6h8Z
GlJxOO75AvGogFjQr/M2X9xzk3UxihI4BWfFP7Vq1CLncGgaASlNB0jK0PlCzHXv9oa3Ov/fke/V
kYJvjZ+OPeA/7IyXgg6sz8A8fh3W1yMukPR/il0Q8G9J921ZycnxLP3qypXXOgs1hou92eHHSXd+
0LILBlxsRa2jnWgV3lusdWZjXOEvE/sxo4rIiIdZ70WNHP1gPd2RkGAKvvXq97e2EvRSIbfhQBGR
U6tHQpF7Z9orJ9TlnVcy9l9OVXvXFUf60rcap60LOCWoApyPzhmmK2D7x/p+CEg5+AKFTheg5/g+
qoH2stTpzG+sfebjIsVkJubxWOIibEmGG5pHcZe+7YAWJsAkqAMU8v63jNfw0XRyn0x0xOpElABb
B1MwBBZRIvNhrukPgsAAxwZ03SsrMT2cbc9FSbGKbxdAI/1/uW3huI0xGxTH1NYItv5vPMgGGEA8
OUwUAPXGN8WoayNmTmIlqZjX9JwUmN4927It7PeLZV8ZQgidbdbMlLjgpsoHC2DwY2H9GRhlAh7v
CZaAncWU8rMuJgiG8wejBsTmIfi0EnioyxN3zki7YHjIqKz2X7d+X7YhiCZNLy16/lA/dhy1yu+t
QvidbnU6DtbpvBYNDQ/2ZlLj8bkvgDeFFuUZeutjUnqtcvlPBHL7BoJNs70jjUtzuMNKTzyEZzGM
ArKq5HoMgoQ9f0jDjV0HOkVEls0Y20sNNKhppSENyQug5CkQXDrv7agO/82n8NQArHqvwKNZ4FK1
FsIrpxbTW4M775lhQoaGyw/nwIjIzTE07DfL/fIPbBurkIQfLRHA/cPgtuCbuuJszbrzmEV+Ss0+
eEujAY0j10FxDPJclqsz2zgJOhwhFAQpW/wbOisdNFg4dvvDgtMSC6RlgIiFdAqXRUUjC+yCpY/5
krKAFm/sH74oabEBTEhDfINBXMDhP4lwKovag6+VDRvy0q5+bPwW0YJkVm2CIHitHYKXfsM2vk2J
JZjwYMXveyfkn4PgwpYjLId8LdZ+NVpe/wCqB/yyRYd45D0Gjmw4l+wy0BPrvLuj7DKmmu9drFgw
vC8bvJciFMET69MC8Lp5qg9NZSInWS75sQfl/ONtjuNKzu+EmNpna/Hr/BB/KMta5Q+hsEwGbYNw
3MRqQ227m/1pXRbNvPKb+Gf2SLjjLR9+qhKgTVtPgVCkSb2P+dwZJXlfOLxkfeYY60WFxsabzNyN
ss2nCTab7yh95kV3SLuY9VLEkoXewbcXwulYibBozE8yn/uJbeZMuiQB6FH31lH2L/tvqFfEyVJS
VMrLti981DGnJIx7Uqv9gVRsSXgWnk1zeED8ykdRydxaQI1QoC8c/QRyzScPpYr9s/4iCc4K+GE9
mcCIfYQgvMk+9DbjkuWIGpby03zdInxk8K7KRSVqemtLxA5sidh9veMbPyT8l+d5kdTJBv6o9aPV
oh06ni4c/PgwW9YBm5D0mPM+grl/Sjd7TfLgkQo/nCBzdliE7M3l0qkPd3eGRPQmj02DIaIPy1Rr
BDE4YkA58s6t1KB4xa/Dx9myebdNQAlasDrmhTOTICKUL89p2lO20A7yLo62NtllGzsQ6br/5xiY
cV1+ozjN0M2NMH1OimliBmW1aDSaLvDdKKyMyTL6VKxF3CpBskXfwt8MUfQbLyepFtInYpLPWxrl
23xtwgrzN/VzLQ0U/jez3zpzOA3w2zExtEgmz1v1UBrdHlhFrY9uD9HpyxrBUxRntSv11L5krCWt
LjPP4SOsoaRRm9HhBuNfq0Ws+T4gjbjR3TXJV19ihTCbRTtCnr/HdrujmmAk3XS5+rAwFlmG/myc
5GYx5R5c7iwM7zSx0nQayJj4KRvtECo4gvnjnomOq/1vX8UPHf966aMoPtH+fy6alSFmzK+/XGPC
VylJUJhiXN/eO09T4+MRzKTIQqphfsCiXddO6yDJ81YaYiK4LANkJzvZT1viBZkAVb6oBWNcbA+R
se5tR+fmTjVKHd0nB3uWzb51zVFIAhJv+8sIkdum3ZzdhejTIiDErr+PGcZGOsYI6CDXYdIIlUrl
pPZMLOx//nsmGEqgCex+9VvSXlzLka3+DHVbCdU9GtctWajr080SpLuQguohqDtzdlQLp0viRcLV
CP5hdZg+f0s8u5vPPYltkuURy4PcwcxFyP3cqq+k+h/soN3D/MTRHhsxnZH8AyP9xmQiF9LaS94b
V2nWVOh/svxRVWS93gP4oKgGYf/49y3UgMdZeHE5zsIOU+0BpSOh9x77PIV0vRdYS/2mYGfWzDDq
HDpxpKltltA936AQAMnlMtGv84VBbOaMJQm5DD8ZGrB6HzQvjSyixOZDWloKyPwZhUbQzkXBNVEX
kEgKUIQFWcQxUjW90tWE2ZVafPVfsGeZ8PZbAXThJKjaGMmNlGOm9n9o+hbG70eklR3SHqkmvB2d
7kRLt8QXa9uagx2gxN8+LJoXOHrF+Z2yWQTm2wTsz8EjPPFPvEhyFYJdGWN0E0VEHthWdQuh48Lg
OqiL4gL50b6yJBtw6Qg6oyvesNsu2NPIxlolUkshKKftgaql7s3fA0L8dMn2NKcaEsNmYem8fe2n
KuyfAbc/Q1bsqkuW7L/AQCgEKVQyjp371H3PK4HfoknkRsh4fa2QuGVGtVTyxHPV4cwHDp/Cr+4Y
pHqVRok9WPVqWESzbvD6Unh8GdeOzLgR55sl+vKdccOWhYze7WDPAepFnoCYX8/grIGupat0E2OP
wxVRMEmTXRXx1D3AWsTiHePVOqA3V2Mlw0fdlH7ywcLor2yS9q31n+QlIslwQasSIHoJcYnuGCxu
PdS4IGPZmblv2+6mBAutXrJH3X8Ka7h6U+iM1OuOePl2fDO3NPVS5ki+tcgtT8vTqmmGsyhZl+Y1
4SulX+Bk+ZtI+6q03spNWsCqZu7Wk4cTLRBwb2usFqAHYlF7f+3EX/C1XyL/EvPI5ef5ebXu5MLT
D69ORrQCjsRVgS56SjNjtHoMErGNKyXWKM6v2j+moGXCI3WdkXVCCQCaNDHohQ8hOPSH3j9R6YVy
yB6lDuvMRCY8P+GBCfAB/BQCaCfSs9sVVrKG2UYqARlZtCDkCuETqq3MwHRZRPLmvkgNFaC6xCqm
bCmwHytR0erz7rv/hXZN54M1KwJukPHAuRRKwJ7FkmrYBY5IccHbCp2YAo59WH7+yx8v/dq19ePW
wOR4VYFbrOFXFuhwG/5xYOA3yKy3Nt6C8mZvOJ/qXw+7S84KtLec8LuPfwGph4rfC+fHMEjCVu+p
Xr4oDQVYByp3MaeJsPEwGDUw61eOjd9ENDj29FYlUWklcslWrjP22ZhET48mZJ6TvFK56hPZi4tq
d9PdsSq/zLd3fMHf/Z4n1gEQIimtidPlmfOnmeLFemFntfzisx2YrTOJyzuKv8jabATVRgilohIL
YMZ31zH/0aq+wtRqRWE/rhrl69HjS0C/+TWt6KLV2Ufaj3lb4j2j+fSd5XytrSZ+EhmloQ5lk6/S
H57Utm5Ms9K7E1jBemgKfEULTEfXz5lUUsH+SJYJfM+woew6zawBP0kPAHGQagKEFIvQVm/eZwmu
11YbYwtF6VHVohACLp92UOpYx+YSm+RGUo6dNfyhxaMYwAsSLqTdlosjoxaumaBcokP4VQgnTkxz
ckETVH5HLTmneZe0MvjzVRvwb9T/35o/cbpibm11WLorz/Ju3QG7kG7EBc8s5NMbpeRuTY4asGxw
aBnqSJbTtdFXgy4EdBop+kJufG563WgLkKFc8OxaUgb95QJ4t6yqzc0Jgws1mITaef0LwRhubOgW
ENnmC9qNWp8bsKoBF7D68zXzlLzJZnNJ0XcARWlwW1wGl4a274IeTQo2ZxsgndosUkMG14SVkWli
ePf2cq1AqDIAnsTR6vMO6HXGDaMXL2+kMucUBqicelbI1RKKoeDNIE2D7c1VNZQGSM+q8fGEAVDU
ziZ00nbHjca6OO11ZkeyDwrgp9oswWdw+mOERElVwIo0E64eb9DsxG89/WFfwezdQTir8vU1e0tV
fQo8SF+z1kIoCQNYwbkqd+sgALm76MzNFGyQ85nXtoxF6vIjew4OOuMtTxWDjo3BWkTQfATSyWV2
8FNNWASDmf2N0Ao5j8N+VJj+eoGs8S4IIA503tMAJCi0vxseNgRT65OIaKOZ0K4GvxC+lwYAOA/G
1oict0ChlQwtoaAFabWaKbcV4v7s7XXZh45U3yXRmVAPJqFn8XIDwxRLK2B1Q2Y1VmjzO/0i4ey/
+TnUdXQD6qcWSOcWL36gJrqAcHRwlf1KuHMyF9RNsPMjcRLt8N6c5lX8PJW16o4iHQK3XT16NbNH
eeUh4eRM0y1eDOSJ6LDbygkPiw+6uBanPGuS7qr3xHtos79NKafsLRYmSw4dDBM8Cp5ndBARtrNS
+MB5BrANivO3OvUvqCuUGFZAg4wZbJcfDdJOUhnhgJKU/krgMFey0qe1KXU9vBrksavsRNqcSfFL
v6iRMpYpTEaE8ajfNiYQZn3gYR0W1CGPJVLBHPhaH71YfXYQvTEYm5mlX+uQ7d9x/veFxbYK8w0x
HfQpqHbFC29dN+mJNdy86dJpoy4maVubtM8cM51ElCkTETNxqi1f4Uhgvvs53mM7QToRxCqyEZML
gXXzEIcowpm2tT4lbDYc47/ug4cOWYvK1lfepXxonMhIc7Vedx2oQPzl32xyRm6B0WAKB9INFwLs
gJeiSWteBE0qY5c8H96YG99xN5h04F6H9HPeh4ShcpLzio6H5byUBG1SGGQNMYxNAHDqtilPKp/p
H6rrZO8mOX92ojTBzJyj8juSlwQk4YlnvnR4gP/f6eP7JaHgzfF7xxLAuGH6bEpiSelnq5zrNTDP
yf5hGGSnEFXZBvn3fgPQwXjGib6dRZDikpOpWHsEMFoW2zsNxee4g9fA0cRNi6HL+6ADdVjRvr+G
ibh06O+cplKrxM28f47ypkAk3CJ7pa/o5N/UeGFpw+MZndjehlOEUvrPQdRRRcl0TPbq3QGOlUxD
P+ogdh51hmGCBafQPMFbNqTcCveK9a0B18QhZPHIuMl0UsxSp9pT1T0gjQ///a8T6Zwh5A1bKxOb
xu3ldt+bdRnSeJt8o3Jlm1n/TKJUdwQ8sv0yCGScEgbLklYWRgGgxEHCRp+W8KBDaNUoDYNNIBTE
ZNUBn0MRs+t1X6mimqd4OcGLztcw4OWjwv+hxw8naf/5pE2cR+9H2kD/Jh7ijuyEzuF3dxI51mTG
pVnuMUdYaKOf3xtvC1hXNjbrnCmjLK5VSdJZRiJaA8etwcOt+YOaPXRQ6F4BItGWIei15KZTIRjr
6nui6XVhKr3uRpu7mSJR5gFluk1ZpwMEh78ADZhn5hROUNaFHf7PEpEbRUT2pm4WbmK1qhVPvNIE
d37cV61VgXZXEV7Bpp1kO73zPjeT888k6GHAshWHab/SReXiYQVoSnMMrf/Y4NNLDBl4tBu0snd9
nybJ3KfW+VqV1B10NC+A+hXzlOhzUp/kGMfm1hDm2A8zqni2Sujfsg7tdKWxZHGarIq7kZ1elEMB
a8cEacl1qxkP3neSXXR+vn/bOiVHoRoHM7Qb7EPM9FerD4ihQXoLwWNdhSgNMFi8e10FXw+xa/j8
e2He0boyvBoeK8IMQ62GDyf/GJHOH1VPvrmfkm66ouZzoATH1kp7VrMRGLl3fMndXSai+MOiktMk
SlkLkC7k6olG6d5yk0kXCBIuhwg5dfTl4aaM9JERy4wjvgtPluqtx5gBX4APwgWGpAEZhNOHz6rU
xU3cNBLBPiz+h4vs34i+5qlgJB8VZR/g8plO3HSOwwbH2QEnSs0xuoAYK31wPVFGZnjJaFElFSN3
1SjPV10Y8dEaQF5yi4kd+D5rUsvn3BhruY7Zyo5RHz6RiitDMhwjOcszDQBTGcIdXdG8vENqg4d2
fVRuHx8bxmVwxdOd+yAPBRpw+UVwTmpw61Lo65D7Qi2ulT21ye+vqP9/lgE/ChlZGp2sm5nsTD3i
yXDTWeeyGz5lJm3KdbeF9kkfXEOcaLRGYutDjkQakT5e1f+ZhvwBb1vHrYz98WZjPnVwZo17H5ff
uwTlo42i3q1JB4+im/btPlPDiRzMxL/X7+H5qJZxyKqboMsqBKqp1puhS7d3ZdVkXyPOWBLfAw3e
bDmmBKly0e1UgFWVWF/rut2XLtl32zAfwIC6J8tBlFfblWQlfpBgtumMdEuIfdaU7Ew25lIqFMEL
VJV/iVkppHI4/4QeewZiQMkt8ZEZK6Q8FaWAUMPxXpoWAZqnxp6jLluPFJ6DZKM9/Gfv+WrLrd6O
PFW1FI3LZbSAWAlmg4Aqs/lDKrO97d1fxhoP1XKOGKpj3y0CcQJKGy5ccefeY2DtJitH7JCA8Oi9
vkJKeMmiiFGfV9OFyJmtuMGtisnzzywUm1DcPz3uKKvhgFuEvcJi7u2kH+5cp+sFu15JGyDbzLfb
4GBQVmPVYpyW9cgo+e6aXRRGdX1EVePs/n4qyxCXd2ODNsqQGSfccl2tvzJyWS1KGib98f1o9rUr
6k/7VwX+5wz5k2+JU4ii6vTz4wVh3mI4+aEn9Gyf3v3CUbD8scEAFHIVyX/N8BbKbLwU8noluBRp
KyekX9cj3PfFt2vrzfnBTcPZI4UFAD8bArjlLkDWnGIfudUrry0WCvybIwxSDmxUryeV1KlmSrrE
RvMaIE8xByOQEKhGbQQr1loWKGLMyT5s6PfcMqUUPxr1fNqM4dCOipxVaJqb56lTmzzejAEemu4n
F8I0FC9ljzUB2Kv3b0K04C5e85hVl+2jDl/0hQypDT8RoeDIS7ueN9GeXK4rxjqUzAR2tfawvt69
wuTzBn0SGKPJrsAqYDjR3LA47qkoB8E9ezmajC6fcEan+m2GTCjoozjARhCZieycDczaW/QRGKsz
o2yfY1S6PjyYsl9XzcfKuYonrbSYAZ6craSKW2Nxd3t/JeSDs8RvyIOI6ZOncpg7FF0AmOMFRaI8
KN0COIK3Cy8cQBnr/drt97o6tJ74T8HxGga1bv4VOZ5VRij3upcHDroudO3NJSN4pDYfy1VtvZwk
uy6m1f9IojwVCeRqkK2MJ7jII0G7VzgZY3toYMiy9VLlZcbFUNTlsKwco+hEgzFhoBzgBRorgMQB
TBXCCBU6kNcpEJ05TnLTR57/LF5XfZwrmmM5gXtbC0h6EnY8Rf+u40+xMVmEey3kmE7m6zPFKgBt
w5vlFiJjCtackZ+U0TiE07Y2oecVMEoMBeAA9w0rgnwNwvhJbX6eYC+L7E1TIDlFp8rdO+VnbjUk
5llklXQbakL/AlqFGBPTXPNI/aW7nOxcfZXDF8xvqlhWzmvMuNs+yqnZFu6SPKqiDf1Jn51LCTHw
xfHuUYGpiwFQNthKA9BxqTfYlT9p6cBHjDG/6FdbxMLMAKVCmS3oWnaHq2LPXORBEZC3ZOLtf84u
lnYB9Q2bN6kBx7QfAld8XfGVEAxm4EaJiUIjA+dWVWN+IUXqwl2CEdL0+mkbvNPoQIJas4aXfM7k
MlYor10/B1TXOy2KN1K0Zgc8bfvxSNHiqnkYuwF2zG+4CHc7qTNM6yWn0i4WbE+EXlDH0zBQqiBl
CHncE6sIJUlFPC/wH3YCKHTmGFnzllL1ZrPb8nLdkhaB7A4xDfKuTkzc3zdYrmpGLCFIJ1WsMpOE
AdObEcpMwrs0yRAy/hxDl2FFyPPKqaD9D5K4MC7/5j/B3sZ7RXtbpuyPnz9t6/XYKIcblsaDjBJ3
/qxBviwO+DpVrEsJ3oOpRYxGVVEs9r6ftxrnNfXf0DAFdiVnN5oklQCe/vKyvVLYHSy5PNyZ//+E
0jAFAFMmYf3k73C9jd9nK+ragfwP4uzA0cft+7adF+MrZWsIrIuult9uBwSgWA/QUlh0/CpleGkT
ZthRWrWF/Q+noKTr+aFpGpH9jL9+n+am9sfBXQ+4r+BNQokhKp9Vlm7jRhcKO5sGfNGVjM9b1N0E
ZplFKWWS2TCw7zdEUpoNjM0CwXRADkloo0gXWARvr2Kfd1k4d2uMuui7vvqiunq0kIjXUbOS1nxS
0IHrbE1M303mR4u95eqsDWLIqgRDoyOsPjqHS0gT2EZOJDTuoKlHOt9Bi/sE+/R1RtUXEVnHZ8m6
PzfPumuXxFylUa7yyZhCDw28VOzWDStMEhCt5+qabjad5YNZfYcU8uXzPYWhpEwodfGXIzz1gpwI
s9ANfbssy6+Kq4tuj6uKhkxwpbLhacbDKTyjtoKGT0swb76IzrJY0v8vY6hqJ/i2CqMgiroCT2EZ
aXXVuhCkB5Um9MFo1aAOXOvv5/bCEi0s1W6lwbYIN4pCECcoCEp22aOr/SV0vgTmCM9o6JscgoCr
F9UdHEr/zuMzFJfjfVKWKlot6vGU5HC3dYxqnfplE5z3PTCYum8JZaf2wDSx5iMeTEuVkSO07QYJ
DQ5YHQMORPj9gZWtRRXkFEW0pUYr3e3aw2Kijy/rMrZUHTnwPpsheTjItasn25v+9Duy/abWD+Ny
/UYGQxxoqA5IsDzwJ7snVb4jD7aTOWW+PNRWjfIG9cH336QEaXLQcuf4cqJV+M2m28GURiS5yw0L
veUv2oxoWQzdIHKXBFxtY34PrQyv4aIGF7HmtlbO8Dcvu7QnOYKuT67XLlKqmVXSO7+3LH1cuiLK
i8g73NLmdKyZfWMxkN0W3sGDXJKXck8FZEvL/vsJIEhZdpQdby0N7y2x2mwgY7fpOXU+A4NViRvJ
FavyZnB//JOoH5MIJMBcjZWtOorrVGPLYSlfL1GswuE2+DOcNa+NTul/5tY0Cl/R1c+rB7dwpWsE
+wFlbfV362UP43c4vA0SGZu4YpxGh1V3S8AggeEZ6lfRtYgCD3Vvi/Aj/jcNSq1LpSowNViqAW3d
qvzf1kHY5n6qknBlUcXoksPV1Jpm7wxTsfFvktHJqJoZPAAix5eOaGte7kkIq1EHTFf9/16vMpYa
SbAYPC8WfQYcnDVxPgmYwrRsIVilOvnUNnwnB0iu84szxLS+ZedAaejCbRJUks0RtsRTmT5M0gSU
WOy7fIqAdUcfgC6hblQ8xa0t5vNmuZG7ZoHq4jJwHGqNVZs7b0Y+LpiKML5YW4DvoQFPIFZpKfYZ
J1ySAQHAbZYhzNKHPsQVaCliL7Sj1+gz5a7Y0G81eNUg2m6WsrzXFwRuXUBHGoHr7NJP2Soe4EJf
AkH7lQ1KG9Yx4jUwOUl71OLsKuQCNBk3hd9/rQ6eQbndns5eFdw1GaeT35DzeXiaLO774LlF8eGZ
X2WD2WDf1L1RnWY+uxhD7en+5XMwEzyq98yeO15GRUZeiPHP4IMVWoLYooUInPZp/n6WhBEvNiuZ
KJs59vWtCVFF+qoa7O0H8LvBeJoqIucA5DWQSFX2ZBahYHu587yCH59Dryhq7+aEQBr3zUl32LGJ
aGmZmiB8DeXJcmKYoh8ss3oZCkRDWHCVVvZqDdN3lD149WLtGaBLRGo2dLayZD0x1QOKyNEGEXH4
EK1D2UW9W2KYEGL+y0WT5f8QAUmYj/mmxYJSfcWrLydcdaHzDZl9IyWOT5NJ2Qj6F0G57qs8ETWQ
g0Sl0/nPBR8QdjsuUTk5Q/MQgkyJ38ieypcb42KNwOneKJ6v/LKQKQ59OQ8odbdMmiTzF68Q9geL
trD9yQah8nHEm8cdWeBeHUDs53ZWjhmqjmhmZuZvUQGqLL+M3uAwC1aYvLf3vFLvGHUVfWkjqL/F
GZoOE2y4KunyaKJhIdpIZzzdvM04u2Un31Dd2biAlBgNG5DdEnh0zlpjVOlstoO391O8g+p3n+eb
P6bVZO9VJ0dGKmmKtQzqkT2hvzYqb63FUbvIHmRR168Sg1UeGbzWgV6pa48PFgxo23hZNW0ZHynT
wZeckU9+J1ZaSVOaaZ9Me1v3ui7FISP3TWmhY/ei4R5WC90LgQfWCO8/H1XDYV68Hth5Rgzl6aBQ
UVqIFBe0vBK9eBVNzgsa5/aSvJMR6mcp3RFFb0dmwbmZGEjWGyuj/XztDdonMO4qpRnYPf+uY/Tl
mx9MDP3SZhPArhT2px6FtRA82kbRcoZPBYUb8RndVr1TrAZa4MRtCcrenrs9/GC/NMgrXzrP1SJf
BIcnF618D1qutduCjhet9ZfC0eHt8ujk4a1GOXGGXBT5m1WzJ1QNQeAlbtFRta6vlFSEmE+JyI/N
DkMopoMkHbaDicceWZ0P5YaznjP18uoNfi3JkeMu9xaJl49t9QsUfpPkwv+zIGyJQ3oZlzEq94N9
Itd4ETtn9BNzdn7EPdUjLv2GtlrZ0dO5tJH+4xxXTU8OBt+97/iEo2TvjbCGGN9TGCbfICqEVK7N
prYsOQ2qo00P4BukKMnKwVT7nR+HM+/YASIJ/TaEMEOhRMCwcMqdCXpoWyQHzxXzlWw1srdeSO6j
7egliSIIW9031fS4NvJYuha3ZVy52PtYbZ/Y6wCijpeXAvBi9miKXUj8O4qkhuP+VDkgxZFeOrRb
oDc+jL63fL00652oMq5JaDBl45/WOx7ttw3a2XzCXnIAZHgCos2XE1OGADvdaUkwZnqf10cfQNxf
VwYNrNuG1HvlZBo74vH9L3hswNx6YsORsUHCNr3XL4TOVbDxdfx5jVoen+ChJYCyqlCxjieZZQwx
AtCiQ7HE55CryARIV/yojpfYuArCVRU+iDiJpZlm39SeKRxeGB4SRXuT2MUxdXQLBRqNr7pNGPwV
Ta7Viwfb2fUOOlxEkIbvjuaN3iUXGUO6Dhdad8Wp4bGp+FoCiFn0cImFlnGE/YjWknIKQV2yBtwG
vDHW5mr+bxnM77P3HGI5uv5a5Wa1VB5ReJbokHraoV9oki+hqidPkW3eXqO/mGmTDcLtSLqlj/il
H8w3Nd3QE4Hwndi1NoRdTYVbbsGzsAFjPR3iE1vC4pTyMvixYk6X3P87lJYJqeJ3guBET9Sb9gub
U5Z0/j1m7PslM3sRfSOqNW/n9Wig+ONYODI34J8bou2fsm/UvgblflARWKdYk2Hf3ieYUad1Wgy8
BQtxZh7YkBR13TI/8dMWAlj7Icdv0aMsEBlGC7IyRnzGJcH/reD3LudbkD8hFznq1Oib5UWQR7DR
VFMUlkycv8CE7cVJ/bMq7IlGfYII/MaieWetnVj8aojxHVcbyASoiRMVjfrWr2Hbad6mnmsPAKs0
nMm8Cllkemxb9vaUrbjJZlj1cRO+ZTJj+Nu8pQOS+Yrmcu8OyhrH8N9TeEIrQM8KLr96Uwd1+PPT
x+w6m9KxKXVpfj5dZxjDAmyBd0vj2TJAuVlPcXt8yqPMEexo1V0T7JLCLbm3pGx6Bsks2JEochSt
awkGsNGcwbCbb5ufzasf6kuGAsyYiZEmLVzahqHGSbAxYlHsBXuoWSfFekRmUwg+Kcl+fohZ2nnT
GfaZTsLoRILLR+KENrZUGQyTiglLmNo2M4zFCqoPhh9lfN0zQjoDXIJS3if34+hQqnjo67qNzf2e
IW4zuu6xoa/6/HtY7QoJGi3Bz7wjJLLPrP/WkD7hgi7RVrOGkyf5vbpeTW4TgvWYyCjJ63KAYOYa
ru3PD/ogx2fGrDYrWeuu4QtaGY0rAhjBMPXMKXd/lM+zNDvhZ3lPLsJhahKasOZMRScPqb8pOiZN
zg6mGcJUHPsvO5FP6MwIpoNht3GbK1StV3ph2F2lqyOwIa0sWsUbNQmglb9xI+NWqkjY2TaKFoZk
TXeqRntP2xEG2sx15Q66a6cPdLQqGUtYNOmCBkq9gn1mv6bHYq5O7o5Dkwez9d5qd4PKeDnLLikK
cSkenv81j4NF0KA5hRUO7qbRcMjcGJ11K7vH/ZY+wr1zNGzsHLCN2lYh2HK0T+659DdCaJO7+Lbh
/evb+AP0txyGA81DP+LlceduaxP3iKcqAtWvb6TLnL3ED1ki+7q1dWuDDSbryzvEnSTZgAyZadse
NPl7n1Lm9UGBEatppRqMpbj9wCRNQUevuN0O58+uF0OjGtBENC6GOQ0hyh20QAykOmV4ZrKtDA0N
XA8V4qkP2LddNnFhZqDcPoygv7QSa9VXMjgbhP0EFyXpAjlqlmJZ95Iog7dOFkwwQZ4BYFqB/JD5
8whoM7wbYstDSG/KX6iZVhDfZllZuUMkHteNdTeYkDrJbIkB+tltWP1AMWKR3ryIrpoSG4+9lroq
s0G785SHwdMjg3rh2Rzek3kvdfg/8KakXce6WbrtyJLlekrXTAVtzmEnJdIUKVNgIIymdZsg4xor
b3bRURLOo5FoMwynPx7qYggPJyJwy5vDD4JHtbEnS3vGNDNdV2IFTi1YJ/x4Oy7Ogj64aHlIhUdm
3aFfd6ejVpon5E7NmStoPGFy3/RrHxg5F8H3REpRMQOs8cKp1aJlYUem2d3XynXeiV1pmWsUAl/H
acyDJUxIUEb+P+tdAqdzC7j98lCN1XCXuoA7Np+k1yf1TVh3TAwdgbEkuJsN7ETeUHqOwMUvRDoL
fRvJH9aJiSHo7HgSp9HIueJWjUUIcaLEP6xd+Hk70iTEAlUgS3oOx4Yj4ZYyADTE0sH5f4QnQVsu
ySWtrFGS/q9qzPvzSQyKFpvAAgueO0CG6bjrP7rWHbAkCWXnQtTwITjZnbHEbVW9YI2oOLD6rOXr
nTqOsV6WX19GdK5Cj8t55S8ifUvS8/Wos9EWU4BpEMklYeXZ/0aXtUAqjhbYGxXvHqNJNP3KHDYb
hUP+jUTDmRR9cp0Z6Ycj9zb83x53a7gSd2iqPLItXjge0pxPr9txB71DRGZ8+EbxvTGKbQqaspjI
s2KDJjJZir5dWi4jojelsSzHC83N+SnSdjPuGi2Z/gx+oUBoALCaHI7MGELLFloNz9v+YJETKOYD
uEz/rRyckf2rH464Iukv4JciRFAMA9nz+TNDKrt2YJAc/9+kJQgTkex9EZPhZynAOyuqH7wwaHkj
yeMfl/pM0bwA7U15B/mdiEcVmf4jXXBsL7sXVJAgra1b5C1u0BevyMNJd8qIZ+Hih8dZEX7S50CT
+UXkn9jcWm/+wVkSq5+qisDQjAF5m9U5Hl/mp9Qm5uYRXnNNBGyKIFWxxFZCQrDD5vQ7wbo0GphO
RBDflapSb5FsVOoFxD8Yi3IpclfP4iXz6ZaPY/6j04+glAz3GGfS2xuRnpHug/U6Y1ixHp0p5y30
Hwa0FlDRuP7J344DTWdpqy5db40jJUcu2+PyldTqZRxU0i7DPjw4SUmgv25MuULZCBVhAJJmQiX6
M9Q7u1+vllNpaHUguOmFhykWRMwizyBUwAxPzycVG+pNO7E5X2SCYjFWeaTG/d1VsjUqM92syjUs
i7atmoSCRFCYrShjmhXZtN6OR4qx3CSmp5e+xecsB52fjz0rREj5pUUqYlbd3D2g3S7vfwuYaqAt
PYyZi7G3RbyRLMsvA1kB5/pwRfIPqUWrl5YgA8W9cWwcaFG1SDihXFSkLigeKmMd/Ogbp6vpRVGl
UGE+/R4Qe5oVjFUsbmZPdx44ZGnj3gPTFD0Guabk8kGqHWJpKclX2XyVA1c6USjGDV8fPzvK88qJ
eNFPftJZXopmyYhIvBDdSdDs/8jU/e6Tyl/pjsdqXmVtcCtMVmSSBOymLqp+uxtPeaSSi+Ln84hl
fsO7wGn8KI46VyVhWNoKs62rikSDgvGBMwqzjDw2NytNGQsEc9efW3RXPzjm+FnN/pBNC3O9MOL7
5kRxdiraZUBxIUBFhmciz+BljsvOBC5gDWkHDhtRW2qP/jZuHkVmk7B8JASZT9LgUQUW2V9nOGMZ
vAeCDQFcS4xUw1e8dd3r3uoAZ140z15A0XZAwibwS2U5h27oxwdTaInQuduO6CCApSlhjYaivhQh
b1k8gZE73lGTntCU12SrPBnT/0UD2g1L019WpzkILYHWs80Y8+/Y51zRcGznoJPRG0436ojapfxt
DL8gjDz1wzPoAeIJUznUdhJ5BjyJJmknF98mJQAZyGnHoJ493tocUOwfbZ7cyvY8CaXkCvv7A3Ml
1NBpifJvDpImoiFWvkjiDlvpvoltx+BVCj+2+HgsGvcUitwhzfGswHH9dNV5v3ZRz/OwiL+kjJJN
W+qCftpwyA7fduHS4VyqbcUvW5EG/GdScICBXJWjIFb4WD6Z9E5er2PNG16YlyRX+z01agrNcfph
KG/UUqUPQQUZbA8Im7PYupvVyLqLdALtNaR4r6Cta20a5dEIxtXUr9OW68vgZIbhdRk3zVH64k+s
+JQUBUAWEcMv+03DJ4QKZOuiUd61zXlgq6Seqh8qEcUwQKp6xHhohSUKh82AEOXn4xbilSVHdAR/
0oF8ad29lApTAwaO3klv99fBMEvYJSEeWmQgwz4Wjr7N6KUxdHXRSA0IA7oKtRRAA8elM/LBO3p9
fx7G6EQmgS18HFApr6XRCWK2CStBUND2Hk1bazQLMdSL33uEZB6EBdn7llPQy0PliCXzm+XMuCZZ
L6bM+eLKK1mJULRzoALqn8rkeneVWO7SlukPrjg631sjOgwxGwA9LJBNTr745nBcBBj2PhVWBXoT
ilHEKNVJYdG7m+XsCntLNOLX9DYlUpI8lH90ApLRNSAHMS3WrhgPc5AgsDTzszy8FeobUIt9CWZb
Do7oFIVpduLUbPf49VAJtLRL+sIau7E3eEM4wTZLzlsVopmn0nq/5qHf6qOOFJQiR/LgBmbFoX7H
AzW6y0L/QfT2yEiq4Upkqs+52np/Spq13mWHmKRmmFqJmJQPWvs/w7pop5huVwnFP9sjbrwDGCw0
M9Y+6IrCzu8c2eULmvqWDK5+7Z2Faam8PuZErNyIuDLiIr+1n7ycgpWqfGubtNmcrxEUnpqvckfe
d/rj0QmLwjEnEO9bpI8p+LwfCYOKQd6byOnu0MqVrsN23hkIHR+6pXwvmUYbjm9NRJpNv5cun2kr
c3Zc5YX4/5gopHhNCf00ukMvHlLfWav7GFgBQUAKcljN1QNvFZ1sc8npuR7UMR1R2diJla8WAjjf
yJXSFtHmrIAhDNaU82JHp0NRQ3kTLjgbM6Dd1fLXtUgxJr6UR0AY738q0vNjkoDEWBv5hXUxa4Al
TwHqjSY3EuNwDoW7/vzQqtH7N6c1y7fqT/jONNC85Xouh0sVoA7xuM2xnwbi/G62qu2vubo5OhEC
FFX+CCfruHUKJcdKI/Dqkk5aYM4u8cVT7cYaqun2ACOhNUUBnIigDVdQTnimSFr4i4GKSqwZeIyj
DiB09+ZauKa7l4wC/AKSwpBTA3DNYPDa3oDISRsFJedvrwAgTC8wSpJnpwMo4Z7bd7B6Nmi1aLY0
vmgR63nmVvvG96OSRQwDlbyrKt7tL4OxwNvjMdsCOBCQSh+aZIYZsc8/7Ocg/lT4baGinrys1uBl
J6Q/pYP6NV/7LyVv/asLi9sciTSTAkKqZ5f50wc24WEhvfpn/cF8TC6Erq+Yk601/jsMUhhOOSR2
AfsJkqJRJ3FXCrJ+EOE7aj/RxkD/c7LTuAWe+u7MdrABVvo167bHlXTl5n3C6I5qmMFgmlm3Odg1
FzYwFPEEAnKYeGLUkq3hDIgQvi2vRUYwTR/Ai6d1/jBMOPbPNbv9OpAhj5IggZ9u/he+TdITgZ45
dDmwQqAR92xHVgHy/v2m0knWEXwUz39rCRVUSneYhatOVrKHda7Gweqd2KwuWnfDRotqndlyr/pR
tULha4fc/Qbx9muu8HIid38XJEbAufWClNodVvwLuiYIbU1rM5WDNW93AuGsQCrcUr66GlL4KrRg
7m2yv7nz4xGG6E/Hzqn33F7ddjxOtqNMfd6PjBbdIudOrazJHqnGGyUcTihxAwGNoqGKl/JMpZF6
9CgHh5m7j1v06rrE1a8uBZoGKjq4L/vgyquDpdVhK948dHTrC2Hyawhmy5asAgU7+ff5Cr0k9+a9
HQX1agyZCgTJJwVTGkgjykSJaGApbe1p7/BCUC0f24Ssa8UNmddsbl1VvaNDyWSPlKyFxFz5aO+G
p1dUU6iKN1gchIV6l95vyunPeWlvcotGr+2mwemeyx1zPVIeKOamfDzhsEpWVGvr4VAUjXd66bA3
1XY3kSsnTgzhBivsRbMyBR3wAGvPj9IxI569DlApUQdmO4yj2tCoj+rqkdDmJ1tu7HewcVvEjVZH
9Xq3XvvC1qqSYJC27gBsp8f+P4PMDtO7iBgfo9M8XB/yGMbassFdKGrO1pn/CFksRolneXdthBVo
CH8b75PQ8LWcL/9pRP/LGzSrKI64ZoQw6Y/USrIfhBBVDPMr8jYzqnNfh79TfhL7r77jqymd/E0g
IfmbY/ywxU0DtEY1HrXeBnPeA8NHK0SUnzvVRD2iZOAWCgFEk+7tvg1hqGGXph3ucoRhurMrL6kF
iZWcSxF9/txl7vZCKbCFEK59qyn9RTLTX+vkIGdnMfRiASG0t56BXma3YBj3RKxtkG1yE0D0VQdb
zvV/1zoKxP5+XmG3FffLWn3W2bBmYMiuTC691uud/YLgg+a0vuz2pY//jMlvKalepgxS593Y1LzM
oICukwssVlyY5jNcRJL18xe5tlho8XpN3lvNxFrge4C17EHkkYMe/DZewpmcY4osPaQQTrf75UTN
NhmiqdKMvV6p3DgxOJq7JpsniECldIgNn8AjXXLAAg5G9QBy4IPIByTW3omdC8V9PQJbJ7t21V6h
E9q97G7VC0mVzvb26RtuG5c/uD1jMHfeA5jH4hWisjDhEirVSGMnqafndvrPxTUDXdhFaUOvHiJ8
LB+jGSu5bJdivSw3RNo1DqtYUHV0dU+8aq2FPOb9v+Dk2bl6faWAxwJFsRlHFml5M5qCqLKFp/Ek
fAJELfGOIcCHHOYOmsgMSqhpMLwW2Igc0jvQ5FLcfCDjHUqNTnKiU54RdHzDHDg4q1aRoBSSZDeG
YQROrrXG6mex+aMRhxgFBeESYE0L8K0/JT7RzSlQ1RIQ4QBujnz4iMclfKmvWYUxVehnQcMv0Qz1
ydqAK1wqBV98bD5PAu5UeGWpWQdDzSTro2htIjWX/101qlI2e1hs6PuiVlgdtmNlui1kuXs7DTix
ENQciBqaxTsTJWqpL6D0jAm4mgWvPSLzfz2HWQ4HTPYmXViYPMmacQbu8Isk8lLTMkRVxoXEQQu0
YS4hfT89vduub2518fmfTpo0C/8DwveYpOITKyspL7CMSFaRmYWu7HYYE+7Flqq2yR4SuB6uoPBI
k74ZThXnCPIrDxnqKRyrBKrY41jTKxcRswGgk+UJxnRZe2yKN1UEdun/gubgy29M64EcXH99fk9p
Homp0lsZiButXgILPcGbO0hwLFzPDUj63x7FKzTorENAzE1bvC0Cbor6/BjZOQxTX9LYXWvi7jva
cT0JBitW0EL2YgNhgCs0Aun1OCZoms5kclTQ8h+29uAz/4p18G9P5RwRKG7aHJOhCgrX0aQDR9GD
Ay50ufnh3tnfZiKhHlHsN+kOl1s3IrpRTNCGykUZ/CRZ3eMfqhkk4dBg8GMx4DlZqotaC0PPkAU4
8jrzJopusjuRmdT376rYMnstejfLPZmMY/kFmNR6K9MuIYzZSdHPDuijXgrLJUnhdmC7IYU3Lq+u
+nenrd8j5dyZC14MIBXXYRI8O7gNBZexoRPODn3wE627gmj0wEeibP72DVhxrDNI0E1xHiaqEp8Q
T3NSN/OWemwvVLVXBGrOhcrPXIllnzOfbZQMFDPL7XPi9VcWtuR7LT7CFpfZNihLP+CW4x2ADr1h
7ze6rCBJI24jPn9jIydRTxIyfKHR7ghp0QqPvr+XzZjKsHYClQBr6cOeYuIhpHBGtwo0dUVY1Kgt
Snn7FFEaN5C+pxsqRrF+yxxHLgX6ZQgBUFxKZ89xB0ekdcWxPXe95stTWd8z1XvN8OzuNx6Mhxwx
fO3v0p6DILj3W0GvF3aCTVAd1V/ukIHP+EMLsnljCFqSn+8OKXJt9r0qgmNXz2JgkppFNBk82hj2
T5N2n/F78jZf7aIYN81KFR0KqMAIpsKRVtI3fxp8bDGtDT7vl9iEW/1QkPXN+PJDW0HfQPPjJesj
l6zA06C4lwveZ3vvMewMzXGx+na2R4RW1rOPT1GkCp0j7CaiHHi0zoIRiJedgTQOAQGvWH/0tY0/
01l9WqBNdbtR7lwZJ3RAX6Uxn1R1g5QfIxKgqfDMvlfX3jL5Dh+Kf2PG1CBiMaImK79mR8F10BzM
vJxAWPz5qoIHD3q7nXmfFwfbal/07H/CPxIGO/dZBVXvse0bn5j9aWeNxffRThpEuAPaFF59a3/j
wEGkBxI7eujC+x0V9/oC19HjinKYqHlVvmF6/U6+8kDI3Y8yXt2BGZbCfa2wS2SORAzvTxorZcpw
F5usq2PMErpAZqG8IFcSgA1SCXAczP4Xynk7InOr5Sxm064j4nrOLV4q8k1hQazhTmAB5gqZ8Qlm
DtY1BnFvVGtwjhWK8q4/NL+Y1DT441eYAme74Fe2HvzkRs5qoAYdq0a5wlziZz1rup1PBSnrQnUL
AV9k87HqTw/9aH9mNHCGEE9WfPF2Pnvyo6V6/BjuF6rT1p50WsgWlXu4wqTfOSooHAlV6IsLr9V8
t/fkbMuR9JmWVUw63QyOt+Lx2Zm7ETiLXqQ4B6T6xgJg0ldIu/MPeJZ4PpBgyXzbkaN9+2UtsT3E
OcRWDDC3XeYZi+POOPxqVyZ5vSGv+Ip3MOSLK26nYmzABi/9TSATKM5v/7O9e9cZvM9sdoZzVp6C
taAjXeFnR4BOeDToSHs0nluPKIBCfWYBVKh6uzDNUpHlPhzEYu/PZNP+UAgB7ISReyxtqDj3o7fd
BQqtpen+P1xhBICccxwZVs1vMQSMu4LTSc8RTF19dGvF4rqPGuLBhRzsL9qx10/pv9t0ovk+ZSbr
bwuZKzHBDG/C//KA9tTqkeFeSyXweokcRXTrbf5RXxQmnw3cim3wE/JSurgTu+Kn5bT4a3HAfN34
Ozuvs7iKJGPCEfE/8/PjLczNnZXDh2CvswOvfz6yqFzPGdu0JxQJd2eTmE/zf6kunLyNO7349tp9
qXROdh1ZGRY45cg0tom/DvlcUeqMMP+txiXP1sC+aUO9SZsWvDDL7kS61wbgp6gn3sVDOQrQ3FAS
3N+uMBLKum98Uhev1jBSseQ7QozJlHzqnjaZxEGmiVQC4JwsM1Qu2CuRL9AFAtIvTAfzuTg8LLjM
UOZuE1RAhtoYNX4k226UZRyylU90dfyKJdF8Ak1rdBvSaRchJRDgrqKo1gcmVS0zkqxYb76h/Mxo
SZ3NWe0OGwdiCCT7CMHy3VOic+KO1Ank7AcjA6Mex6tQ/0+sL+0CFdUZ8ulvpJZa7p1m5LMbLCKz
anDVbTH9UKDC5FlhZ02hAO/ML93zjByMN5yHx6oviCv3EvIJ4lm3VAEve12fFQkp2TWi6FyRWXb3
oLQp29b28+PmJ1B19QzyoMUMr59EHoGaMwo7TrFWSy5lfnwP9N37tvcm41WvVNxMCdrQdhDKCU/Q
kuVB0ro+Mr+vIVPLfIAVIGGWadzhr2CR+W62KouXWpiUD0qFfV7Ljz7jiYM67WUXq7qdLzqp6fqn
ZxJrAStGen/K7Us74SRe7QuKBfZ3sDYYMlnGPxAykZq2FVrPKcNSdwMJ3vuzEFyu3WvZH3Ed4mkW
vMvB949cVSZMpcit56ECfXX+dDfz7ie9iUTM2doahNRgluuI9frI5wTlXVowyggnfVJhvDzI/KGe
3K99/iNykXK99Nvfs7X++Kv4JbR4MtwDdY6ABJ16ZQ7OwU2ntiwlJeQQk+KoYs6gAxILqezExHK+
Dlb5akIfac0OLw0lHDpg6UUUQudlMJ31ItXdVfWE+f7dd6FquO62Zv24d5iKka+WxP2FWGc7Plm/
nwf+HDL9BstiJMzQjBnNZqbl5lVE6b8RJ80eXVVzLftMBO47gbIWE2l7gSBnsX3yWQ/mTYPB4plu
3J+7QhzfvbpjB7Tu5QwV+MJp3R8W/juZrDjxQuTlmVh7rRVbAS1DYpjeEA3fTDmLC1Tld0+Qm61m
JFjn9TpllM1Hi7qgU2VDPZXyKnydk3jkViTbGbApV44z8RpySXdbF2qqWP2eIUtrKteH3fxWolnW
VenrijWq7JxDUjtbogCvE0gEAS0wLoTYMD/ldr7I/ee+zpZJeKtY7y6lAQd9l31hnc/CMvY4ND89
BclRFRSbaMttE1O/uJrUt2fmimlXP0Whq9ND6MXoJjSP1awIZFKp4moZELd9DWN6HlIWw/zFM2RH
4lBjU3LlelTIkV6VuQvuViXJthgtrjpvUDOcBLW57h0ppaMQFd3wyGuatCpYYlz+fbp32aLgaf3Y
oAhdiMKI/4hrvu4AmBVPGUfk8SNe+evxkHxw0beD8VF7Eirv2k0JC8LcMmbKpo8mINby4Qt0LmUy
5y2iYXW66aLlo2vMhBhDOYzrH1DAxHbEvHaRvUz7xhc5kEDI9PK8Ef2LCKF+iRRRZSfT/YlbSI50
aukX9mjVFyzxtgsPRuOf8C6Ox2fhRnc5v1qM1jEtSfv6CQGbyrTgSisirB/LUpw1Nrlx4R+1F98I
+ifDVC6CGxx7upMsbFN/DDfKm+4fbsU6GxHe6Sz3iPrhXzV0x5OESdxsXHjruHL7TQmm4JTq9J2w
lHpPbvKaFYBv0r35t8PQFoRsiZtAZWN0TPktSret/gqIaBbyogunkoJlA2KcQoQS7xawDKRC8vKE
BkZKhjRlWz3Vj/FWdnald+1YZOOhiC+F6DXy0QrwOVb7tvDJZ7PKQ0brf4tZ3yk/WwRETaA5VkfL
LaERTiX3AOWnUdQ4nE9XjAklb7K5/BTy/H8lAkC5ZZEFfgKkYZ+SsYx+wCII3QX4bXrBSorOKFy6
TgR8MptL9reObjLMtVhTdCm5NQPNT+QcGvk2Lqbdnh9R+KJaLvCZ0rXz9sqscRjiN3MM6+du2uXA
dMt4iIvBj2SmS9pb6DTp3kmmLDhY9hPyBhlNKrMxbD+3oDa3GEug+QmPlRkBCBKRSBIVuAvtBJ4K
RQ2l9Zp8qntu2xBzXs3JMvWEOmWQXbYhWLA2HuB9Y+Fd7cQY6txj3xjnW/1KIzW9yefjMGnuS+69
j+LxwHEzDhX8dfd7n+WwzGbfYqlwvdGaYotHi25Mt55BrXAicCa9wZAAzgTH2m5JoEWpOA8xVRNT
EoXSSkdyNV06Imk1w2v+1tr46qIUw0bt9w0NMpv1fzpRipMO9dsN1GmuZ3Uoir1hvj7R6wGQmTyQ
wHhwDDLIoPOPqvFBli3bGdAI8yuWzC9hdmrZezMkHGmiCdceHIqky//AfetT1RSQsYbs7xyP4LOz
iqCzsunRhCz8LNt6ynmqh9CPeoq50RVdMhPGOGn4gY+B3UmIyS3BUP4anGKv5QOxPfyyBpVZAcCq
qMj3u2/E7przaCmBmXysezwCTF1G0ELxhVk5uC0akJr633EFG782EUucsJ1IIY4fCOz3TUUiW4RR
xMZpc6dq3f4OXFDyN9OCLZLvwCy2qgAkgLEJa10bTwQ5xD9KRDnZ3gs0bfI2I/ErKDOVznM8vJYR
bijwh4m/Ivit+fcfeJK9cGGaHS3tsBBePwS8YcgU9Kh64+IzLgtIDcyEE9aDxqyRVRmdLowjghMF
c9aevmf9Bz4vQ4kD7PZ1PKQkvQpoALgUGirj7zVFuHF9dJh+V2HQv7Q5lPDfTdIbguMDvR/RsYa7
yYueLoJEos/n/ozjtZZvFZlnknFbHhjsd2rbKNlDInfPph4sCgKzO4/6A+JFavIStKlMBHmhzYSR
6zgxp9I163X0bWcK3TN8lUEoXNM1TFn/4pqnAWpCp812B0wB7Ely2+dqlT1GxMRkoDBKGoPewLdN
Lm4iS9REHGeckIVhAGWKABFKdiOTaiyeURnvizdtvMmGDfXIqI0JUxoPHyLqteKbN1Pvh+S30UXT
vhadRKcbrpKLMhPxzLJNhQHLWDuSxarKd6ykVDAiR83ZvQli6C/pu0p7xM6gmHqQjyE+dybtI6kN
Uug4HuCYvEnaARLjmvkODphzDjMxWj6tIcpkh+YLIcqnKWcm1xINHUmRJsmL6bHQuoU7ZA/pi9Ui
hcsCrf4zSuNrb1JrtsQ5UfK2vqT+gTLUOsV84oMbPlJcdYaGsfneQw7OGm89nSdd6bKL8WWaFw1h
aJLHvv6kC564zn7JmY3Okuoa4cqc8O0QNdiGNhGEFzxqPNC0c3dGfJwoeqa3w0pMZh7Bi5vTspkP
hJ9FIqfeMaV/k3qiDaNPlKIBn5rE4hW7hipivpdoshMFeBnINQsJi1CmCCuVpYqECaZdruG+m4al
GB1Z5hBhuMPcX9NivW6Ye4jLssmAHmR/YO9itRw/oj504RyrSI81W5+ShdZ2fVvyAiFcZZGN+nxG
TZlRGYaAVN/SxOUkYVjd/lA5teaR/Fk7K1+EYrSaqW2mNzK9s9HJXDYCLrUQVka35Tgw/3rdZXTA
N/kXdcdpiIPnhQdGrdROj45kxB0Z1oLUZ580qHTWgVGYOMuYyDu3goQ7OKeJmSa7f+N2dgmsKhq1
Lk3WlXO8q6rJu3NwsJc9zRlmTZWL4S2+k8VZCFCV4POwflSIXTKCb01uGbcEdPtxoQubNnLEgkyw
OzYOK05AOAj32MPKW+142pSOOrih67xRMiFnFU7CiuNaZhXQJR7+eflJTpDtQiIxoJ8QKxRznsPM
UqutRQM35wppqJYRhQgPzLQ5qOAXFoRvWtNICaTUYCCl4tz6UCXVUJeuj1c5tmkdFtkR+3AnArvs
ho4zZAnq7Zy3wTr4l96SSiiuHl5ZLNULIbCy41EpLxa38eGbtUHCugRCu/bGkPa1v9LugOF+ToOi
XCFlmivj4rwUfLyAefnp/+qKSIXyZfgzJZAXWadYE9e4kaNF1SJ8tzDXHs4d7aU5PrueXHsn/8MZ
GgpaPvlDeprv5lAU0q7+28bZAkRZfOLjeCAgvbPB9fo8lNrG1yoPh2tIqGTVWEMxAZLGGjnugfFC
kACHlctunWYtHJa9FPBRY/liH6z4+wGR9NWbeijgO7b1R4dByFeRBX8ABBRz/1cJ/72cBAMdqHIg
rD1HypX2BrNib7xZE3m6i+d8Q8UF/yRUei+GVbG9T/f5d3QYuIJw+l2255uiXRFsqiasmDUElD7f
J4ruaNO1OtXLwb4iNKQZW3juLsC/CViFljy4owHXaNxLeEOPzOu7bQinURsk/p7WXa6xtfon0ZuY
/uHYREzOuVge3sMQxa8FqVQqf/UG2zrvjcuaQCo2VfyO6RxdPl1KtlifBz8Xek9QNRku5iDUQ3gt
teIgKaYSv6/kAHs+nVPbJU3eF748fnq8aTlb5BdqJmUDEC4mb4fA20EkDn9knT9Ay9MEqYV+bKeR
fN2iSb2a3UfE/Of8k6Wf26e0YoWqFIOd6MtLzSy0Cc6Zp4OlzLQuTV1K1QPx17ic8Q40KisVW595
uGxl2+wjVKNlswCyUqOcirqUp1BaKPLSGe74Lb1wAVhQK7jLxwbkKRWJr4YlRaaxY3wiZcriKcJy
d4mJtlOGfXnH6/OIhZ48ZAOxsq466oy2Zl9Wf0jXeP/aq0TvbXQU8NfRmK6sFF037cj2DhUpL+Jx
R7fp7uY48rcfmpmdwpEDteA0l3YZkleFX3ZGIx1VqizvJ/wDuFRj2IO/jYBcX4fV3Bi5scdl5NTg
D4aYwfBypreJtYNxAxUsvld0CtvR1sUDPIgC968AIWdjbGcuPBJecc1aYNXxk9i81LPBmx3H2ehU
/66NCWHLj5MVfU92nsDj6oIulgNN+pEtj/Q57MuXECn7Lc4XuJXZdNBGmcx1qbialFiiWvN/AijH
p8aA0C+m/d46D5n6aaicK8Mv4HDbUv0Gm+MZXpNPkQSjw1SL5qAF8OFhqIWBAdMEfPIx+eLJjvSO
LUFkkGE8uft/UxgpE8Ah51E0a1aPLN5nbli4ooYr5R/uoGtyXk/wVJuZCEEXXGSz6Vg4iU7hs6E5
DWtb/MDnLlSkvFAO2t1JNB5W/+aLU/oXPKeTx46BBY6HVQvdYoV0/emJ/J8M/g4nvSBJKvWDVkYR
pWN4umgh0yKJ+H5RVSMtejZlgtp/1brQQSJA32Fjzakr7ztkOItArI73t4sPoO+aIhBavmAY+OI3
OAhBX1esNZwjW7NK1FOJTkEoJemkIIKMT86jqxj7w21/XCFDayMzjcYziwnHTMBYVEZa7/+HvDKd
Lj/DEvmBTArtkBudt9MlWD8TexhAC/k+yvX4Gld950zSk7Uwtit/PxTiZRCJBJZNrBN1fosYcoX9
66ybEVGn0+bLnLp4ysIPM3LpgRpq0xAqc8wU5r/t3IjlzXPnZAy0JFOcoGtUpZZUZwreowF1FDne
+8Of7vJSU4kz0rAbf8a71HnA5iBj+2Ha27xPC+YYUnuez17Ol3lRWe3ImTQEh/SPciNnwe8z6LMd
ocilLtmmyxelTNMAfvmnD2tdGtoI3NX5qvZw3C6WYWhPbLGUndlZyw7oPFRpeynG7C++ybHAYVZ2
HssxHOaddCz9d+Ayvz8a5294c3B9PBTVEokHSJdEM8VhnI9xUSakrYIR4LpNPQsOhfgjeftvZsCs
TOhIUeJCpGklCljNEIiBVVDRuJU8VNElzm5Zztc6n3eF7qoRD8U5/FvNIlDyzUXcOulvrKZvhdNb
jl5Xovzo0gmTCDE/s0Tf/9gc8hqXrc7V8A6UJdDZmoR86II2h6o/JUw0GMcKYmbA1Ho2IKWpTRF0
raC3kzp1l8fmvaxIZRAZVhzgHnuFMVwgMyRmw+EB78X3qEvhbsnp0S+a3S5iU2yr3hofcyRqNuTw
UAof0wKCoxZIBBGv2lmfgkHIzpEA6Ocm4ST/5dTqKTOibC7KsPUEl3KgzgPOVZ17H3K+hL4CgeS6
KFMP4B2I+ix0LJ9/aAIFckHhmNkmt1Phuu1vrpvmaTyTlOWzRZDKCNCR5BNyf9pNU8JRXL0cx1v5
wB6dVdRGX7Fc0/dMc/GBPEHK/OXPVSsQLyF75OG6thIAO3//OS5EXZnN83lQhNZrJPve6ycgn4Ns
Cyw5PSF/5uc6ssqYnD8C/FMgJopslOC91Xk4kE9KBWUDHMc1EzktAKSilHvPlIUgSwbOUYSrZMax
u7CAz2pIueoIbl+e9is6atpMBm/J2+DAvQntmgTw465yXWEHNsukgZNLIYQ1e49M4eZYEL2N1lFv
iAUosJHeyouAEqwZooG4ejQhgkMAjgEBXYtWr4i8E0ClUX9yd8hwx0l15CAZyBGuZJkw+2HV45QG
P6g+XmM8MRQ6r/NX/R0zH2/r1O6DWH9DlXs3X45T4eO6D/YhRAiziReATS/mNb5Cpz0E7IHWus3A
sZKKBI1lrqnexYsUnoihTfe1xlzpHOUEpS9tnRgv7NtZlMV8iRbYG3T9/YeluJaCVmt0DHgaP/QH
5YNDYFdNlGlri4eyqOk82nP67hQ7Xw8An3kQXrXHmcv0kgWhD6+DF+fZ9e4ghlxvld9qwLiAtUEM
vfd2OGK8/BPxeLrwVfbLQLDdOUyqLU9j1DsiXf0T0vXonqd+quLYethYUi4ZPGNJcIfqN9pIxfZq
X3WMFSBmAXRkRk2NZzGx9zwso450jaQ40MCnazA+FH6ybba3cLoxVZnXrxaypbNj3rXlt6VMRuk/
aG6rnICvwNwnO21DIZqPChPQFGFUgweNfRnfOixfKEHJDOV3MqXYcozRjW+74BegImMrvRa4YDIy
TGZGxfXAl6HNGxv1mS8nBXB+eMbZiNXDy2SH8oEEnU5INo2El3TO060RkwtLv9vvSbw1VBfgRITF
YeOoPol7IWBsrG3zrvgRH7qzYAUc9SwMxKi9H8RjoJSzXmGdyh4fyre2pRJ4BDygZ6tzZ8hHrrOF
AgtJ4iyEV68SYQA7OQ3sUBKIBJAy0aGnZdsb/DvwmosQ1+4VIOP6PnG4iHdytwvUgJtsuEhYqLHq
hwJTNMsfsEpytCKChOX/LxYfyoEAtsajdgxhIwiZ433M316zHOt1nN6IqOjjYP6W8Lt9apLuzwEb
06sR/oYK60PXnNexAFtgCYSzUGfL0+6D2fzoUJ0pZqk/z09mr3y0JNaK2KbA21TY2a9OAKSYkL3I
N5L3bG9N2hBQYdJLn+5LHcFc4moE1tFT6MO+jb8TofsFtEWi3xVQL5t6JI18Df1Lun2vuOml6xqa
HDe27JodkLZFIK5tNS9xLeJZpLAE4x/rn2mQIVI1L00n+ZT8myvv3cWBwxMAZ4Vbyt0oFVwog/j4
cDmI+L+jS+Ny6mS6RzbM5/3VOLUUMYy/ZBJmd2SvsanbijD0tXTTIQycOPGuBQlFyFTDWl9Ic9R4
PcfQLubrtvxc6vgrAB49YJQhlwpfAJjohwKU09yfKruGGNP979S7JLR4Qm0S0bpih8L+zrdzLlrG
9BgaQmpfc5cy+SbAuek5fvWMEbPLHzyODrXyz8W9aK1w617ubCRuu2WYrQtZFqjtOYHDZlC8irXL
l8gumjbSQ11LiJy40wQjmWjjx+k1GedZjx5FaF+HC0DjMDcwD5zGIqf60Zalh0jAaWsRsHz6Pi1w
vOauWoJ36imk5e1qFIb50IqL/XBoVE9iNQoVrvF0WhGXDscTUCFCoUhNVgJZizVXOLCeLjJTCFO8
iw1rw+IP3fSwMU/+PIbumezheFGsaNjAK9Hupd7IUA0reercFQ84cCWlLTqNk2bbMkZqfQvKpCTp
ajUBM3ntnnCVdoI2Q5qjWA1Si9IOSqXkbnXiriomO6ebhpjzjK7DHJnriwOS/uprEuJnYu/VqUnJ
VbBdh0cnuslUzvvBduMDpa09QCmRafbWrkYlD2HLa75HZm3PVAKbU1tHyP8b2zXi+oievV8/7BQI
JvCwA8mEIeg4FPI0vip68yzzNjc/FJlr+qVrzPOwhqYiEO9F/8357Tdh5XrcIAa/7HJm/J2IUHqf
7EO7uBUbzY4DTIudEC9k2BdUymYE/BZe/Wtm2PHSslsKeWk1Wn1KjDtoPgRqFCmYvjihwzaL+V1f
WirAdPcCz1Cj8RTE3bIXc7aJ3T8jO7xigr9AQKLuI4TTRNbo3cOnAH8/3SVB2fvRFA5hDuReir89
/0dXUvGcyICIUrvv8HoClRwXGL7fMkPDgJoJegyNXRHZtN4jf/OT+Omce6r9Kv6K2QLIgup0EqLS
u5+7DLG//gKoOTbgbEwgmgtABUdlxZzgs2FBta06bBey1krqCp8DKKu3lvwpu6W5BLSD1UrXpaQS
nKqXbHbn/owcVN8BLtMbbBQThH7hobBEqb1bTTU4LHV6SXff5g4cdOrYb0XI2/EcuKiyD//n2PW6
EkWeFmkNEKnCU0G2L34l6hCrsm1R81Ypco/X+11x/LjPbp21i3JMsKNRs1cZZDC93zO9cggpiuHh
9aDSTe9d9KQqEiHHZyZyx+S1oN2hkN9aHCpz4Rk1S/OdoepqlV8PI3myhLOhstq2+csItKMtjI4V
aNqJKPiZVDTtRcJSMfv4VKZKGR4PzcVKyEV5CWsSIL+KO8eYGxLSxjAlc3FDIvZHdlJY8XZLZ/MN
SybzSaowR8wC/KnZZLFo7CSH5gOKbYsuhwQ77xAfHnlMKLO7v7Mjt2uqJGfT0KNaX6dzfJ1uBm2t
LWfu4kODun52mrOisMJyS1gZ2e9vSL73tCIARwFGTFbP7ojJjAsLWnuSV2CC/NpK///BJ05VX4eE
2B1vZtGnzrQnEXqHYhwspNdoxKs1C6unsZzcQYbObrI9PYU/27rya1p/ovijdZLKYbRhbR9oNuFA
nv0kwfUOQUkdo9BQxiebs7aTG5zpuc72CxWyquy2GgvC1BevuJGawiwq+kIpPDC94u4uynBa4apI
mEBdRcUOfptG99RDedHm79Awzz/+Hcpv1Nu2Yjy/WjPQpFpDpwyIuBC4kilbjHdlqprPqs7YEBbA
5tofLKir9Mf0J6lHgZS9FTL5soycrOq5bXEOiH//5JuYEZXDM73YO42G1B8LhpO4Am1v9OOJRWSM
4Zbn3gvpMrPES5ohtCCT8qbfbsiNKI10i78P2MBBw0MiDYqBsBfgXtuEdO9MniQH/dpKB02ptFi6
4uPgM2tuqzqkhaAEnLOSpI7gAngbSvesTsAN2VL1t3sjgEi8DfwejGbxjsvW518ucb1XsUccn/7g
j01ig3FrsbZdIkkG+5nWanUFY/+LZHm/M7CD0Ko7E8hT5yhxq+HFsasSH9SoHJU5LHLC/V0AaSN7
QAaidmpRZDYYszx8oWM8C6EFzneH7bQu+0uaWXBnAp/SABRlqSrnsSbv93o8aE2oGDUeNE/AxpPF
/RaJAXphl3wbOx0gzYS99APTIJI0KQyaMKFOaSA6YMW2p9ZRdOocHqSiNMTdS3tjdn3tCJDE4l4x
WVaBHxp/jnCs4Higr5IzMTo5wAtkdIjJR86aeeUq43B7fA+Py9RBjUd4FlHivT2wPDY75zyK6I2p
NOxpdU5D0LLQnM8VQp5c79BvLwCz9giHOM/jOorrGaf7Q4GQ/tZW2bTDwfxPWuKJg0XVbrPFkFAL
P/B9HlNl2MijpNurBTGhHaUHqXv9Drfg2up4UL5Fz3apUBVbz1ZpKT2MmKEF8G6Xg2eNojiy6S5B
V6+TzKD7XldD8kcvUQN51rAMm2g3BdTlL4pgFtmw6VRnskIuSARvHzfFNflfdWgvp1ELEls7f7m7
pqDdbhsoRzjzdjoW2UaHr0c0QUq3RoUCeiuONf+/1CxwqL5K0RU76qbWAl7BxC8rde3620NVSMP1
B9AX8J42l1+17kqRspM090BjNSMyXbQxGdy/m7sgyPVB84eOq1On/gYk/TUpcJdFj7vVBd3OzBXq
bjnCxsMJloQnqWtrP+f4NGgWT5WcwOr+XE/JKLZDql3D/0W/jIed/8aYdNkh8cJLlb1A2BTb7faC
nz407eNc0PhS03QC0BuO80H8T2A1PEFtT7zg+GV1g8yp1YTdrjjM0l9cUhE6zFisYx4f+ie1sqRZ
mj1CrW8Uyyeu/viH+qOus0Ims4bVPSNTLTQbhVi/VtaE5l0WVzaT5Nf7lXkisn277YSxxJfN8duP
Dj0N03phmxBIrsW2VAFcEC2Ljder75Zs7waDBY9lZRxRP0Qmc3ABuq2FEuvogDA/CrdXuqrsWVy2
dJiYPOxP6fiH5fiMXM7GWIOiV06QkwoketM2wXvMQ43pZ3DoWs2bQgIbWw20YRptH0mGtic9ArCD
+3LorvQJdyFB9Lw7T40TfIqwdPJl5UEpD2C9TU2bZZvJlsPyEfbSz+MD2xFEdtWv6xc/TrsPA54v
f8xc8KQ8kh+/cDgep7YERp4psMxNMsUJsfp4dQ/9oHHlMvniu63mMQllMw2vtD9N6whglU4JkS8p
usmdtB0MUOthmCx+2bVAUbKljPeiWEt7uGwPXcUlKw+MnqNqfKln/EBKSSzgM6sRX5zarZ7ZVo5r
DJI+SCNtkXh73K3awXO9Q6zfow4Nqr19Jytp6+BBJ9QCudbktCo6kIuav2CMGbClrG71HUCSbirC
1tZP02u9KVveWVArsNQRFmoK6cGM03n/uaEpqfaeWW5lL/ZhaxgE9iH4w4JA0yV4Y/eQ+Ipl0tU9
4nnVO8t4s+vuD2ZUB2ijIL5qsv0cLuY2naFC2CGccqa2IcIVJm0kPHV2EhN70GoEW5hYmdujwxe0
xBqZBM0U1PIhLmWlSOdiE79fFEeNFoSvPIOVP+OhAJziyjVfEVKGXzjifSEU0t2WIlQd/eezL4bH
6x1gKh41m3IlsZeVDXt4AzPkkRFNCjr/rWhmcimvGtbkLpf29GqupXyK0rOPAYlDJTyXjB6aBnMX
RJsOl5GH7ZnMcNhhK5t+e9+DP5+yWKZyvRVenRi3VNBoyyPNsQ/7VXUZZhvRb1U6LXexqQNz2tJy
WsKyKQXT4tkufJaEsqn46ofTW4jl+StNRsJ0OANVWEsUIRu7jPk8GvGkdKoxWq+gl3piijjG1MRt
CyB9rAb7GZ9lhCDabrL5jNIg7OVH1Jm+Ckm1QJOnTgkfobdYLOXxmXRvqDfXXvFWqWSxX7R+wuTF
N+a3qdvgrxFvY3iG0NswZm35kuakQLsUVmAtQ0/xEXsqGSAQkWRLc7gQfdvLS9TMRfDoQ8EWPnEZ
rMweVrlOvPDeKO/LOQIiPUGmXGygYsWuzlH0dV+e5fLbspANAcZ8LmBhstYUxo13SowTym9AfFmC
2MJmoG0TMnWmdp6VFO9rxmRr8WSYeP61fgN9IQeQDUfNApX7KLbsRIRYH4U/QB+KUAmezHyFmio2
0/K6OhY6HBmdsuNpmi81Hw0jfGH885EXZhs8wFVaPMrNl7gwdy1AAXUVzdYFOwi9OpiNquDSxjm1
NgferH5XvQmr+zFGQtl5IDkK2suuUpxwyBYGlLXSQjSCPhlgdIyJdQIfesWjaUQ2vYHxwN7Px7Pz
1BPJLf0TQDL4gsNhUaWuQEFgoE/4Y7J67MwG5uAIHznK+X4EGLFQsfFj5J4ah396o+03VLaot4Km
Po/3GV483pUAxWTawXn+mSlPcPUKUIqeYp/1fLCn1tCIxtQhwjVn1+9VVJ7XfhSklBUT1u5dizEK
pVs8Hz37Dp4JFWmZkdRt+Ul7NHwjKli3N9LLnWHDFiDRTjfvzXjenCmdwBrg7FoW7BZLNqCEh+mw
E6qbPRWWghkFFcqoNQQBEFPxH07WDM7gAK29R5lRprNNor6JCCYaUjLxEuVKFHGYipBW4laMZ/lt
vdUnaLQeVi4R6FsMI8fhXZtE2Wcxk1PBAALOAWDd+yW/V1C6RFchLkPjsRxLxEUeeQ+uRfyXDhvN
2HyEc3gGmnKOOOHBYEIgOvx59KjQwng17Yl++CRyHlD+Erk10/enCRb0Xdc8ydTuTBmZraQWgoyy
m/kbvXNMShbx3ffw7Bwa0EyzFmVSuPpUhjvHPEzntxvlAxKRkNxW0McHaO/qr3FmJvG3NRyMDJiE
ajafQR8ERZw/lbv2Q6NvJBf7RO7+Bz6sPKejceBIFnGM94752C8K42sdKHv9H5gcrU6yV/HpaO4M
JA3iu6AAZNSeuXSdLYok1Tl0KYMKX8JTv/bKSuT5xNP+Jmf6H+1j0i6CSYIL5V6H6iS/aYw4HjQi
UqM+DtCBQwsUFFOmuJ6QtHOKwTmTE3zeLEua99NUtYRclqIYWdIIWnp1BpbhPUHWGv7j9f2gZElN
hVNO5+8CgTbY+pMFeaIB0wo20JxaFKIkt1YJJhVlqjt8YkxmqE+p03UmFRP0MPAKrzo5QyE0coDJ
LpdMoQgjqD3Jv6bs0dOAFPjoctAQnOXfQHalHLVM3uC5YtwnzYx7XnCZlk5mT8575gmpB4fM+uPq
8Ud/72ifESbEJIOqHCc6GL5vODUIB0w45mzUMFVzvloGwteR8PMa8io6gDgMCoq8da9SybZurTv2
EKaVc8U+3GIU/aV0mGTQkc+qGo8A1ar35hJhiLoUJJGJQ2hzTWmrWiQzGYbg3w9o4HlDGJ+v2+PD
E3lTRorTflNhS+jyxAqyQ4Bp0w/M4EtiNcLgxXAcl0axBAcyKncGvfYF3zNhK1ndlCFHvwZ63HDq
0KTHwUNUv9e40pbdc2/mcCW2fQ2V8m/4jB3aRR+/m6jSQCg8HJ0Tmy49cii6RBjBZil6gWLofkGU
E+90bVQKIrYmPofdxG6JqLtcuoaBYxiG5kymd9Dic+ILSasn7jz93pacJj/hbytOB7/+umlWNl3Q
IRedqcW+nYNR4uPmPBcCfTODPYCuEHX3mXi1VtCsaa/7gNXiGFIlv9qndMC3Hbz6anbO3EuLHMh0
VwtrRhblVmd/XNElxX6jhAv+1mvyaAPuceN9TjAm4qkVHpvv6F8L3vBWHfwIedo0f+N/3O5R4ZsB
5SMjewC6PnR1HP894pyyBbFz8yMNVrDCuhoYAdyf8COeowo7vbTTC0CIz4ERNinJiGnCwD/RasUo
pxzj0sbX98e9HxkzReCMgW1OxZGFHlqjdhh764KuOsmXd8bVbkv0DWe+njZSnAPGW0BXHY11xQPz
1ZDmNd3E9ZAU5wsDVgQ93otgpfeTuRqeN530XPgufH99yyBlSO3LAovbt3Ev5/7aL2NlA3N1JERX
Z8fuTik6OpNulMwAOuUese7rdyIeMWGsio9dFnO7p8IIxuAecFDVfP9nRO/1eqnV+vBNQ+DEfaVf
SA5D81GbMb3nMhvo2qBRUe7AysuUTCCbO0SNHhJ5QcJU8L1OBCm8EF0rpNES519xYZs2rhu8tGhI
L7b36uOiQ/35h59TEG+dih+wGjdHu+HNBE8iAWKHHTYv+Cv9BpPPjWRD246rBKDY1PaoN6RXcClc
RaMt1VdVTouTHIfPokcgqWHtjVzuT44tZn/fAkHWIElJ59a5fLnw8zQTMOeky8PM88RHqSd5V/+O
B6VN04xJm+iIQirnZFms7WmZbcKoWBewsPVcRQs71t+R18Tg9uIBfY7GtmMOD8MZRh5pJZYCvCbl
4QtZUfI+uT3GcPpKVsuR6TNyVqKOSPkucHrh0v7ifsDbTzzrdAfYVZZUXQi1XsUl2jQY9y815MTf
iFu27qIYURKScC/XsCIeZ0LoJCYMRnGE9W+fhrSISM1D6XuQtj6qU342apNMHZLyFdlZHr+mu0kq
IHCgIQ/GlIziaWicYncDISkYPjad2CukY7POYZeXET1xICM6HNxSbD5wKkNgT2+gkXJ4IGkchAx8
GhafX23376aixKfajaG1oc3lH9jy+qHDLXBkox9ocyfHk27hDvOqROL/h0poPj5V/JgNwIS9IJSq
qskKFV7E3c3n3pFJ54mrHpxwYk/Tnr1Vf84kpCvMq/0dISSyNJxvaUxMrcO0PySZnJWRMzxPreJF
02NxC6O6kTLFCauL0f0fiuUwPkMw2MVu6N6TK5R7ZJUrWMm8W3CdzRrsgCwXlgSH7gEcp/iKoMij
Ut52TTr0R7X26VD5AKNTrKKpXOXNZncFbjAx/Q16LXr9QwTXia9my27ui6QX07MM8JZ0pwe3WE8U
uFg0PSzwVMR/bNk8Kj6q57WnLZop+RaMz1oXuqsodN7Np3OH6VQsPCeSkZMReAp7x2FKtDzUpX/p
r+DhMA6iYqu2vl/39NQ12ml2z/qtOIqgsCGgqD5IkOibugd30yoEHyQZUXZNGq6kgGTqajldaO1A
+zpYZvko3LvcuzkT4Jl0tRzi9OeqUHlkpCOLuvyVAFtC//T4gUgPzoviNOWEucKUhHoRgqR/R1vB
7XS+VV30uaFOV0wAKDDosVCLNHAQfgiaPp2FTDL32qwPTIhc3hVpu6fgI9xc21KtKLG0txK5XTeC
Byw5uEV5V9V9bZj85n0FNaOIcXPL7f+iPVQhlQFvS2gP+Om1grM4Y5+ZfiQw7trqLR43cIWXtlQs
78ex5wd5WleHEGRqZ9iP2L8FfgjWWDlYkdl/So2fKRfDj6FPvTx/kF8LFzXglItp80jK6+doDKVW
I7s2KvNkoxyYoMJ1meFT9VSmKCzziXTKvdsFYbg9ejga9eUSJFVNb6Rr6sHDxw6UHb2Jco6iGawK
p1ccYE0pCKrdKDVqtKpuo8zFgaGJBrs1uZGTCNmoEdlgyJnb88K10Kr5IcUW3r2y8mUudKEJLqpZ
78DiTqQWK7WlzmH2s0dAlP7NjhAappl1NwRlzBBvYvWMXN5D4+cCHvdptuY4BNS08Jy1o6/4md2X
/7BkMvIRYGV3zsTTf0wnOVv5XNjac5Dk9fca6DMNFjEJgB3yznIFAgqobvCkCkV0Q1hfI8FNsUeN
Mg0Cz9kQIt0G1sgiVoueIP0itM1yMG6dhQoS57pg7YLEB2xVVwAIc3r4o9nRt9gQkKWkRVjeQdPp
qCwuAJ7chQavy+RsgcPpZQ/iQdSEgDh2Rp6qYvCGWLHQwsR02GIdS0/k2cnIntB0K96eL/Orutup
147LqPqFLSxooMs2C8EwcmKUi8+7iRXOFIJWLrZZnkaV1n/6RP1+5QTMVGx9n8kxnQ3IN+d3UXnP
4XApHSlknvUilEy0a4Gs/SYJ6iWXuBHI6fRsnFRVY7X53lxVcNi2vgRZdNfDMjWIN2+SSXQiBDI0
EOKh9Rbb+PYBYVVtnsh/q45IR76x+YLlRlVMyJR5K5ylKvqJmaXpVuE7bKAwLXGq3uDEY4xTx4AY
R34sk8bgsoyaQ9OcfTakZfG+wVFqB0973KDXpzwDGbN/9JB1Qnfb98oDf2MYve0YfeJ5dhtBP3Jc
r8yFaDC+rU8kMLX2jZW/Su+gZ1lvUTTzHWc6Mt+8DbIi25MixCp1GheuHix9COnDE9R6g7dow0d9
gNgswZuGNg03Z5MTgwxDEjNCnxflBP/4eNZrp08RQqDA60JG8MBBiQqS5eX4cS1c6y0alh0APvwK
pLVkwrNTdwlwt4C8VKZM4GLBsL2TRbHXt4P/zscGgCU6IHbP/T/1on89UbMeZawdUkurOThUEgii
QqrIxjGM4Mp/dIneqJ2bbMpSCj0tu1YNdccA84CA6D/vbaAZjWo9MQafBmVd7tEU67+XuiX4FkW0
utZS3qsvX0wkZAUVCXOgnZ987CGtDnUErROX+kqtdUDjnOS/ovni9NBs22CQRgFBgyjww4yGg9cF
622RJRqpPTIdE0OkKrJR406QDX2p1LWClzcvhHP+5wuyXw8nurlbHOE0qiMbsjSClvSXi+diE9HM
jaQN8Ptc3lCUfGx3y5P19CWvT69HPfSpGLrNVAhbtJA5h0LetWoNCQL+Uw2aEbuBkzj4wdpk3HvL
Fmo1qguIyggmvcWokBULxctJUzINO9SXDXoh5dtsOxK+ZXMdcCWvuiahN+XA11KUEbtibTw94VNv
K4V92fZXqhew3dmD0XN29C08OJWPu5f7LKo7qigvxUFi8rS0Z7uxMOV4tP3f6K2RtR5hssmYpyVL
j24tWQ9xI6mwsIF1gEnkK5ER5vj4omYndWC7QwJSM2JiW9GvQ5MS9QCoAsCxH2bEJzLvZ9rDFqyn
yzuOz5h24wMKT2l/o7XyC3FXnDenMXjdgjrKh49lumhdcPND0EAA7n7Eg1oV7uEkTAEAWqr7nkc6
n61slhxjCAEksE23wQRaBRLX9sfN/nXooHIfDrNtms+5GJQ9TVsg7dOhxvARq3grLP0+x78M4Kxp
BGQbfoLJbd22cQucFT3oq+IKGKn32WpY3JX/4hAukKqzmvieFkETiIsFifvtPsByzZ4ozaE9fqb+
kqxKwRJxV9OLrU06M029M0b8RLUNxRmPdO8Sb3YvToRvDCqBJBkc4GL/cpRT0KTuD+zMQa96fnJb
K0JPypKaI9XOmjP4GBRsmD4uDUBBTJWXlBk8zGmYFmxa8ZPbiajnne89LiuLChnjusFb0W+1rSFe
c1Jc2JAa6YjgeRxDRsG/qpxiYPyYNpqeq1Wyf/tLTI1b2qv80bza2ITFs+WDwJRPqbHoQOgwcxCP
0Ynv+VBEiKZ9iEIKqDk/Pcn8PHMt9xa7obFMy07uE/tgyoO4x2tL28lDAc/wOz82JB54b9W+zc94
gwBze8hmGldZyjsb8ZXIctnObbyXACr3zNMLt9yxEjxCblI0r1ibi6K/wxU2WxeqJXuTFVkNrwd5
Qjc4Kte0q7y0wbOld8P66E/8XVf8sms2J2AZEpAztMpkHWiWLi92+dHH5Orc+6LQAAjCgazTw8gI
x2YzO7viyxrTXWi017UuwtU2HVtzYXSbCjAc+YoYlW6eaevz7LDGOJqYZV5VGzUWmqQMRLNRv2Hs
4Piuu7aki/Cf4py1EbtDISXM6FH7ZTIT4itTMLxKQ25FPdDJqbK3rWpMs/6nGHdSJuYShCIRhBM5
yrcPxIs3mo0ZVfVrz3L+U9nPyB2/UJaWA9/F9fb6jsdKeBH+Vy7smzc0wVRBMXnvDdwtFRcSXYCf
R2P+9zKgo5hhlMqclRTlDaLuAJyIluA+okkf3gC5Zj/FY5f6hKYeyNUqG+Ibk9aqWwp3mPWDMZW/
TBiQr4VYTz6PBlZ/tpVoAHtaru+zRlYVDiTcpE7vGepxnddr3QhAMxBfAWoUD2dTeDddc8wL9Y62
SqxfMKzz/yavmXAJaxQGc/W93MecJynbnvXc8i4xCohShGpNkGZtgHnJhZOqqa/gmiv8ueZBrTx/
/jsT+3vKeLLu1+T2DVqgzUVcRHy3xnCvdi8Anz3Z8lvi7O1zMvR+vAyA0sz9XQwpAEFIpUQqbI9i
fLG3e26nOLroCc2btbm3B6SpKNAQmGsbCREhCOT2BubzEAb8K4LG/Vi7vOI1k9yGXk/DYOo0QUQR
CeQArvAoJTnFGP0z2lVgYBbJ+gEvNtKHb2OYFh1TyEQxTQySsA5ejfUiZwWD3ZoM7UG48CNujM8Y
qnA8tp+LZjefzfSEOqFXSCpNHnujaP1jtG1AGoMLCl3WdI51k92C+FrGg0nUkzYVt18n/1Ol3l3Z
wxO4mya5KbBw2rC99+fnCHEuJM9i5wipX02LkAECSbXquz67Rsd9piRfhgRfECFdzVxnPSoZxk+r
2Vv/Px3JNwpmljd9CxqL6WTCvqG3W9NwU9Zvkxbvde5098Aav+0rZ0vSTBOLwqXhwqHELeLBndNZ
u2YTJv50o1S65gM70iBVois+pyJvQfd9mXxMAgD90Azl7fADN2J+2hDY6AFiZ3+kDr/eTcRANmgo
t3YKRDmONqWQlq7biln6h5iTM79ppg3tlZcm/KC1tK6CqAkPdbcQcG1XByz3xJ4wS9nA+RMYPjXc
l6jzVJ1nUlWvz3gqv8umEpSzL32ACC480pmWLCoGvqyxapgJFbNjw7ftitPCb4miuSiSAfNUBKv3
qhrx+Wa2OruEsHQm+Yb1NSowK/+8N4b6dgEFFZUnHVAcUze7DWGo2K0xPZv7fZ5jIn5jyxWmtE76
9YV/7wFUdlc1wCzY8KK+K8rqK/clk4umqB7P2H50NcSykzHh79sGqSJqYhZL4cKvRbu5wJnWPyLp
iow2zFiliaDQP/yRuy8x7xR5asILWos65jUgcLXQ1/fdn4lvTdNBhwlyux4UBi84Tc3mquSVo+y1
1zOpGktuFm0f+HcSX+uhmLBI3qeAA6+qJbmG6mhZw9jtpWFyZM5YYKe8awmudNN0t1V8IqZeKGGE
R/8mI0weyg+u+PbDa/90V+Df6m7ZoTTTA2DZdNoK/vwsBAJzqg1OBPvVgQJwSZaJ0bquZ2unr/wV
rIz5gwcpeHc58OAkOBv5ilV4TtbEfdjCrqHWX5bN9yHOElPvND1jvWeFhsOnl7nWxYeMJcG+Xowk
tA7uIRiVC+cqM6MqvPEN00drjvniaOCrTv3B13DVAq4qAM2Xh3aq0ZntTM19hxQ8JcWRBFTjKuTu
93oT8mO47Z8SpBgc8+GQOL4cX/Lp0H01f7RpSaZPpJkan/WWLrttFsZ4oGeAfMsszP03hdljK6c+
9/MuXjtacWrHzrWthai3+j01TbuIER5iymCRFkUl4ig3gT+NHxGtnaY0BzNIsSXFEyvA67XbkF+g
qBLBfprt0kkUBuwZGZypeSvkbEopdiLeTkKgF16M40K1fRLzqXJwXCDJ8eQ414nHC7sMkAgHStKQ
oD+VMtJdXh8feAcxRYJInGJRWSPi1a/wsyVij8nhx+x8GYidWsS5uDzFuvPuwtXK4+ROfU93dLxG
3fA0JBVxr13/Y6DhZVRteuXcugJYaxbCE2qxuZ1lrG72DxorFwKIcA2iPL4ojZSdqdcO6kt5IK7Y
LMIlc31NZUgkU2yzf5yGJAoF6ZotQTnxQ6ZUvfYz2wjERmDOfsGViI2MaCy1gXgSdW4xIJIh0bci
5n4pEvjvuIsbQncFQlGr3UFoE1KSYqHl4OOte+uKfakzUwPspe29ESbPN1INl6aauo+ectawW3mq
JjMGPeQ/kPi6sS4fWVdWPrWRVmrwX5AYrCYHffeEO0948PWbsbPRTKEH8f1pZ3gfkkHVkb3xk7lV
vHfd/lZ+lV+owGWyPPBGHmaVuYyDuiAfrGIZwGgX0D1vfUoet67Imt35UIT4iVKt72a4kYYROnV4
TrGPsKRl6bzK0WAoiVr5Oyi0mXM0QSv1XbpyRZ33G7PsdPgr93xuFvv0IABSG++qZ1YB8ox2/v0q
rYXbGEPzanbMYA2BTGIsDys/pkBO931HKf4A93dCFMQlEHeo5iEZZYg4ivO+IHnvebZQiRaWOh5M
AjWTNR9JLxdpxsCcn9bmWyNYioAt0UaVGuyjPJzwgxVkzKNZsM9N7Fll3qsOwpG0QyN39PB19uEJ
zPFhKWLETkJjCPfyCUaKse1BwYDS/dYlJwlFu3yPgQuvEcot1VIZALGf/+pp8CXW5gSvjixsr6Wm
JHsI/sijJWy3qVbt2jJPjnfIDCAAhcGl8xlEt9iNEXk179GZ1JDWiRLEW8XAlS0UjEiUa5jzIlma
J0JbOXVSQ4dz44iNdizwN+OCtMwl/Pg6kQXoPY2b943hWW0YeZwKIyY6VvrkqsSmziE1sB3cuY3K
Rjsk79Yawskw//Cqzx21140I+SNadAZHuHRlOOEnktlRqSkUk6UxrPxeUGbVi9JkhS7XQBAzngPq
TgtP5QZzjfN4bRO7+kstMUtjJWZ67PkK/KbJjQa5/qf/aDesBNPqX9DqzgVOyvpRMxGVktPbGwXd
p1SgSmnwKKHtEiWDjU6at0W8freTxmH50THuuxjxPeugo9ypDnr3n5Xwgippe8VQxNDXKkfdORfn
qEogwawN7s9N+xmv8BCaaczk2lwLt7oMKJ1g/aNTYxqkGW2lrIwU9cO2J1lzYsW6/HcevyMlwtVS
3X0jsp7dWbwy1uj9FaUqoC6XAEOzJfQhFfzG/4pm5VcHXq7VnI1oXsj2p/KxMzsQwxvFHRRn7cVA
HMdFMFqM7G0JLcphNgD6Oy9Ot5zxVXwj3s9PFoB+c5bRNmEvs9Ff2cUKPXHoY12ldBAul0LYNo0k
8COfvHX/6bR87f9uQmCObus2s3ognPfcNV5sFrlivi55aBCyPgufS14693Uv1bzj+8fYFh6JQUl9
jNcoXB5KiSUl+GXnLWUcuN6Xr9s9iWcE/aX+Q5F/l954Fh2FYKP7yyd7gLW0wB2j0AteEfWp6vtg
nC6GlyzF/89GsYk7pv1OltZHlZE1+cgkEDUga4sL3SRI7Igp/6yHjOqhwplCeOdpDzYNN/EiLPel
Pe450xDxo4vayB7/PDexPevNxucIRStfveYNO+IX+8OI4BLxFB/LT4IMOzkxkyvrYujHTnZoXv9D
SIT1Dc6j30OLqx717Bs7oYU5HtfEsqC3RQ7yrjabBue9xcQ8IgBsrFtSE1DG4INjAe5GRHnvwA9R
iUNnnBndTwxSd2Ax60dqzcMK/7n8Vc1CXxS4J7pXWFSEoJlvYupyfMqxjF7nUo31y0pfzPIGcyDy
7SEssmtWvGJheorKxuDZhwJ2qWtGurFxDqmu6DqfCtkm7S6OmIOl7aspIxhBiKpzCdTqiZn6E3g9
mCJRU9l4xpjhqtufWVsHV/PIJ6EpM7du/bTwC7ZFSN7DgDfBR2Xax61d+c/VqW5R1csWYsbtY6cY
IEKF7QJo6gD6tWGkFLm68IkBy4nv8zg7gxDJEZkdm8P5qRwtp0BodA/bj9kc/2khB7YcKzMu4AsJ
ozEOo7vBXlxXzW0KeTrPwRqdwmiXEWofU8eLCFK9yK9uIUzg1Mho74yuylLRu5g6huVH1xreZOrc
zCum3j6+N2ETw/MTHm/xyFa2l6A666/3Jjxo/bFo2caI2UAF6A2kVQ8CLMFa0uESwwEw81+2qjbn
Aws9vW7p7EJX5zzo/idEHCimaLpsEmFoNpCmTops7UaaEc8D5LbR110wzWzNAuw0iHFac8EQb0N+
jH1oqcatD+kK0YLJlNyOsNJTiLQuqaapAqSPfEtGlzK4Vhki77OLNhShb5CTAMMTKCxNm3Qi+Hk3
t+BFA3xQ5RjJH0Ff1Has1/nkXvFQBMuDWvUSIC1B1X9/cpl/gbjSz7OAFbKKU22NmLEyFW/FSQCl
TZHjP59rlRJ2+vv/du/xwUf9Fb9LMfPXt5lrawUiMUxjyCuFJHFqeipanJAZGLORdoYVWNGADo8v
1hLabGulMqdWAL6zMs45lhWPtifPkSDOfOZUAFqGZAXEW8pwxtTKuumM7Knz+TWs/34rSxUrVwPO
f59eKqT1EijMmoAp1tZ9Qw/SFzva8wh3KqcMQsDbZyEjCZ+l99Ee5DOh90fzr/b9pFWANj445YsS
CUfIBuJfeOsh0Wr5w54qdSrVywIMzktNXzdAXI7WemGSxVA85hOHmyHYE92ny6oTlvrR5Gzr46s4
chweY4GIBhWpgEAaYLU1paWAN+P/wQRfJRoGzF6IzhyO4nlFFVLMxIfvA+rG6xRylR422x9ntHwu
4QFLZFyoPmYh87KFv5Tk9OK95vy868+/dt9zoPiDc4Ew29PYQkwInJw34WAU++EXZF2Jx73pDIsW
t1h0HWJ6PvGIquuezOWkrIbfkYhKiqkSzSABHALIAO6OBkhJGQeZbQPrOjwW4WwMy35/9X6AAnmx
3hTX7DiznFgNFA5MK4GgikgCVgIM1JaPvP33hzZlwkwWMHjw6WqhNspPq68uFoHeVmE/wp3fpPjS
QLQwtBHgE5of8kVYbDPi61EKsucPI9P9SwX/gqeSSm8JCb4wywqSfqH0xgX1nfq0mGdw7s8zOXmp
ffO7nB05DQgkh91GMb/4Pp2NUqUIroOmJrwWdzZMUJNUtL6Id+WKLDWuHMvuZrZimoIZifd9tJE1
xCV9ZYQDNc1QbYipGtK3pdTHLfK6OAFdz++RPx186uk77pDBOJgmZhUf28KerqGTMEnXVNeE+IDP
b6hrX+/Hnnk+l3fUHn6NwAKatJIBJ9JTudP5gMWBF+ZOU0LIP+wnK2stI2xcvurWlMnEPc7OYgEA
IlN0+5YBcgqKdNWv3FplqNoKi5zQefxEi8SqXzFydGnsrDuqvfto7CAAbYIPlwWpnszxWyYpfdtp
a2rahDT0kSTVzutNojMwkp3duLf2w/ar51/Ln0ftZkm1fee44dvK6TnnLc4mH54SnPJxtjuyn/Cs
nggzI9xXfBhY00tAAMcEAEje1zK8cS5lQjgSifGl7gipzXz2Ru0LpPgoP0p5om9kdixUzDt47OWV
V5fwnnIJfANu5QayYExh8PPeISJ57Gi4CT8UHs+uIZUO40ceyO8tm+KtPgecqJp4tmxsxSHrseKN
wfkREFpcBJEPdUXgE75iQytbGQZKS3WZrIC02+5w5uQZ6xLPUneWKFC1HoFpHhCbBJCsLGjvkY1h
/beoYhqSksyy7K97MSDn77Lo4TzBPb9u2dkLMaHjnRztguCtpo2G78eUn2pvL6Io/mqTfkCm28Sw
yKbhcENLHsE/XTbN+EQ+jiZ7JorulvR5CFn+2YUH9ypeSGqKbhG+SITP/kUhIUTORtCttzVao9lS
Vl7T/v+zCK2t8imXCuULrTiovec3fhkw13LglqbTeDHs4x0IfuWRwk3QTwJiyjzrhyYrW3ajpr3D
RK6WnEfVbmltGtYbp5huym27qSLUhZ8RWX63/wZamis8slIUvBGEJDXxQLaZ6dRGN5xc6/xuzUxq
ZIj2z/ampSCiUhbx2d+QbowSfBb1tuBbNmmVz4IVSmc/kG+V8ovH3bzxURpSzyAjcPxzgwBFIVV2
3tGurnOtmAqbmsjzFZw1Yw2aA0m5eC78wLAu+wKKtm7kI7bIyQ/SIJfCukGZcHzE8JQ0SDG5F/87
reBa+kspmju2pqRLU681lOZ4xqs9TcM6PuKTky8zz0H0xKCKXFpH8AOqmc6wcc2S+xVSJwS2C0jn
eiamlUAmuYB0lvgEx15eEV2sbYWHrG6z1cheaPxHh4guX6MLfZjdZ/l8CH0F9LT10UatS68YjYBw
MxH0/YdqCIYZGQmGX5i5LVr4BQosbry0tmQ0g0meNckGtbWRln5BWur/DqP0qlHFeB/Xo4UUCTnw
B3UutKwSkktWLsPJRvEHO9spjcaOmNELjZW3WO3l+JQQJ/I5kWfBZqu/rvCPjB/SyOukusvnVh9t
1tr5nVnrg0R2RP0OWJNDEUx3GiIa9Y/iMoAx9nnREdohTGecYfLB1VOlAxwJOAbSD6hTzxu32mrs
rKQlSYJKs03nThCdQARCH0vvnbVfhSNf+ZmRv1SaZ/l06LMhEki2IpVvl3T08Xgd02BG2gbdTqyS
mDsjUecgZx70M4XMmW7q57apl0zrugABAlFDMQd6EvRZYSjJITUlOFdtYn8TMP/nzCbXnh+Ombqm
CoNx97UJE78EBK7+/24QBZuaJwZFqP1udz0piKw2d44bCZwjaR/tPGKqiTKpqTOv6/OPU2HYXl1G
9CuPE8LjPR4NLSLRJIsq8sg9HkWFtY8MMOlUlpOpvz4zi0eNxN8dVKSc1V0sWTlE/a7iUjhLWsRo
UT/CfAL1Z+cvmDdl1VlzmNh+rcPhWEPtcOU2vH/v6Akg9Gpwim0VwVjk4n+mIHVoP12V/GpQ9ZLY
Kvn4IdfUokkAETLt0WhiJ/JgTPmK/4j2qAE1ThdqZdtOvRpnqQCrDV4eBBvFWQzJ4B8C66XDN5h1
W/ODmd+biX+/6DjQ9Ue/fdBUxTFK29WJuFOzkHlm6jARQQshZgxzT8z3fryhlLxYz0+J1E/r/rAL
C7wp69dA7x50NW/QBi03/Uwc/iHx7RAlzwJC+wgHhYnsYV5b++JiGN/ZrYFtPGQ78g2u9JlGKTRZ
Piv/2OSzroQ6guIsRIy+hPIArzopIvgR9ZpbYObCdfrGs3YktRsbDmeqtYhB4MRGZgomUemedb9W
5zS5xVb1E5IyBqbgdJyZ1oSxNXODv0UwEF81RZD/dQQKdx1/QJqcVWRR8BEf6axpbQUPj8UsKcdF
9+vr/c25Be5FG8A3BWf48aUDPfF42fgOdAG2otRFMHZ9QLyMqBQ/8RplwqmURdzjsT+7i/xvbfuy
I4ljF7Dx7BAdDel/sYlFng0yLa5zrgh+wA18MzUf092vBJr3xPzMslRnukdMd5WS/J8MceJx8D9B
G+hddyrS6hVpLbRKXcnWAG8KMDkyCQKVW554DBGl5ahEyPcAdsERRDaG6K56Qi2JUeoT8tvksDaa
fHRUeTei6Uchpvoku2V7iB31K+dbqUCUtTHOucoAsqFD2RJh5X/XDJlPZQ08it9LqwuHUxq6/0q3
/SviSP4hoiLDtD7SQy7WGr7y1Wz73YZRzWTZtEhy8WgdLRGfOgHTy4RljI+SFGbm0lQWNPIT28r6
vjdNkTNI7rYsPdZLRkDPU0IuKdvsEwv6WalbgIclMkrsYIiPbzVJhNiNhVQFLhYJHfJWi619LB1k
VMnonq2MdTyJIh6trlm1BLHDVRljjCg4AIHpv3CtXkOzkNoEunbQKbG6U1OJnI/ALfeyfnCloYHe
7rVc5CI01zYkvIGulkr4EY/HrJbwO0NXXgoD+uzs7Gg0jxeCXgM9nMm9ikrfUucq/LfAf4mixy/a
h5ls5x3vfcaWDbpaYubm0Al2eUcDlH3cj+DB5j/Mm3HFzbotxr8yRHgKMJ/OxwrZFT4XLnOUhDTl
BwCu/Sb8ecW2dFkPFQB8seNZ4x/7xXnr7GvEYKvB8u05z9G6HdDIZU8UzMPa5vhB8whvJ9QftjnW
SUa2cm+o6htC9jOZuzjbmMKwCifwlFjXW8JhL584/QaGZ4+LYAaeOUbQHy3tadD7wzEEUIPlqoUu
NKKCZS2E/2OrbEucwGKaGoJMcTK1qWMGPCFOMsBuPhgvpwzR62eIb7jM2Ek1iP37URBgzuExOqQD
qCYmK5KJnZMQICqjPREv8QJCwN7TrKGcbAIBD4KtI3Xx8idihvXAUqxACV45LnswCuHXS4svB0XO
Wq/+DHGbkzZ4LuYfX/9pdwzXAIFvr5WIYjLvHOjwtMqkIqWqpb7dYT2WfrMR14FR/Qr+8E16Y2ut
OYvV/FH/JXiuL5pjkLkGdxFl1zO3u4rsASxo6DLCuQNVSMofkzHlr1P0f7D+qo346Gfcb2CAAaow
ZeVS/+7KF9CVkKQyOORZ74TetpNWA7GzeZKyhSL/1/GiXyuU/wTnPazrUXVha0rY0kbWsnLicC6l
5ZzswAdj2Xzo/R3LpHc3MhyRg4qTk/oR5+cNen+iTnkPeE/a/z5Nd7Z1jg3hbCj6+B0sy4+/l0JD
MUCiMUVBZItdcyj1v7T9en54DKB9pLb5nDWGUdjagx0fjRmdf6WHLNXccYV3rB5Urml5W8PTRJEg
awJAaJbCyGA0QJVoTEZ7vq/2UTXv1oCDn7reDaL+cEwLlmZZizv2kpOGCCV01CqWFKIROOJNvt9+
5u2ljMLPvPEHyaevbv/pBfznCFtifuhLa4tl5pec4fWpdBI55nm8mmjECKUBUstBjxknS9Xs6gcW
0eTSGMrCJQ1QrjMy68Er9Tp4wXE0/p5q7nLwdO9rtiwzz8guhSBy0phyBLs1ALPT4fN6HuUhagxc
HRPBwfZ96iBrNEWpg1NBHQLlN58G1oMfXHPpWOeJQlrPua09ROVt6Gwso+vQX69xUuECrmoFcyNQ
SzmRO5SrEwAM4SRA7W5s8gWj/w6rmYycp8af1LojSVOq9nBfJy0YWiI4Tsc31xL3JCAhcumccc5o
22XbTg9QHYOINThrsKKFtZJ5xJHSpnYmaXoLEmwbqwGv3Yg4CjqKX8pjtxJV9JbmuHUm1nn4Ip8g
piEyuDlFxgGZ2T7iAiWy5AiMg6Xw17pWLvRIEuYl+++qkWlGQkYhJX0nBjF4vEbQ7HNeJ42N2Kk1
VTmDlmA5HTAlS8NzK0SttKEFY0MS3vFGXcZBeITZ8B1ho2zwnxIlQWUNj2tCs9CvaHHHcKppz2FG
8nugXTeyNv1Qk0my5pVA7+1AfljVKVe9wtUrR7/HmElwMKsHHH4wrrzL/PTpbOMfqohfo+7NqT05
3+81NF+YYwOJ/8bgxuzNHBvon88I+jTZi0SKmN3i+SSBJ/O5VnpCgdJZTaV5OoY75iR2+PbAJPIr
a6sAEUYmXtH3oV6lDf2tlEeBqsabvHZqD2VyBcFGla3SCMF+D6lVWtJpbggVSYfFbgtBjIQfU8oX
DzH5kCZzMvFfF4mbU2oKvkEOF5qGExuqIsAEy5UGnlq9j+WWXUtH8szjKhybTokrYE3/DeBg/n5a
aWANhyJ8FCVO1EfBkpexRf1MdpFJGjUZl5z5hWeFwOZbxHDh5ZJS1ExhCojllPHidIXoqgGiQRLS
qi18IJDZLba3vaq65MKmo5/QQ2kAxizGjz0EBvfah2EhY3DWYf5U0rWDecDaRXGWIDAb/gL9Rvg2
Z9LbgFVjzmVGWXNEq+H7PauQxTNLUfmbo6HRW8YnLriVB/o6DTNWcbtyVHUP6TQ9EvtC8WZI6WUa
3C2U/ZUMCCz67aBNXRCbdJdzFRRBxCkDB+/FkTCfddgK8vPiuemxSM11lxyocfjnlzKPzynIagHS
gw5cnMsXv4ZcYzLuZSHCkxSfSAZ/b/K9Mk8cqv7zvHVvZBIvdI7m1bNhpMp9AsmLqlrhZZ3ODcuL
r+6skl18+TjTVkV5Pc/IF8a5c6JRGYW9GGRhZJF2JeRX0qCOHgaw7IK9NurxH2j+6SvdJ0azDspV
+sReFGHr/bZSTJkwHm0fBWSkvT7wS6IjjbpNR428QfRB12GxtDHawnXx0rlpZH1pZK8RtfV/4AfN
exHLeDIi0fcBVnPXqOcwh82vjchovJZkIqGSfvfI8tNBFV+X/Kjzy+AxIHxAfIGLMeh4DMPefWin
QSpTRCabvwG69FzuvuFbyoBT9+ThNWfMwiinEn4wOSzsbP64jwm2W0Mh7QjmYFK7A/ldHnibd3c1
NtPgR13xkRQUEOHjcL4X6Vu54QU5DwyA98djSZH1D6INlGgpxHWqAqWTvp9PrWD2FcR7sotStQFZ
DD43NjW2PLBLGfFkUMKUAh08UbRUAMt03daAWVg2kA/7Bm7/7ibktvaS02gxFFyagmDZcAHv+RxU
+3XvZgf8x2X48WEFbzlzKDqJh20yISZY99zhAH3qSsnruHHu8xRn7ieyH/H2QbrSZmCtKKEUs37h
5N9N4tNsIyWo5A0lg5dO87Y6ns/fBYslw+nsFD7bCbcy1QErErB5ul8+DjHB2JdNjnk5IUsAlAiT
z3x+h8nX/JtFTiFZWkY0HKjvWKf2MYjgI2Eh6OWMFvEt2JCWYNxR83ogMCweJSdtoN3HCzkKo7HG
3Y7UXveLJtuuJnUAcMYN8xObTfN2crk8AU3xW2HBYz0TDnwX458wRlkWAEFqVIX4uDhCyowSvbew
0WY4WxJ+na6+1JooTxfZVoGU99dWhaIZpexsWvlScoqV3WUh9h06rer/o7W3jT1iLan5rRTJWIui
WN06Fn3MUAvhjIBPqNujPd1tLomFAPKnb7+ZaaiyFVd3uobvUup9xFwXztELzOG4DS8TITJ/L5u+
jpJYNlPLtqxUsS0Y8zx5DnS2ULKGT+r6kHqaLsWwg0gFeeQHDuVKicmO/Hhf8hX9AhWFxEvBNJzP
5cmAtIbVGpGzJICHL78y/+HfUUYW+0+DgRU6OALszIjvo/XM5Av61h9kVsq0sSlP4KVGXl+r5Gi3
FISxYgCffjSTtK1+jEkGayMDeDT3EWCxkx4NxHFezY53RtBe1vjcOcF/gaMdTymh6UIriM/l7x9n
Oukw5cfCvdPoUc9befSprwFwCfyhzr3u/YBiMYx/ZlRuDrAd+64C7eaq2QLUUAifMy8e2Jq28YPq
IRhql61kdZP98CggS2p9fHa5wswEtip4eVLmW+4lm5isxmQZHk0sT4GT8t53/hV4ZYgopy8H8Sot
Q7X/fvQFDh+Nmw7yCHK+wSjcPb9EgmSyM7xQ5V6C1Uj21kaoKJ+gsBrjYu0QNOrq4mYtMxGAtD7r
Pnb9UPUJccpaPqqFM0rVXJHkXpjqFwy+h0xCNm+I4WwslJ5SEdvFUijf4ndWm76HIX6Br3fKUvEV
IvzCJZgOVDPAzRruu2elRePKKl6F53a0/H0SO1uCYAjFY4bIVYbWpb070C+pN/dSSfvi7S1JsZjz
22CUfcJ6Ulc2Qdq6d5p7FNdSPmnTSOzlih6OPYVPcERRlihgPFO977tX0wNp3U5uJNo7+3KsCjmo
qUhxEOqgZwGPiV1By0u0Pbth1jcdsTdP2IMdcWO0bAuYsQmvWwwqCzQDGRrbgGhhZjy7a+5Px72A
UDIcgjKiAYeXwXkbyz196d76P/Tww7NrAbbT/OlW0ePcY4him3HSzyVY74aNrMvP7WtdE+P7sQQQ
OZvcUJLl1meXPTxoMMqfra7VY5H+EyJrRUmXPSn4iOADF+VNVJsn3G77MQszbBKGej/e7e2ieeM5
yA1QUoZKLd7xwcfPwQXAPqQAcU51ibXQLSVzwZFbAeQedbKUXtyo+HeSphq5tUcJTED0mJ/zdY5p
FpHIIwCriXL8qr3vzhtwW80Q4RH7IygePRT7Ab+PQhcVaT6N4oAAluzGpcykuIsJi6h6Up1nkVbl
q139pZFVHooviNzusp1OxbDC9OVqidJcwY7g3DUHpOUPnK4KpK6xSqtNofSOnpwF0/OIE9MOsqVV
XYS9U9q9JwsKHYv8Y0S3dzPoaFQdnUYGFrPQD3nO40G10hQBG9hYnegzckLxwm3c9pnBooSLfJCK
6wp67bMAvkrrJdy4IZfHAQSjqGlG6I5y3z8nFLymfS0vMqDgUirxpKymQdfE7Q3OY1dzetbp0GP2
alvbBN3VAvZyIm0FTfvWhORX0stR5Z3rQ9j5i1JOl+f2La/wclQPtycYJpccyfP6lSQI5h8Y8UsY
QPK6HHiKYfPA9gChsWfdOvyHPdzeKTYlRuTjMnRQ6PVFW+xEZugRpFUh4oBZfT7YinDNGmEr3XgI
k1P3Tx1fksOKnDCYePT4NXhg7xvZH+r6XtSGoIg+L0FSLaOYMqDNE1Bpvu4V5Clgbgr47CR0+nsM
zXt/gP1cPlCYCyj5dB/XCDYq+g5fFPRylQnbPCbBlSPohfT4EOcrFdJzn9cHJsX3MO7j76Q4aUfn
TBAeyZ8oAorYtfGK7LzX+IPM1E3HXq/VKDUtbjBjaMY/Fw3ksutpjVSIIzOZz75S6Ujc0qaAouDB
SbN9vj7nMoXj9Ybt2Rv+J0mfbq+jcVwOfbVzXAtVrlKHax7T0VxEFm3wk+E5FQUba/cHWMmdBU8D
3ljAOgM/hN8tZo4snPPSBmITe9/roNNrwKOUp7cDLuVB+tZskPqZ+FKm/hjl9XcXtEh6lFU1tvDi
2CXP8Y3dO6HysBGsFClBD9EzH9qQjeYmXRxSVkrEqHKj5gvocH0w6zMZ9hjgh21ikObS/j24pXYU
uXaPkMK38bcVLff/lUCU6bGgeBk72kgKgttZZbmTodGSH4r5VATnYPn3kE+H5iiLBvTPTf5Te3Pf
sYdOVjXZ8AysdGqXYQIVkmMUCwHnsxHDqxvosiZ+LqHMxkUmp/NykfLMPnlhYctI5HrW5Pq+bauo
DFZXJ+IOjBZbl++2Wu4baoUVE6C0C4LlcFtsKJvunbpDDR3yuaSr88QpzWOJWy5sOG10UyLaYvYS
TW137IlYo9StWnwDKvhJu+Cl+hvy4RRNxwLUTizp58I1H+KDYh554eoblG4duzqtggE5zXI+EYco
wG+bUklJ3WduVO/7sdgzk1UyaAI1Is2F+vSdC1DjnDRjjnXeTLKVm3aE4guoTOdMMzX9/xLszyvy
G4HoL9b1aighYEfvdsglahzY/bDMjYdUQF1J9U8wnjV5qmP+dBmy8gXXLeV6pbBLACBwpL5ptAt6
aTFZ+G2SJ+VVQ7djcplfSuaHD9S3givsy3EqFaUMNwXQOihl1DETYS/xI+3GBtYjw8Rl887huPS1
mBeM74t86Q6D6BzsqGbRqWlfh+OIMy/4LbKqvmWnXnoSsbXnLR21gGJa3yDSZsR7htwWblIMzDOH
MGkfiqVaz44KZSJPjZ0GW+1CfaK+jui4jvoebfOMSDU18JHdZGzPoUqldayA5iFTRw1+cxQEZuD5
JgmdWh1KQslwROCXXx7OlJ7Txgv1/UfU91M/eaTgMAJ1v0t2UAAap6oYHaY2s0ajw5JL4+Kl/onS
/J1B/A4Aq0rCvq/jpvwQZAgwKaDpNujW7zB+53sDvrI450w1ublv3i09RxJdX7Bk5Tb7vjW9GjG3
XJ+5ChtQjpgSJ2k79ElgryX8jRIGwfVfVijLtzusmiF13bfjPpUaSFyFaYu+5DnH9QLjfWq5M1/8
C4l14KJ2GFvsekZLzu3kCi1SuFPyUDnexIJjU38AoF5SwTsB5fy/xhJlbMdVVAO7hbpKJIRN63iu
pLyvSGqZQGrDyicjRTKyUhnOSi9ZvTy+7No6ekI4/ckPAD3nmpIOGHI2IXcbZZ/07Fuy/N+q9pil
CeRIqpK8Wm25QfISjtxC1KPooA7tVpLnS0c2QWX20ItCyhFP+G/tyqqtUPJxMuuUYRbw5SDTuyQ6
ND0eTOOs12nlkbjlmvujrafr9bjsoU1QC3SyBOeDNVxiKjFJHzDuBcpITHhxYg0roH6IIZmQlyOe
TiNNSWw8iJNmEz5BV1BmlQpWalBDxW4Hu180YIwQ9VXT+Sq98hhJQM7rpzhTF9vOpX3zBn5O71cj
3i/Pp+sOB4WkM5fW+8F/479sXgoP0gnffvU10kkT7scjr7EgflhWT9t7RT4FvA8MhoNR2u0YPRzj
MDm86/UF3eZ0gwDSPDjoiD5qCpzZEr0Hw4uxPdx0zeidxNKf2SnRHv+xQ7fz1uBkvpKbzISzbplX
CI7o00rSjDKM6gw5Mvk9uzxWwTk5+gGl7yAuzhVMFj/4DMwXWCTyzdYsnVQdYZRgj/NRQXTh1LVY
r0gElhiYWyB2o31/cWTfB3j3oWnCvy9GkKjA/LenUJo3vljN0Y/Eb32CvJ2aGQmR2OlipkNO1M34
LnV6VFuoxYY8ORuVLQP5ffLTyrznwqknSHFxRS+IYCPNOiaEzneFCUj691XyzwhLGY4IYR4pkgKx
FijlAiZErY/YQDrz3IBMYIFmLh1yV47GO3NOJvGNhMEvGPB7FulLtzSyaZN6XJmb/0jQgK8HM8L4
ATStPzHHwpkVUDm/Wl+FCwMo+lQU3OyVgt6F3RCGZWrPvNDfYxjj/lApi3LBlbZwUbdBKUePItMb
D+6u0tRaVlR5ZeIjlDoVYf2r5NOyr18omHzeRZ9R8XevvXZtGy4vAgAG6fCXAWheTs1W5hTPD8Yr
UQrrHQgxrmckFqv/y4gcQsR5TUX5+rVDml0uwpJZLj+bwPmx4RpvtLFL2fYHpLFfZ6WwCxUWyXwq
osR7YyNfs+LrvPXWamYQ1s8rHLm1tOWp43NmJV3udnfKgwVS0TKiz6CaA3O8TiY7BCcvmz1EU+jz
wMxEgdG/l4t1lM5cT2QBoSrpxj4AxSkNpagWOUHA8lBliysDygoj6R2rPw2M3VSw3CwqCJdH3vK9
E9uof/fm9KVBxrzmM7g90ubQ0vQEJeVREqQub5HI4xtTtqV/3kdZmtNLdsntdmHmHhGgTAeY/ImI
xYy7opAi3l8QJkg1jA80FROgPsad/gGKJBVvAnC3hyubqjXBFrBpweKh+IFQRHac9g6F2W4FPUxR
mfkq2EYsV/Ku022w5eIkpaKUs3nWaYfgnYT5VIDm0KoweG7iUy+Mdacopr2hSbGOu0A6dOHpgQXe
NBYlG+FfSicPW7eWmJRAdZR1TFKp0U2qvc64PR5T7pDvt0DXRljr4DPqCW0OWTtGOoA2gdkggwcD
voerymGEZFi/0VaEnu6fOO6yP2XgH8Q3nzBTzpT/mGO6h6/a2HSxcT5iKMIQlp8dFM9a+Jg9eAhV
hWc2raahpgGCw+mQzAo4Q1P70Vo4pSHWqTUXZ2R8AHZmTFaKKN/RUmYQAOkUJ89Y/4oNsEsRWW3+
lsDsFSdMPou64wDZKfPlThRo0o2hZPpOi8zwr5cChck9lxFx5T2F+13FTmhmq2yZHzBUXT4yxYGz
E3iUErVlcYe9Hv/baxb8fqbvtS6n6LIqdjjbhCqanfoZBRrneZWmS7GlsrMhMnbC4wZC6JdXu8xl
J7VCtBnTWpt/9Zmucpea5cryn+JIRNWWZsafla9gTmkSr07eVMGvLYXB4AAutN3PG7JUFxgqR8we
3j+spFvh2ZORTNJsH+pjX7arSuGwLJc079BbTte5J9euuMlNOJJz4ridsavIBNadkiMHX0nfK9ab
pNXh6t60Z0uVv+N85hL8OowIgdujLmHYJtcon4iS06XuTh1ABLAX/Q7nB4Opbl7r2J3AMe53Dbx4
bwaVJCaY5BY/1F6F6Ajn+FOnVz1o4Ui40uH5L5YPQ2O2Toa3sXqrlwsSb0h2CqXlKjUpg/r5ZHQ/
IVeYEMXqwN+AT9H9cMpOnadw0KWyQYNKjcVs+lZunu5ddNeklotb1qRY+ulpiQHIsqSQC8c6t+5f
9Xfj1q5kirze1EOwUPg1VkXeNGkjJ4lZHzMFtrX8coBGnGqXgx9CU3kizAbXI12wo8/1DELx13W2
Ul1ZPWqpAJ+ybAqksbk/M+HuC1vd6uFrx6HhwFNe1rDEIfaEDHbXHN16RwcwMBWf8ot7SWdoIPy6
ZxTSLk0v5C9QVzs12DYURUQNRNJrcGw1qI5S6s2r97yaYBDgF3V41KT3+Qgx3W+JWSGiGPqz9+Ge
XZQ1zoySQ4yzwXwN30mhpRVuaMXiMwJsUzevjXmBCWdYIK8MKnxpIRnkYFWMuKO72vsRAS/tldtu
J294eTnGrpUlk7n4C9e1LV42O1Rur9XqvKECiG3+dEkWqBmOf8eXb+rL33qFi3olQc1k+Rs7ijkN
x6OB1bhf5HUbi0n+viEjCRtf6GNUi/673pY+zEUGbiuhwFbe5z8/kApJkmA5Th3+JgyxYSl62sim
wKTuI780VtUhqbdHJFatII+3aanVPNoZXnIs3qy8s2SMxCwfwmmuUHM/4Hh0B1/rKeekawbrFY4f
dS25KQZyTDiqrMxKzCFwDFYqbrmrgC1f1PHOZ8g290l/3UzIYKQfdiyHtuJEHZKa2perzHbAwHr1
Fck7cGSB3XrIu1MwhWZqH/WeB3XWyOpzWVHY+9fKpGQ2C1/qZNI317xLB4RkGupQKBsnNEiB/gmc
6JSZJhDWE3nTNGipxLh+zAr9nEOS+C3p/egKdsG5LKaCDrvkB0NBbczUKtVINNfzLgJPz3epSZx/
XJuzYhWYemYsJd0tm73hsSy4qnZf3DhYXQ6AGGoqLJmEViO6wFiQCD+qOxOLtAmoUjgkKUH417NG
VuhfYaGMlSxoJMpytoSA29oTWI1HuEA60ClLwsxtsY+tXv9Wx2vqY1maxry66vlrDSUF/PZ3oFTS
Ajv+nprzwpmFCaobZT+uP7SyPIyZEhAmhpyGO46F35e0I581rddCXvvUs2rp09hsgsJxMs6iVUYf
eYYza20pVIC6xaLvypXhI2tetSC2sHdEQkLcPDxCnutetiqas/lt2rhUPNuZz3MXsDBarwpWPRG8
AZbUD/CrV39ekfiTsoByskjj1o46uYx9cZYZR6eQvRwd/u3vL1/4u+ftpbD1V0NZIsmd219qwXJp
6i+zT7bYzUCUhO9r5K2BBs/Z4/iUD/gvX0/FD5o3JoPsqJspkT+iRwSQSaouF4V2Vw1ER/Sop8kp
gOM7dMKypNUz4hxBDdrbdL9cnwupsIghZ5nuutsFX/PTEseMEaurLni2R+tsEWjUdBnhM0+zmJu2
iIHQSAvFqdD5nJGCnfXxKZL+ii8SN5GQdZfN7Q1tEH30xzcXb7x4tc8ic73ALAZ8YllJAmKsRpU6
Ku+iz7MTAeLq+k5xDM3pZE49cxNsTWAb/aqLp5Ct03cmWnW/sk7nuRvgagTBs9iX6DEw04BiM6RU
cJJf+yOhXnOVRN4g0U34P8g0aGmXd4P6jhH4W7wyy51jDL/ySQTjQ4N6psI2ZZFw12u4+SPn6Odl
TYRR3UesP0g+qQqUjRX+x8FfKAa08RUznPVHEH5fTPfAI3Rz8w/eJmcqB+fghMK47NPA7b+AiEuH
YKV9K3mJbzp5RpO8oBhxHqTk3CoVsX2JJoH724wqfUN0gnqozow2PLNBdYj5lUXcZY2BppJhupMe
DCeX069YN2YQ4opSOJRQqnf56hm4LXI8N2Fa/QJ6+q0ZPuTP7EJBqUQlfWJKeE6juAbvusMnrSyL
k6VV+EluOdcGKEm4Oo5SXBUE84NqKMg4/6MPFsNcXZdYz/ToJ1wI8EIv32We0pUvVds222tp76qt
NwtYDACj43gAPT9HnH6Z7f8czkjwgBFF+IWtb6jumkQKcbciCRbk3zduzJrbfE5IajoQtwFuGPy4
KsCT6CJnaQG/D+vMuiuXazxh0K6/RBALoDPM8Pv0PezTTADZIfcjBR1UB6SPiQKIJFksBQRgfvrY
5Fch7fMiaqv2pizXzZ9q0aYmoKhTbnuNfHpVzcn1RsOvs/rfC8BPkfdhlXdsZosYggC6yn3S+8sx
fZYgzXjTih9A+Mapi/YH3cXkErp3XZUQdmbb3VEL7MZgpwiBfohhkTCmauh/YeQmLRDPQ9K464cS
NxE+FmoUG4fTFxoU62AxIxkfvlm3ienGxDcahIm08cRC6a4AP9/QsRiNgDtclqiL/0MxE8r3LBhp
z+iYsclPfIwYL3BK45dOYCGjVF5D1paOH+r4JwrxB8CLFxpSSAUdKpcFpjEuAcs+V2Ys6TF4bezN
ZBS9o1gO4G8cu1k2Uqqe3qfc4VOkN7lxCVQ0QtXf1CNkLSar5dRnqUB9P6tOgbIs5GWkfzIlYwYc
o0ht36R7pEToFTxY0aIQCf79GMj60xqYdvac8t0Ha6bbIKFBEd6RIEcjX4kHay9tvmNMWxG9PuFW
HlGh8YokW6AbbbzD13DtT8OMJvBs90XnS7S8QZ7hX5ewQF9L/ivzsKhS0DCA8fkcNLHkKcAqgJPx
CfaxaXMAxDQyDmTilAToUVNuqI1i/Da0vHFwZA2NRFrWaWK+YMgjpyNTfpTgRackwrleoMowa2yb
ZvB3ApQAFG9IdEqhajQqc98VGCULC3G0u8U8S1L2GXYkudlTcxNd/s0GgBIvpH8xhq+7eBY0L89u
EaBo9QEkmZJAJ8n0+bJ64Lcja76h27Hfcq9dtz12CwbBrg+EZHVIp62CsFoHYfPelhB5sQ16y8L+
BJU5t9vy0wCMh5QJamTvyFmbfdX0FsejuMfObFyFxXX9pnpY8KwpkBa+wnemHQ5iejXq7Ys+G1QO
PQJsmIAu9+3sUPoLzQdnY7PtKSGjIcKPfKdxUCamgq1lz3xlxjRy1NSaXtK8wFBy7LMT7WN/RAMq
dDK9xlcZDtUBBfeQlcabhi2igridHRyo41pSClvseeSGr43U8k5vxd84Ot/OSGlVvPIL4dc5rp91
KD8fx0X5jxZ6ZW3O6EW3MxpzU9ONVrCZOhc1e/0iPLwQnwO161LXBpsEmuCaw8tfHJ/sW+llBIo1
2I7KiIpPalvU+c6+uDdoFMDBeE3rfrKhxJaQPLFIOfTj0lCstactPL8gHEMtOtaSW/eI26xJa0e9
dU/PlxGDjBu/XRFKXx4Qg7MiLshit2vTahwdSq5MM7DkCrAYtqbQ2IWqkKEsaeXdOPpYQC0caMZf
XTtYcWL6PFr0gXburZTYT7ZomIDS34ogvzIWt5F7hM1H0SRAik4tUXxe546G3AU3gy4cN33MlTP6
NS9d1uaYSPmlhi8NFTbvtPBABZlLbgk6WWlaH4fSQAf7f0gCTceYyfHI38lJjhJZXwXCLeTnyQG+
T7vp8BRXAPiN3QN/OiwEfQ3+MW4pZX0s2Zw8qJRPOFaPh1E1AgrzX8+ZM7ooyLDUpvNPIuMvokSg
iMpG6CsfrnfKFesaKAE0Clj6mIxkbamtQfKB3IBaoR/y4cuDjrK60ftmw5IGmknFEPrPESQKbE02
ZBaG5XTtGTLn8M/Eo/WBG190DzH1qSABskr6MZr2TRmT9gERfFxLGs/ncEpZu+9EYlo6W2VP/gSk
rM6rFQWEIXoKpDl7gmuX1KOA7hklRxx4+UOJ7RDUwlc7pNmMi1xbu+Ls7rtSnFYtTh2ax1EZCW56
fiiER/Dn85V3eWWxydAwlYlD89fiGKHyh9p9vFBlORZxYo1BwkO7llfQv1E/NdS9nj8/3rQpn3NV
vIHAC5GO6XrbYJgBB567qgYgKsYLlH3iQgCVJA50KZcZKioJKiX5qMqeMpquijvkkGqQl6Sx0YmP
mc29ZX8Utws9wmJSzqRu9vck02iSatFAU8sjg+8ZgPA1+JUx+K7uC2ediGyM+mo1hxgYFiXElDL+
qqAqRITL/2ZphycbM9/U/m8ZEXIdK8kfg3/zWaJOdv4cGTyNpea00AYsvu0y9IdpOik+wwCg9XEC
2gr9ro6rDE/hDPQ4VE3wyi5NOYnibVjkOwBkL5tFnVOiRb8s5flmzITelvzXt8aYigDbVRZ/mJI1
N5gjxj3gF9ld7F2SnqHSDhYlLHB+dOzddIKeeAF1yj95i5jU/ZMqY6EwWdVYF4fhADpjIzHS/p/D
lP9V2yU1mvMAM3SdWFjS+/vNaaWcyNw/M+Zmnaj55RleaihRw3qvfp3jN8FHi7V4762MchqZ3tLY
m+UUfEp9vFgT+cy9FBIblgo4MsU/EL5IEFuyc7xP0ilBrSm10QgVee3QcWCidVmHX/nZWyPm17u1
lzlqTzDkEeQMUhgCl2EF5qhweX+eKUA23R4bjuP3Z1ubSClGcqxGMVFEcQl59a1sJqXPRulVFwEU
tW0+G52UJsmx7zy78aABRXazf7lt5eFx4bbR8j0fL990pW2fCQNu7Xpimj/wKdJmGohIW4MgO63U
1bFor3bw7TnH/nGMi08FldszG2vLGbN1ZlsmAbrYjmadoVyA3C0lrFsk8RIlnjkmjx3BzLsvGo+B
MI6fkylsVkAIkinxe6Ek9rOtTRe9W5NwiJK2dJeb7FcegOKWRFbbQLzkL20ypSA0ztiNJC0qDPNJ
86HNwO0voCjD2fQN4+Q0fksbHrWa7lMAjxf3mz45pBku7aiYSoW+mZlXwoh/WqKNwEwf1udyipSJ
ihKsi81hNIUNyBH4bpHxQVT9d4ik8kGz8e8S8oqQQ5wT0OwCY6uFPiLryf4J9jxRxR4SErV569zj
3ADsI67W7yjyDqzMwEfJGVlufHyqawqHMX9mGVTQFLVrtAaQCj/kpe4NAQo0/Is8GSdoo2ltWOl7
r8B6/Ffmrh76UlfEr7QXyTOt6NSSA3OJ+1OZp08h77UrRIJaCnuSOeBbM/9fE3amCvzJHBJbqJzh
tdnx53iaUNlfUFILLJiXwaeNdwdeQwQdKyIXhtGZr5/Q40EOkax8HbCoS8f11rif4ADeb0AODVrW
r/hXrn4zidEEoCoVOMnaZr7rHRiDIktkWjvslvT583PMnSNPWtXvfC28K886IVzlQ0OJBhe10dIt
PvhnL6bRwmnaOKGfToqk240UgrqW7IfTisO9dqEUMO01uPpK8X4TzaL7vjV/DfCUepvAVpeAyXth
nAvpU+g+NyEGAupwRRj3tcZf32zo6v9jubyLGIPgtZTM3lT7AMlPOacrwmn6NMZcPT5bZMsCPEzU
UGaAqw1A/iUlcpTHG6tmstVTlv9aDEqtyKXAhdn7jgKzjwabZz/WESLLiQvqqam/Bp1zPoe4+Sy7
8ErTSL/5g5cp4qVXq6rRzc18DMcUV+aoCIecTq47bj1H2IiINoecLAh6D/kTPntUfeSN9Wjqj11x
wFG4nn9MwdkuoMRbNaP+cqWtF4qbHdU6XTQSw4/dm/FfPKA2+IGLU5SSCbHMqF9PC7G0w2DSyWNT
k+wMW96kKPDNuXjGZQjePJ6uF5OVV/H/nqh/M+orWDPEwBlroYEVjF43pDDjRhMEfIgjcHSJ0g/O
OwjP3SvH6VfC21IGD85zucG32+ye+zcrYSacLhSGPvRBuMRsVWRq/kvNTDEOEOGclg7p6k5InQd9
at/RGznybEqymmimfrR/kt6/EYLpzRoHoOqNSQoRVGPV3WVyeKsmCKdSLoGvSgHA3dVCk2ViVs3r
SXQg1O/HkmWYByFjLOVTIpmjiDut8EyUHBNpMT4L2jh2qFf/U9+jUM8+3iO1Rfza5eumWNjcenGc
7KnjP3igFtttCXPIpHxQpNPpxMlyLm9/00ACsALh3BnYLr5/MGFYwvuxoc+/WA7snoQqBb+j6iWT
7WsYvvdO3C1If7rDpNnh+D88eqWASSyRvVn/cKpBhrwjeKqFe4k4omr6RK2cg6yWuFFAi6pH7FAF
AWmLrOYXRxUwCtEccbN7BLznIowx6ggvoreBRxpKdDgsK7TLjKUYVUloA0nUwb6jR/HaV1PQG/ux
UugS2TDq1DaybsWdNO/96nTMTarHtnIAzGwqZpdAuf1347bsrvhWmXkidwbvUDpgKCwqjIndNHgF
Q5lyaARxPn0joAbt3aa1aqElyBDs+SfnR0QGEgFqzEsx/z3bd+XhXufFooKLmNfKuohL487FcwgO
6Yg78rE1YeW5NvymcxaddODztSM62VCT72zV+ebl3zO6gzynAd+W1yrXjfyFWufJPWmvqvZMwmY+
4QnP0cHXP7MukkR5rSaWi3PRhByElMtiwgqaZbCqQaqP1aKTxhPiu13bQHRmDmrCnzYyMFFnxn8P
KuquG5ifo3AZwRzSXvtPr+7GM1lFiHJKBpT6ADloezmy/+oWZhxIJN10FYg1oZe695RoVv1K7U7j
x/RcymRXG+WIMTb93ECE1uel+DxF40wV2D5cgVdNrflXdgIUwivaeh1fk3rN/8jWo865W0NgXRUU
XLe2dcqI6B2MIgonG206bnHk3/HWOU2bZ8iIGGMUvEQy7djS7RvTDXoIdy8lc8sN9r7bib0tuEU1
rgaRwB2kzy+0d13sahOE/Tr7zSxcQbaeJRwCYSVx3sADRlUqdEZMecYYIY7nIMFyY0YJQizjdXht
T/1J0TxDxoYOZ/8rebDEOFPj4OYESh67/DOpwV064xJ7uR7bOx+Wo9wv8q0rJTrCuG6be6zRN9fh
t3afv5AMeRgUb9pyOH6SsKXLkaEbABLbstWP6m+12BojelozB9V1dx6+LmtA8F259Jw5gCvTmzt3
Y45pqxxkB5ZzXgMNt0/LPAM5MkabaVZTDOtyWScJa884+0zkt9BCie/RP7w/T0xVFRe8LEt8e8tx
um1+swWcx9SSdXjnnr7cEUkl6aolLyQVzZLRqmYmTKFj1UE7yNr446+icFjfGG1pV6bm7FOx/9lG
myl+6BCJae8jgSCEvve6q6mXZBb+PG7Rk5BrE0SMgvKjE+MjxQbwyAEAMfkaa7EvyY0IGylwVUn4
hauf5p0OPHIXR5MKRafrr+t41/NQlB6ayvkbVxj8Cdkbm+GsBDr2icw7fCbeSv4f+mIhEeGOfQBn
nZH08wDk5wpqh3oUOXr2Aa660UtytM8izhDEfrNIhwUL4aWdvB8BSRgtl8pKvzcS8hYXQS0itp+8
MVLlGPIvbo/ugBW4YGgxQWCMZ6RQUvAP90a2Uk27KUaNpIj4iuvWa64WYqeTlUHDQB1M3j5E+ZJ2
CysZbIgsejupvobtbGYfvxa5f4JASLOaAZ5JoWgU5x5RtRQ/xKDiVgUMVT79lRyL5qlskyHeR/iW
WBM10zx9RYjCtb/LdZ6sDJptzHdyX+c0+Ho0tp9/MLaul90yz1F+MZkntm+k5LYuyw/Et2SX8uCH
PezAgDuVL97WTO9BlcORUOEEv5UlyAQACq/VeuSkvB+wMbBZzHhx3tHKTzyu4p6S2BnwlWLHw/Ff
tLTtNFYSr35KQJC33UhLxRaadNePdNIlKB2YK2n8KjLqotNgn0zMpuFoTiBbXDpX5zpBONRf4ACI
JxKzo1AbhwVhiknJcoebBLCJy/G8E0vxIwjbgzCD+fAjqiYFkW1qa52GC8dcfnmbimrppKwvj/Ce
HLnoYL/JQeIsMOki3CyXo3fqLzxTxGytxDkxPKgZrnQ6T/WdTLmjuvAP64Yqyu5CwvYyAPYvBvAY
SE5qJLD6QmqdWFrs4tGAZBWkSFk+/uesQMXL/tuesEpItjYkOm3/Ub3S4g5npNwWuMhuKg2n4uEg
6KtWtiem4MsApPxUMtJiySVS5Mgs3FDJGBxVZz/zECZQJxTDAdjPv1X0kTe7mRWR25ecZQhOH18t
04wEWyLCJjkfX7O/YRi7HmvHQZBux9Ubqib1rGOEV7JRe5rjTi3Ge1VAofLKPTKjHbragHITqDYB
lBoL6plFUYoaYlpg2B0aQtR5KUgz7CYplgsioCVG/yorApbKBVac5/ZZ0FH8/qljbpPN5iTGzYG4
AkHCv3qkEDtwE44BPWuiVtmTKkfZq5uBDKrZN5TNt7TSOw/zZ77WPYPPB3l8zDyrV++rkOBbRrWM
zoTD0tUrYf5ygSF90Yv8Wfim5ZkGcPS05+skcDvU2EjjjjT5bRhA12YyHJ6olbMPBmmdm8sqGmtT
zcwFE+ig8lxUFeXjf6DdCXvqdv4v7k4gLWYZDE/EkWTDYgKakXgm3x5Objw4OZcvrOTV7y3tFSMk
1yE30D58uhGhZduh0Heiye/rDAr6e9qpo9S6gCxNqq3UKRRBeVogT2zll4ydezzh4I6V+IuUqgAM
d07eiDXS+HI9qxa/eDbwDLiI3PbkcR1WzuLFPkZ2E6cbbsmEy3lCqgntPf2KTGW5wYLCG0/HgbbD
Iq/RQ7Il9IIBhGJC2EHzTc3GiGCdMyJZngOyDBNCRjM3/I+dqeLehw/+sSfW5tk6b1tY0WPUKAAi
mAtjrMEpBkRYVOuc1AQ1El2Er5miNNSq0aSZFN4ChZWKA+HX4eRycCUfBFe7Map3jJO/FVlVhLJi
Y7HK0sWWGuE1OqtszAjgjitQNAHnRQnxTQDOur90AWISUI5ED4v6R9miQPIniteGKmJkWTideNvR
T/2y3E2LUc6RzYgdwDb0c12xsd/fB6bYs0BTRdNw1EGJq6zr+soaJMtwpIGSNswTI23QZ+ONlBKH
qnFWWegIZo2elV+M11EI5hDhKaP2/NsaHDLaua3vysjvrNZLkms90nXDJ2EyMKfmi+cY3HMoZEGt
ElO4HHPE+44xpy+jstWo97TU6xzrMVMUKmhR1FFZP6GL4RH7oGnsPb+mVhwdvIQIf0+GwKlLnPv+
csqof4rzLXSnWvUmlc+XZAv29ABzm3Xni/32PmIQx+J8SPbliFQbvVEi2qrIGSxlC3wk+7m43QTx
HEtyJ6w++nqqIl6yaFl5ExSooJsJuPK4hf3O/JtmV3mSHKVYK7FbTJxcdVocwj1qxi3ttV3f9j15
CkmJazTi13kByxPw/CUxHltmDYPbgH+UJyjGbpVxREi2xcja1E63CgIV1xieMCCkwQEoJ3uZY9RD
V06C4hU9sNZP+Cpyrag5l8ZAoV5i2A8+sqDBeZ1/7oiCeu9XMM/Z/LsFLPqJ0U1+YZZpVlMhq7nL
Uthqr9rX7hdwbA5ZzPvF2ze5ENAnpwnmNaoVAcPzy92VXiGbeCyE4dDyyJWEIOob6VeyLMaTWAzi
eLfNUJysnWeT4KoBBKOB39V9QzV66nktGkLB64hxB9q4F/M0xMM6X2pDP01WIvR+FFIUYWTIlRYu
5abq0BHZ/KRVpRxHX2HGmD8XsbQSC6dGWVIYDPfzLff/wDmXJ0GLI4g7HDoGkAxT7ineSCXLpcwd
W5dWuvzGVfl3gN8oqfCAmfQAcEH0pfMobzpBobnB91AiWKpPkLDXp4o3TcGZGvmHEsMktTi3MOGe
pgAus090zJssazFRyOdrCXRWNbHyoXXUEz5P6DHO0nOa5jAd2TGuAlyboAHFwYHsK50zxtqeuuCf
nw3HpB953x2mH/EhpKFiKqb4RTyOgztEKWd3RUEByeik0NImwxMXlClz+NlTIRxFWXeFWAIxmMMo
OePJMWWXWwomxssfq7nr777YnxH/aEnQgi4mcD/7ejCMK70+JycpNeYZEaEh9VPvzmqkigJi+Rlh
rS5enCx7Gbu+VcFCuPz/Okp4vXZ17as8LUFQ/AHzDWoZwsISXEYi3BEA+9h3SflOzD86b2Q8Cjmd
aX+ABKG8n4hNK04UGezNvc9dnQwIDY1k5LGfSrIycx7FYFPMWt3IE8Sk9J/kG5uGBwWKzxB0gj8e
MXDY/g8cElhWpOIiZRwpOJohytcauCcgGXaZwD8LUrBdcwQbd1jWtcQlxeE63tbSUf78OHXq9Chj
vuCTh+u7V6oZlH1tZLu4uRM3Zty9vLgXJeGHgkLDG/w1vlrts2mcgePv+6SDylzRiqBQtWd/3WqG
QhCg2lQYZXEEJZB/+XrRrZfGAKCasNIcxJMPHY2v8y2/DgNO7tIZbdP4MGRFBGU5WhMLkDXKBkKZ
4TxMJKa6Rmj2ED65YJdefSqYCI7CAuKJv6BEprYiSYsY9vgcXLNnT/SwIOeLVywv+dtf+mF9QOLj
lm7wrlf98cF4n//VIkrakyqWG/lqM/UgT/i5S5JmdFNb8WN5pFRygpsuJCsblYp3IxW3ll/jNe6Y
2TKXhhD2D/0sLiJQx8E8S0fzZaxIxrN8AqTH/0z60iJq4zZBRHt3Zm5SYUu0m0ruvQoDe5W7IDU3
nkc6ruSqPyLMCXkpgYWrmap90cei2Cx6QjPF329FEkHUe8AzA1Oct6jbFC9o7kwMidPGjCqiFUN1
fFS4ngwFObep0H5E4Sthsb91bK03kxDQ56OzYY3XamAudzIYQg9YFHjONOI3Qu/J7IXhtL7M5TM+
VAnx1r1s76ctn00Xl755JBceXzk5RCCFhKY05BEpqDOjEt5UvDzv59aLt3dkqzQ3yO/5OwhOb1Zu
tOtqNM0kj0DZEBEWuOmrhvIwhqY8OGxqeBcCUcClS3N7zc1gsLYZhQGgLqCCbQq8rxoZH7ikCWs3
EPkvyzRZqB9dk958Qg6AYkESsMzKqYgto4fPkEfDlUYWJ0o3Onbs40p6d8dQkn/n1gJmkgxFDIFD
itZhS9CwMp1xG5t4LQhqwp5tCZbnhUXHpNamHWoGIaOG8oxxK3EAJuLbM+TLP86wpKaFTF1Sv6XI
t7DZVgBWP2mvJ4je3Wr76yZgpu4Gsmkkpk2TVnU6hqkFXeXTBdi/qyBGLAJfwTyXMVHSaWICLhEC
LEGU7SLAS6lget21TZ7Inm5OgLN8HxrrKpHMapHlefvAFprZva95+1BhAUaK26ye2TSCCB+0DGXY
aVnaaYsa797xXj5DqYzmzDALQvJ5rDCuvuJKmxdScDC5Dl/gBRxkg9D6/wJ/s4y66FpYfdnp/n/T
KSmezcFiEXbMBRlZ/h9x7+mU3A1TZJMfM9nRCwbnlSuHHiC/conYiRoqJGRf4gzeyMQk9Qs1wxBd
PxtwhsFn5i53L1I8R9m/rqQ8/BErMzJuMdgOubOdwio7VJFNUYT6rJ7j9HONQtBjvstnhmF85f3b
+wXl8oOpI/G3zSEj26qPl9NtNFxlLo8eSM9OqpeSjnNTv1wrqeXap87AklReucttF4RKsbkY6bUM
F6IU2GfGvPw8U7QP2axr2EK2BLxL2tvHcp83CR1XwmM3s88Uqob1jeLajBEa72IsmyQJkhqF+1ph
f/kHgAa/YXE47R3mOmcOcK2JPV/23iAnG2CetM2NFSeSnTnVOXRi4/4sOWh2ujshhoGBcoNEn0NI
QlidFzfBEsIvfPgY1YHn66V2OiG20wRpTiaOpQQ94BJq13w3gpSDa+GBSPAYFe+zCxls25BuL6Gf
NDF8+GEfFGuj9DmsCpb/zHVSAHLb0nAvp3T2HA4Ug+wCVRGVKi8BG3HjCSwhLWCRq5tUumG2QGKe
FxKMyyMAAj45GRVXvVgjZyPfV5Ta/DVKVVC1UpxTUuqO2lM5k9bdPvDW3iQ1TnnFsQZL32JXKeVJ
rPnheJ9A3Ysb6sLynnBTfykXbQpg5OtwB3szoDxrw6VxL4iNl1fM/a+qo7e0Z0lVDbvrpe8HC0gQ
M8u4QBXHu74t6TW3sNiM4g4JBYR70ApxHOuXoEpUHl57YO14GCi9rYKRDrWeIUpyMBFhnGwaMVsE
DZ4QAtWZFlWb0oWwCIQ+VAwNnXHIZIg2FUS6KQP7bNopdHSeRrreUrWru7u6nIG5NklZx/i7yqxl
v2UX2h2z6Z/+nzPCYVRr6NggCuz/CQ+vatWgjelUdlLBEoXV3bLbQfdy76+RPf13HwUgAFvzGxGy
4kr712UnEGEUVAdhUvL9+GrHxCt2DitFQvmcUxwlQEBP3YqSeQFHZjByWVIvL/BBztjtC3I7avag
zMqxGJl+LkqZWO4Do9Y+BxPqrqSwzeMmgImzdyXvCRzdCRb0R96noe0brqHA2v8vzc8jt21CALdf
lt7NlP/l2y8PiCshRrGaQEItgn/0inN0K2XuHS+o3yW1MEOm5OQq/ailoSqLeH8/YQvAqKqt3Idj
y1yjHq6DivRDQ5lUkv/9EwajDlAxleU9UETtmDIjM0NYwfwNqmzXWli4J/GTZLKo/YJnxJTCClZz
JAL+EL4Cqz1cI3ojf/QFhDN+jBCGUmYe/YAo72hhXyhv/A+rXokIYcMpmf8s0aTKtclfdjTNMq6L
PixS+9fycjfkZ9TE6wrBgI8c7xb9qmkjnf2JU6ha9o7Bdt3JfDzlE8uBbEWqEMJjuPbqltvpMRAA
co90ibmcIuCiRxDXBCfjBZiogPiZxE6ShSy/4M6bcze7dLdQK4fPTHY/Pfn+9J5lqp+dOB2DkRBL
rlEtNq/GPdgBMgISIW2QxvgxNfbujRGYOfHX6CqQ5ynTNEC1t2U/H06jL0WWp37YcclsRhRIXEM1
cS3pHs8Qxbeu0E0nGA8VNv/8G6EsyP1RMi++1GmECTXGIDqTVtyvxQ49wZNH6l9QpXnis7deobFH
yC9o0J1PEhw353UHlbZCWGnXpj7yJi1zJigi4djML2tVD8aj9OowKH+E5trZfmDcQfARtOqtqAXv
g5n6w2L22MSTfEtS1GLFNpHa+8rRVwSNCpOOYFqR+ad9Yqr6faiJZp2vc1Hf9IHJp5+G2j//Nz3i
Pf9yeEAQ0anwjBnX6WSt+O9ZL3K+NwEtigRIW7J93lSUN11OsNIwf2inSmPwTuYxoJ3wL3Xc8tmc
PqaVzBn5vrW0eW/CWvKT2aYJli88aBxh0nngClLROpz6Xyj1sW7Ftz/xzAkQ9Jb9KSVkugcoLswg
APip6kJAYodsN5OcVmxtl0cx50WKnyglnbJrEPHOWiubQhseVDqlcb81/Pimxce4zrNDu7g1nzcS
HGbZiutvK4akTYLBJEQxJIBlKS5yHrd0Dkvyqduw/zv7bpmtX8P23Hz5IB5Q9R5pSsPnHDjNimns
ww6bWkRHIXq+TrC61htrHhwNGTLdPQchrDLNistp6fGEXx8bmJxlIF9gC+eN4oYvykJns808JX/z
ENkbCQNGK/jb1M+wYyKop7ZxBD1UUkslKNZicJCX483YPBuSu3tc2zKKjYOuIk1gLAtU+9WfAo6r
oUepzOZLquvMq4bmZ7637ySpM607DyFX5LdJ3w/WzcWalLQxGoiUVefmbmDbUu6TQmxhxqocNTN2
TxikXGldw9K2WwvJ2bgwf5bSfGcyFscfszFt7LuK4DL979nRAFh4FTSyqPc6RGTTznB551CsXGZK
5swOXrSg3ougfHwPw7Z/bGkdKqAasf1fmnbkveEgPmEPoHOcA+Xt7e4lJjFz1kYNtkUbBFF6gtX7
CU0G/JfO3kdpfdsFTyRH7FcCXCVQz2PGdAyTCfl7BsBvor3CgKQ83cRkCh9RvNidtFN/RqPa50Lv
4yH0vI/QWX7PlnQzMr56qGRpE1apKgh0ZZ37/2MsukHFjR0kLkP2+ZpEoiNC4Qfv6BXKggyUQH+S
LiazQKcEpXz9EeNlAN9PdwhT11jF+T4H0KTrx71lT/zvvWCOed1AhG+YWMOH1KoikmeNd0Y95iSF
KiYaBtI4HXiOYNYMyaCLv1d2xOaVHFYFJN/AEP5BTPHiAL8GJBmy2uY1SWJIGJmgFI9XuqMhvWeG
0obKKjaEi8vM3sDUJ1ZqYlN+KenxPYJNfRZ39S/kKSMEJnuWBvQPUDUeAg0YNty2atjuLaG9p1E+
IgF0tk8MLos+/Cd84oMF0Bd2lkrDMMfIEPWJiALzzYTMv/mYMuIeWWhiIpejkbiYHc/6f/FgKede
Uzpdxk25QKV9jcNCv8RKRQx/GOoV9oGOnMyWnNd8VyEnMr/EdF80N+GXsQcSNGUn6HFc56Ow3dG+
0efv/GgsuE+5Z+B0or9UGF10MyNgcfTMrZchDwy1YxN3UWIZYi1rM/nTqkmqVz4zj1+oTC19zLe/
oiBERBPRb91ELSQBBFPK/9SJ/ZMeZ6+gTNhdZhIw/no+/QtlK8n1Aed1bsTiYBJt+12oxTMew0eg
Ol8xzPLXHEI09bV7N161eFrw8q2SY1tYukSn2dJJBKqHf3tSjSdOjFBMMRppGOXmPgUlnWV+USVP
U/zIbyTwG57mat7jmHsqLNMtr2naz/qZA3sUTDC/pOTFQJNhGE1j4jAFxEjPl2YivvyaGl1N43YM
hEq6POtOlBqm+z/PLUGvWFOfkq1RWkcsG88YUKNj12MnQGCogogKCMleJHPF7/hKI/UgD02NCCv5
LPBRRGNerGS90EL+3vvpLak2acxJzDnx4fTJuQEy2+st0Vq3W+ZuUYixN6TI3aroKzWNZ0DZC6+v
fK0vlCI3AAud2zo7qJvtmKxKhP7EHIKdsSwttYXioBz/WnWq5ZWReQyhD4MZPod3Nn9p1gqGT3Iv
7Y5JQA+t6HkNU/5Gh8fwK4UhTlXjkvSkQKeAHEVHFQoN7j3Z+gc7ib5WlO44sU+9nCdUcS6mN7la
ADBY3qxXKveuneJemNiSdJa14dk2Kr85WKLyO7Y7VZc+ZBgY/DXQysSuBQ+mRtAjRQaP61FtFtU3
rkvAi4cWz9vsov2gSLvt74YYglUVUTU0pv1xTNfrdL1Ua5LcquuiDyFxOwYWFE79WVe8EeHovaKu
HfMxZoUdILseRsvzNJ34LXZ7/j7l7C8Mw269n9rz/4Ck8jSnXUs5P1IVrM9PIuWdG0cBvC/Pbtk7
JWWcyYlsuwjFiVbJ9WAXa0abCyCnmzY93PzK8PBD5j928HRuCTPctSf8WAzV1XZuVDk4ZOIe2YzG
UfO9qWZ2Lb5kRF5JM+1HNXMusBAz5fPusZl2ekX1OJHlHO0BsYXLNcrTuyna5tSuC7zfqpsUgxBk
2wgavwKrSyANTY5Cc7RK+vwr8n91P5JZkiTBbpSQdb76UnEqBdiNGPD1WSGYxJ8XMnPBVBQsH3gP
wlGAx8eFZ11wqWi7B9DgRmuRUhZmO8h2NsBcXk9UNprfnBemIWqD9tSbmKXmXOB1Py0Go7pwf9bM
+t9KnC1M9yzXvMwix+QA4aTssKCnKUf0GVJC1CYW/qreh3OOYjzUSpGaW4ObyREpQBHGiegezQNl
5wbDWAqMEtZXWpkwrMYZeR5BRGyJHMuOUtlrtMTdNn2Ln7a195cen0xp3HCzj40C6WjR7gK5Hhll
4F6oQRcLdO3DOB7lQ7eYNQ2jF108YvNhDxAxhJfVLjh8snldzPFqlX16M/s6S/xx9Kg4lGKJb1QR
2ojS9uOa0YbY0q7aIkMkBwckjDC0MBwfwQci1qRwVx6yI0HE31iA46tx1rolV1coRkiqK++JlV+r
YsXCy5twg0HRDoRx9W7F7j/D5l6dNNR099c+sQp7GJp3npi8k0meLEgZO2E3AXpZXNlC3NttAO2V
qqG91hMiEnRAv6Pl2KnoirrkJzQhbLa7XfMbeFDOg9dKgqdN/M1qvKd8LlgtE3IArIG5OSIQydLN
7FmQCFYCcYl1nmhP3PUbeO1wPOBBl0lZuJ9/nUyLHPVIoNY0R0PK4AJPzPrr4otQv46XCgqvImil
D9KhBmjnDqXiDfLeNp+E0EWvv8y+GDdtLIcXpBRGrVKd5aq2/6E5H7pbrvZZmctA10JGwhMIQVlP
ICQkLpu7L3GhyfxnAt9k0LhIQPv2kA1Bu9LPBLUJIk1dCbv4ZhrEI52l7ucaY2VkpukKzk8efrAV
q6jbH5+T+wVd3R6QGMjSWL6hiGD/d5ntLlMISD0cuwc5Sw4ijiDE543pDo/S/mZNeNHFphL4DwXL
RTKlo6mk8YGEUhE01zMeOI4ulwYJ+RNSRcg1chqXasSuBnsQZUgbLayAVVn1lZ1XvAkFUP9AUTgT
r/4Yd50C4U8UFkfqtaatmmjeENJ/QzdMEPX9SlKQryVXJqXYWgpHPIAb/grHLOpP9HKpW5zVoYO8
47pHeTG1MHMDGOlwRGFAyLcrgcs8U9wXevRIpIrlTkX7r9t2L9SZ8GlfHm5sKR7qx3Ga8WfAVcLW
cJm443+e52Gg0t8tCGdMbMbrTLGcQBj66UDInLgLtDxOuQmWNesC6tMawHXgJmsb9OFG5JR8Scp5
N6PMK6eNC3tZ93dWekj8VAQE3+CKM/SAx4/motpygJxxySUbsrVthT9SiQVB5oWG/JQmZJzRkblX
qkNq45wMi3kht9AUmENmjhxUfXM6vD1of0rol7hVoVSCZgWmrvLvef2twlPWh2TH4CBC+mmWeuH5
HF0Ij9hb6bBYISwZlcMg2vBKxKMN6ecOUtKaaaJButy86O+WvGdRSOg7GCDCkikHH0mh89Wrt7Zt
MdxWSkRpb6rlRJeofw97iiZAk8/eh8Sb/qyYpy7CXWTdDW+GXltDyJefLlnXnl6xMN6lpkHYnB6Z
RIXAhphMhpTdu24ycVPsYA3yqWtW89Xd8fN3ooYxQQDV5VrNBXlbFJeZqh9XYkolDHp9ndBjYImD
/WYawrLWMXXYF4vjQwSVSrtm/cX+skU6Y7rLK3qGFFRWT1TVVaXRcXLRVlW+wOnJpODkiYEugVqM
TIuZ88R8oFZGjdmdGM107Z4T9QkXNFyo6fXl6gM91aMaqiwggh2fb3Yq+fXoZWSuTnEdypi1d02H
OuG1MaG8MRKIkpZLq/2mg8ccgHcWyC75heL3HdFHcrQSbcKise/WODiOTlTj1dT1nfz77xakerxf
zWm43G6GOBi41hqC0SnaDCqsRwdnJGtLKZlqHCuZLbAFT4bC+Ia7ayRWFXVtfRib1midfAsUPFFU
sAmnRHPiPafTzITky/pCdYEq4iLh/M7FxowViVA+wvbV3XFE9r3NwzmCD31YsYYFpdR88E5eMorQ
ol6LZYcwizyCB/ky4crv3tmgK/Y96a6fzJrC2RNd0WIs6Aj1uNTiNMef5dd9WVBOynobg+dWCt6i
MmItXqT9DXXi2swT6oytIdxRgKLLSEW8+dM0y6LziErA03P6IxH4hgJ06dgrDMVYSn0ZbKDCWzUy
1k0Y9f+kpYSeHq9Vwg5aIhriABEg7ZrZbpvPWBfMgSO1FfHz1Vj7Tx0Wh9kZ8klCImkF8bH/d61p
hHDL7tRwwPeVdiqHV59dHBHpd2O28Cr001wzkzxN5Dhfs2jd68R7p2HiWvKav1h3MugqM99R33lq
Yv0i+L4LBsrqyW3fppmWZxxul+uVzmj2mlj9VycgZ+S61IfAq3Mvb8SMyyPx1yZdHzyz6los9sAV
5+Qp3YhjTsg4q9yMRLbeVuhkZPuh6ic/hyZ/fLTiNqUd37GqGMPVxNHwi+c0SEBK1M+Osf8/5RcO
Jn3FqKWvai10XeXUL0+5Cn5WdHYBIvEB4NxB+C+KbHcZ5p3vo68j0ZCBz6CKjv8FHdZ/OHLHQA29
5AKz9cxw/aQwxEBZoggTJ5YkDDVRtayD9RRso4OLpuCj2QvIwqE1pYqzv+V/dSYzv4u+cFxIlBx7
Usay4OR9eA4b1EG0Z7hPTXaDa+lshnUD/6p2haZ6oDnXDgmNYaq9Rw8DJpMP+alTyMOMb7V3sIER
3M9+Z0aw7s/QkZGeLi6mi7TP9dLHAfJb3rD32mVOyuCNiseQq2CbhnkyPFB4p49/3/tYi742sist
Q1R+SqBeDI+qJ5UKvIIIjqqPXqYCs3SYTbh4M1Py6mJovWpxjiy0tOK1r78lvV63zVkD9+Yu1Ap1
sD3R8XlW5if4x/u5QkmHYkrcO2FQFrRac3YaxJZ3J0xzHefiot+YEKqmtAS0GHXCVDslIxiZxS2b
Cch5Q6TvJV1S74dEtwqIgvflRFKtBoeQXeXgNs3GCHO4Mkv60l0mVd852RxRtnpJgSNT1jby+Urb
UdVm6XUUQ3Eoy3QvFHDX3QfMLoxdh3vx6yeD5XaDAT8Hb8Jj0ARSHTBep5GsQyZzRYUhR87Qm9PX
sMs8Bdf6RkOnf2FK+WfiXo1GcscG6kKFcygyaSORGCxVrW00UlzjJYllvpaiSPH5V6/+8fXVIByY
kG2CgFs/0EJ0bcbo50UewCNI3HiczJHGlMz6nLW3cuH1hHVVE5BXW7GiQvlM0Oj4kAoXDWV3ylP8
pFvpibC6HJHLp0S9Yp8nLGj/Qzf3Tq0Ha17FeBFP9BQMNDvxXFRl3/d7WNITjR/KgAxlZ20Kw0gc
yFR6AIK5ekR8L4QBVx0uO+yqwNQ6FhsFmad4LdkCGGHTkkGuM/DR+CykCf4kybH9EkXSJNSk0+T1
fgyyiaa64EYCGlfeoN2wHCtct9c9JFVXaH6o9mcHfPEXBpwFbUCUUSEJyBNkL61JYKmlOe48jZca
kEiORTVQhCa+2IHoZFKQ62ZBej2gSa+pMlVtB72Tc0IvsmUnr7X++N+15+SLGXzxCZyD/1o6E+g5
8b+HuFdnrOZEvVPV431vzez7jsDA41QamQJCswapPLrTvpqHIGjXTw8uhf+wZ2kXIbIm/ZURWzB6
+Y0cr15YkF9Dkkazk0Ld2v7uf1XINQHtrkqk8TTyNHoDIJ67W4NvJj1Xs6NVcO6FqTzwExUjWO3h
c3U1Y0MmUqIldHd6wCVUDWpH91Y4Yl6QSIcoxOZUTRwQM6zCzPFnK7G1J1FPGsHQ196s8VeVwiow
nGVr82N5l5gWTCJSpz3BIR+mwrlj0B4wb9W6JxWP+Obm5qmPUjEDl8L95LG6rpERvTZBO8vDQuvt
z7FONBwxpt4WOxpJMUpt31Yw2M+ckwkNCCy2dztdpHzv/djRlzaKdasJ6xpt0v1EsKgf0/UuX7qE
DR1FU7uHWmfIAX/ECFM3kmHOLJj0xIq/DhpAWMNh1GQ1i7h9DPjt/ib3ZiGnfYta3wS3zut1s2eK
ZuqiBhJeLV/wrPYKGA8CHx6FbXthjZq8Fx5a91sxHomKCDdoB+sz4yJX9e33JY09qzssXrdfYOJJ
6WCnw3ZCQZgxjvn2ZvsvhmpHFVvGdZJCJ3zxm0wYRsbjbA3LrRyyEAE8aC0leL1mFdEJ24jVkGGL
WGy9cwL2L092VVzGda6BwA5jiEEycK4t4cSobNENgCocWKkUyr85gidV5Py1o6cM3xv2x3m/m60c
2a2FbjW9WbpwEjgQEnncL95AEAOVUS6mzpREaoH7OJ8yiInEmbcZfQpPb9dq5pTBviAXPd+Wr9Dj
TsKbE1TmbTI6quP2wwv7DMf7uggJ6AEU0alermbUZuN8Mi/i5E2ctQpAsvXsakrsU+qwJt2W+j55
vQ7avzYB3SUnxoH3Mxd8a/FYLsSWg0bn8mm+a/z2zuVn8y2pw7fxRCyOghtQEie6+hoYm4wED4be
yHd8yjWxdw+skH1SaDampGhz54SFD3qzR1xL0BxoKU8NvK0+5V4EdTRFY+YHcQD0yb5VyfWVRB8M
7e/G1aqJ/vJCAKslQd8lumn1iZW5Cq7qmtAoH41EpA3hLcLjaS+Ae/Z5DkrufG7V96GvxlwAB4DR
4EA4h1jm5iMBKVfTtcYeVeSR9tZsJYPapTRr57zKdTPYUx0No8IMrmd+ZaW7m5gBg2BrfcYJSlH4
73T/1E5KryT6y9LdYF75HuRyoU0DkLEmaeP+pG+FbkwxYJ5JmVEf0lgUnZVdUWMChTG0qG2sS5+k
ei5JvxhQQ6S/RFf+xOtLGDYGK5JmlUybE1mB19mUNR6xeg5lKxHewBD5XbsrrQkNTIYP8thYJn+B
Z1ASIuDVSfT7ecqlK8A9IQcWIMkGGBXDTswteLL4rDj4z3WTqYAfYGL2N8dZa8bd8Qx2bnPZ1LTE
o6SlZzsuuwipDN3prMltnYVn58kAtIalFFKpj4ATRNcQjyX3LzWjTPBbB6oTdGnFTDZ0Jh0019Z0
4kb5i4kYXXQ4P5kGtuKkgDZPdRcKlPaXs7hJh6+Frqopsat5Wky1RTEG1lo8fn8oLbbzv7cEUgL1
N4Z02cqkUy4duv4loo9PbzM1rmBXXbAAVsRSarqQY4s5UwtdYgSAC25gyhSokOvRVjazMUUAa6mm
4DHu0PSGiKGekdC9NwSGAZImOs4EuZDVAgsTfhVTFV8IwA/L/TdjQKC00n2uYI2dhDdMOy35BI2q
N+gHuSOnSF2a/Fk2RKiDnJV5fCA2vf4mK6/PpUMRH5ENc+Y13zWVRmvoNJa5sHo2NJeOca6fnEJJ
F270ycbIE+ESkOSDFAsLp6XkEzddrxtAVXtqLpk5u8wVBhRgfjp5YHfUy5xYz1nqfCDQpgC0qcN1
sqsGm8LwIawqmn7iCa7TyCnka2E4bpWs4vT6iSpNBr2o9QtL27+PvbF9+PbeiTnrK4HqsazfWJCK
b6SKh69cgHheqDr0jWqPBjUEDj7Oko1EgjtPiEQ/LgqjrvK9ee/zI5GsFRrkuUsFwmo+6mCE4f+R
7wn20th3Ov0WxRoI//iyV8olIDgBAhNQuAmGhiN/tzoeDVyDzx2p8xbjf/fIkhA4ozjvG+srakl2
dm7qdni9LPM+M+Wo6i5+aChjDLg2WC5Kesi0PulFkc7u/1IstjlCD1AVyIf5QVLmaCyifd65ku0Y
ccljgiDbq9NIj1njtpgI6K2mCPgIT6uU5ZCvjs4vGqwqU0+zOEHuk57L8Nnfu77oxO1mD7fddtOJ
vUObE1LsSIo53SDJV5qUXFPPQnxNG8pONhw0rtPNsGAREbOjgo3qo+SHjG5A5WtKMqR8nsT0d2pP
hJc9H65PpHxS2da8w8pMf5QGv08NePWw9mYV9n1LTZkjxOpQwTQqQF5BMgoNNwiugb0Vg50wEWfA
luJcQD3l6QSGjGXbALDL7LImjgIW9biN9RWvTTzCpzB6CmOdYbDEQ6n+Y5asCgU472IrvNHIVuip
sUYoAa0Rl+VVTWoqGUUFiHy5qVl0wUjp/YDEtsqByxXyCNfUInSE2oiYTzKVxLKgFEUJ2q1qOhRX
f0hGsZeJ/bFgO//ZJwPgRsKsH5+c+a+7u6QPNlYsGRyqOxO8Btc2h9P79/lDvJMBIXanVG50VYOT
JccQt9cyJD7DWk1twVntwPzrAY0CJOOr+SBzukoLKHb1k2DZx7tY1wV7FISipClSEg9HDxR5tSyW
pM84iAVSkbcZtRRDpUs5cri2HI47wwCsjlEFwNFk1Uujy2lL7tFQTog+ZNmtWzGbQAhHYQ6iIZdj
qm37bLGRcfXBN/Hb7MklscEG92aoMZHRjgosH0TOZbk8IfPOy1I91ggJL3nb00aqvSYVc1p7a8SS
Lj6WL1zdZGXq8kHzBumi5ErY/idp6zNWjbYLAXpS3NcvIp535ZI+5Oj7dR634f8sjuDXNde7Ai2z
xMNA+HVe68GaaHpH8EueEDyZ8O+mvNm3l+BWTV3MglUGmjuwX1MefJi72+E/XV2mlrkQhA/c0y8Z
HK9GeQvwn0J+l0Z8zws1+xSkpNboVqIo+D04sTInSCnxOWBv5asrXh7G1Jv+QLALghVaEpfNgUbO
4Fw8a37Xgm7hRwXj+bpPg/KoUl4JkyOlajBOTSyCPkcxyqbZejV2QM1PM1jGUqimvK0m+gVgWmDP
SPJv/zUqEfl0rla4vKQ7n4thpgLLMoT1derw7TSl8A40m2zEB8rjqH6pLUZonSReWRioIA270HJb
qOIqP03RHVWE5xj9MGIjrDikqeA0b5HtpB2C7As7J6v9Qs3iYvrkSdfPSqICqhj25HgFB+EpgARr
3jXYaUgwpnOXy901lP877N34lzGT0r69eYRp+MuYIzzMoIjkq8cj9MhrQMVYYFh4B+bHcezirqoi
+JIsmKyclINyJkOyx34YYpQwEh/hHi6H1rTkvhJtF3rJLeDo0h22UOj5J7nHUULfCUorjrEkW7/W
BD2X4QM1rqdj+BXQmxhU/aPIi54aHwskT6cpWusSI8evRxCegWrDm5jMyxfAI3/4Am/m/VAdCoo2
IeYhtj3XOVtVCGMal5yyuUoQIXv/S2RPYWvCODSoOJ21GQnzAdD97dv4UZZaxk2/koIs/d9jebPk
V4w1i3AOXVeuR2e1TLqxk0sRGkwohufbM2NJAJvW0oZwW+8Fg6i9Osi4OiisN5EARqP7p8I1UTQk
2/1lgNaNDNtuURDLO8mBviLEnqDpSyKC5qpWOyClTDErNVZTzBRM30OMPdShQQkmDLiberyY8APy
ApGmtTiKofnv+3+7jvc0+TO73lDcpTmD4CIp9rWVkY+lmmY5gGBHId5rjOFcrWpPi82qFRn+yuWB
Ai3Ngixk/tT7zr1uqCQfuTb11LyLnHenmuYSOatskB2ZTlCdCAe3lleLLR67MjFNpE1UP3HlSaPs
YSsDJfaTvSgghXeZVsDe4t+lDFsvOdRNLoovAPbrxhe8OW/XG0CBv89sivJ2U6KQUeFhzIphj3/c
KCdYdPIijDP1b2LaNtaiWzEu78Fn96ymK7kL2rNa7KmCl1pTtv5jf3ZsiWwunDMeoi2NaXx03lBZ
veZZ4BOZBwUOMyQpJfe53lttUH/s3JxeBrKGcqZ/YIu+caSh1qjAx+sYxPNfp36+6QiDKEw36Dx9
MYug0gJ0Wk3ln5BOelSy/DhgQTrU/SQHEnTWqe8DlrM9SkRoPYtN29r7EDbEcHSDoggLvAiVHrDy
8iL8MGSi0reoozG5dKAfC6HD0eK8SLpINIp4fowRJHeOCYEK+jnBN8amD+A87piMwMcZAgEL29P0
p208ktzzrIyD76SZ0jOhGsuJ34q+OmhnvTYSqlAOKDgvYiM6C6OfG+KJERbaXJu885i8ffgKIg/f
Hae6SteiDl/29fUyV0TQh5ousmZvrrhbZcYakSY/T/iAawWR/OD/PGDssctRARXupBBI0EjrAkWO
Cw56bana2UtSEj/d/ljijRWpHJlEZ7AzJLaIYb8ofmXaX39tMDkMvnm7EFgddJO9qpPk6lRa9/F4
SJuB6tKBS1fy8EYzd9U9SJyu6gL9Z2pF/7PRys9G7QaGtzVdIwG9ufKwwDvnG3AHJyI2m/eQbIGr
OhMJar0vCygKRNrq+ZcqMhAU9hPb1jIHzqzxEpYZrQypxNmiCIdgD4raFtCSobbAWD6rCvADb1aI
zBi/eje0e/omukGTkOb7Ave/Vb/jjmAwcR3An9clNJBtTBD/RuKkgcwPW3B0k9DccBpu0BDb1p8m
iRkwfgxu3MT6vl1ulb8AEKQglhnX+2V+LTwYY/l82zQUlGItjW1sSs+HPBVgOTs+PqMwOK9aYDDc
hnLKSY6l0YYTyZ/IeAkjYtdo+MCQZ7IyhZra28B2apYCkr83Q0uT/tzb9rWqe3h7uiTlUgA+rIPB
u+K64WjMSj6Kec1Bf7LSRRpPEK+tz5LfUEVFl/rScJGT3TEwRGXHr0RwHmHiGs2xdjQu9rgPXZRV
vJDoPZaZtW1OaVs5MqC0CGEuV/azSjMd/oh7vURGBuXEO5Q4X06BH34zykczFm5b5Nxa3qd/6amx
jBrnFQo4SkFdYWIVHxEJDQcpAIadiFD/UqqmH/Uhau3eczTkBxZQ4NV8O50HYhQ24mYmee9uRKOK
65+zjHs+odTWfXCXRtYFaJA81vh6IamRU7bYTurS3KWUMAjI50wy126cTz8c5IEK4vMOKQbskYy5
5eMW+VDVAyYhozRGX8YMFWL02WY2gYfvr0elz4oTAb8+LPEEUxJnok4ohb0AbdUidGvMHzChRbC/
oV8xTcMZAuUjr493Xj8Q4Uf5SDoYGe6d7sFRbVBQxNV+Mq7DUJsqrrapmatn7bOWxji9YbmHF33e
GvXA9o2dX62SQdB4zo5GYbjeAfftEZKLRmM21k8GoiGpHG8fgPYa2HTmmPCuqJfnmgo30Ylb9PCR
m2fiqoR7as0M0jTxwU1CIQlpkYqqLoFti41PHa6vBfGU5Hda3kDmafFn51PDiQJHIFswn6002kXe
DFI3oKfngIexBEHz+R1ydbG0XrXKX0RSXGDidQ/bt3Ap4fuRoN4YDtLWc1bOKvKDPdMmcGhBn218
vKIT6B3RK5QyAb4kZrDtzq33IUqRPw+/Aqe5SfoFyQ/3SrtrR91DDUOzx46tiHWHZ543urv/gTBI
LS0wNvT558Q1dO5pYzjaVTxIQESpz4B9S3Rwbu9HmNSY/27SxRfG9yLtbRm+64e5u4zKayUe2fE5
7rupkvZX9rnOQUkBUJ5goi29WBh5Ql+yx6zX9Bbg7HxyPoiHlsLfhx7oCFwep+EtFWYPMOSLCxHL
M12aBONZU8tKtSo2UYBA3x2hU0T+SvX6PrVxXPeWoEn9yIS0hewqQXxVEzmRwgrhCibkD+3hcfLb
Ybd9OxzX9Fdl4/K+CiXC7UkjHKH96nJnzWBCMXKX51qjI3UkTDtvoEVQQYggcYXtHU0KQE/qw3Ih
LiKIAYccmA8j8W/mNji/DMh8Hp6gNzBQBrW/gRC140ALzuWDegBIXgVAELZAhVn34PJkf1jMRR1S
OSgkoj5SefSlQD0hQay531M/c9iyHrRiVJYqSbWxc77BEgFvEtOSjwUhaihwUxcmDFlLP7iGuB5m
I8it67QYqWA+k5qAHoHoGlJw8qb3fTUUAvj85zLBDYIRQbU1FLpSOPgj/j3L0f0eEYKie+EuRsBC
S79eU/a9ObIp6HYbiKtHK4XffbEfTWndXEWIvGPsGZ/uGo/ZGpsJ07dlr4oFs4qJ//LbJadbwQh9
cjluk01ki8EzPE76TTUUwXooHEsFIqdVWGCQMSgHjNyH5s+sdFVMpMm+bnAj5+JNSCUZ8/RBOx9s
yfsB4FNYdMwhE0RSqWlmFBr0fI97qjZ8wR9PvZsWxAVyABzy1pTUZPtWAk/JvcMwTc3ApB67Nblq
ypPFj43Dw/aS5EDtOXbGPbpaic+2SRrqO7EX/wUO7OYQ4cySP6XqIZVvBbyNkDmR3qkcJ8vwnWg9
Jc1JOv+G0uIBp8+IucyUJxzTwUBybWONcSRTdnGVEmIed5Qq3r+bgAs8SRFcATHz7KBVDXADT39W
iQdFaE7pLn+VTN44bB0AzDu6ACwG6LSoh/Vx1ntaPmIxiHs/zS4KSjtd6Jf3NUpAMJx9e+WnyY90
m6NsF+qSqTAFxrZ67aI5Uxnd7SbjB7lVJ9cju8aUi92MFfhQoTo3aLerqLXXcF1TtNMqPP6RuJyU
AMT5Ar0rPGrtxyfg0xgaHxDkKYXXlCkIHiCXq4YUrAvG8uOKCZmOBKvtqJcPzHJCG6o3xGV3XESZ
ogy+rQAmFj1PmArQZOV96YWDAqThJLUL9QhWgw52MrY1UP69IVuhHBZrkny9f8Y35eueiKVJbcn1
DYOILAfql9DOsmpX7kFeLgvc5fnl/a9zgx8x+N3+kRGuIYoq+qpRokgzpuZnT9nNcV+2Zy2Sfrif
Lx+HIXbYBVv7JIdXjXN0gGVsfDivOo+RxXBQhIW6J761xomZA3NSTaPWl4MH7emn37xysBLU/cl1
PmPJ5JTPudOVktL57AbQsn7eRRJYmfJKm30v6hcs8+bB78alFQChldbH3RgDs0PrSMgjrtpatjP/
XiX24qNd/9c8hL7Gux938foMQanzz96tNgu2dKwYwZ4VF5CRDYbd+x+Ng8YyrrDXZJh8ysZPZhpY
6W0yIM4ayVZTedNqpQnXTsXhk1IUbsbWklBl3d2Q7ysVCpugD1DELci9f1c6MJ2WVSxf5c0FoxYl
q3RGyvB6WSA1OQJfQ4fTMgtkaBsyjD6oljcuiIrVLr9ATCTSrlUmjv03z2QNxHA/8b9U9xUoXCuS
KLaZkDMdvbOYn8ZTOmUPKLbbqZ17lIX+thcZXkC5hVkBiU6QcsFGVec/iqqBtdk97avV1knl93OK
suZOZLFj3UQGs+TQ0k1g6HPvXHeEU71WC4d1M/FA8Fb7sNCSI2hxGeVKpVIRtxMZ/cpouyXOmxFD
Ob9KUAhz589dN7S/9AG2f4f3H2SMY54h6mxEMLggJyfC5zyCUm7WEIOU8ZSmINeudsytn1zGIIHB
YOh7NT9y7b/GSieLieROq9WT3G7nFQIQR7CkeVV6z4myToCE+nnIICDD79Gbk5aPoxv/FAhpQ4W0
b8RikrECDO5HF/J60hF/jV0p7XXUr/OL0q91xGtWEjD/aacFS8bOyYpmASESB/hxgsw3rDezaERl
vmud/VUQhine5st+vnpoM/UmaEzk2enh+/IcYfF08Qr78ZFiTvN1eUH+eQ8ueh317+2pMwrLYafO
rQG6ayA6UELx/ckJx0jcF7b7SMwMnMjfjVziqVvt9PuVEYDb6VR5pXpH9raVNXDDIH4AwniO118i
gqk53SXP/1SWVrm2tla+W8MPWgllkH2afm1PoMMVSQgfG3MQjPSFyz8hTfm+VW0EbWYNgxY3V5+e
JQzSfpIen+Dhy1KL4eOSNdXmnn3lmlQaT0ofBfnwxMS2oDuPRjP+X3cKEOJ/D0SfR6v34fg5g0hQ
8qCTEBWYnuXDglXSfgjQXSOO57dwXmDAutsDGRMxs7mbz+MOxdEMB9o90Th1AtWgeoj5pLhU+3Nh
4dBCLhZToIrZZpFy3JR374GiWl+/QVlZNzCpY52bVYCdu4B9RyOubHC0c/1crIVIBxfEwDMkhnMJ
yDeEtNlQW7U/hWq/u5L/z3+dqePCIqctFCL/jlRcfD47KgURGMpanfqedCpgReZj/lMj3K69/SD6
RCG9XUUJcZo7bnlPv50kGKX6s9Rtg8CgRT7FbEpPVpPVbFJnQxRZ74u2m5vmQYBdRPfGu+yaqL9Q
BDuStDs7klxEfrEqPymBZi2efcuSJYzEmhLTdILMcYfv0plE/Me7o6lx+QAMoAdrtbFX7QPFI0f6
kU8SrEZcdQtjXz69ikonQ7SJz0/gft7V5RO6GrxpVRqaVvIf3hxXB4FA7L3tg8GW1Vu3TYykNiCb
qkiaQBtKqLND8/1RPw3d2Cwn4WhIol2P2K2O6ehA3ax7jZ8qbfTUYWmcYX87/keFRyKrMBBYsWvE
mNtS9saerfnjAx27we6QSJjfmUaJKsCNTzCe93nw0LEXTsYGpxWGNf3T8Du1QNA19VYXibrENeUt
QundZuabdJgUh9jx7+9ct+aBO6vmblMKNGAQ02zwZSskM5V8grnvdzbRHZgz6bfTio1Lq8YSxKTb
iTAXqzRwY6T5lCdsDE0TiYfRmgCwh1FYx0GMgQRc3FBAa5LlXWxNg9+m4JP0kBP+rwUfqb9ndv5G
j3Pwyk+WYvOiQhylgh9rGHD//std+WhamKQUg6wGiQN9lwutIZrIBbeS+ffnMuFMZP11bb81xBsH
EqM4XFlhDGJ7TvaeZMONi0aZc0Ds29A6bL+cQTeyThyMLDh/VCzx5Qd557IGYD+Q2ms3KHS1HlI7
5t5l/jjFLdXAjWWtMeD6y+9ZLVnd/w6Sfg5PIQgY/7wQtheKiQBDhv7k4HEtFL+3B9qhzOH9Edxw
wdORy6ZABpgeC7LakPK5VtzKQ5KNmKEYhs2MLLfRMhyBlxGeP3FIeOHkFOdp09qzdyxZKU+ZD1j6
cCUxIHWAcDpo5UW4AaG7I4fOYbF1lB43skAlTbGIS/GxMrpnCuJtnKNQXBdtrwYz5jXvd+UOmVCB
IjVBkb3b/hRX5r9lh/11iTOpm6YOB8sErUIcT9VUFzEglWcG7w+YhVO6tVhbZSKYWN/kbGhihOLe
I6BDIiutNVjwdVH+Ky3UIrvGEtGtDjocOA8Ip7UDFtaBeucuiXXWJU7reQW1eBrhdWAAyM1nIpTV
zmDuJ/TE3pwyLdKxMycpgDAGAixhmZRvGf6TlQVTD6FCl3v7MJIbWVpTH2KWS/0tl+GRZpRaSrv3
azb6YIaRfqKy8cbNWIpwRkvEdnF5FfQS8hjAtn9k81fG60xz8m3KiucgH1XPfDj+W67tg284YuWB
DcFdTNQXzKcIHGuP1QLTLOjSbLvsFyln1aGbgHGLrCJr0IIRxRzdcuX9lUITOx5RNxFCmAqCRpUD
UgbZOt2z6eRtZOtdAVM4DVBdFRNArKq4s+zcWNdCfPy3QcO34MEMB2pLwmU52+ifDdAeLC7xEpAJ
UdYSN4G9aGgf6fYNBVc0VZNZnWbZls9t+ScWCvXvxr3VD1JMTHpOYQ51rF6cgmYE6kfeb6eCDUTt
Lo5LLQVIlV1DmgjqKyTop5bZrDogVSPTvtflh3LuBV0ijTvbnnd7ixrjBUq5cnmYkbsnn2jgo+Fm
aA5Pxl/5uQ4/K5Uf7PbznM2J+2Hpf4GluYqnXqBOg+UHr97W4SugRdvTdJdPCAWhpcsKDQ5dbfzC
sqFz2AHksLIDv1ftB4Gq984gP3nrmHcGVn+7ifvcJw8X+E0hi1qV1vCIizLgvNa6fkGnSv5AEEuH
9AJIcKRo8+qiNrlg71Qd1gsqbJn0vn2CBbt3jAxVWtp7eXEgVxDbJunxMe5jAVyJOaJzS/LhsxZR
C9wXtrtXJkwOZX/y6VXxLAMxzVG2KK9rKjR2KZ1NYvP4d44GnRAKb+oBE0AdFHEAN1MKxV57LeIo
v2QROPQp+lhQtkqISveAOOhQDpl0zpw0HicwhVf7O4BbDv6hC3vXQDSyXHJGzrT1Yy/W6BzPjGya
doqOM2Z9yoIQCFFmt32aSP0YLTncRJTwbpirc5z3Rl9FFbHn/tlky+sp99cVyki/EBC1iruhTQh6
f38AMz0fY7KAbTKWZ2j4oUmze7gKzCUkHSSgL0pxiGl2VXQZcDNW+jQBUl8UrMMyEpImwfa3uMda
WyhXtQRjse2T7v1Yi00D78WblAWvj+Mr+FopTrVijKsgkbGy13Kb1PiLSHTwbbAxN69ifXgRCiix
DQXU5gt2WRuUoAOLTFElNwpiINKw3cm3NQOS6dO3acr62ij8kpktnm5GPhXFAFsEuVybzJrgVLQY
v23Xw5yEfbmf4AqfrAvA5VH82SKV3ldmYSV5H9tkS9EcwXZC1c3gojAEx2yElcKkNCwOWLdG6xt6
v2VIGWeoiZ8DyK9zn+0zCrBk8jFGpgM/zaDa1S0MyVkIvR5cD8KfMIzbqVn7eO1F4dza8pL1Lcaw
/vNaj0XWwk6DfJZvr2z8SG/L3OzG/6lYCNKOZnKWdRWmiTn/wuPKCKeyEgDU62wGLIuz56+37Kbm
2zDxwvzLAY4l59KQ74KKPUmEgvuFJ5pXv9Jp8bhFGX5d4dY3gn6m0exNGFu+XTDmxpJtsCsZQQhu
N5GKQsjtVapTTXWoChDYE1VWRVBRoGLjM4ExJdyRtHQUwb6wQYBiKmvNlO5fFALIxvCYmBGGEvCl
F7xnvOcjdH0XVUy9GHiTDIyQUk5tUtbnSq9yqf60uvF+uVFo2p4EW6xXVAMeNkFg8+5VN5j2SyYA
hPX4opCkXKGOqBXvXaYGqVGtHLvxHEdrPVPnxVo/ZGnuolr65GtlgEYjRC+VsEABY8hwwrIZXDvj
D1tkKFtjthhJ4JJsnCpDJ5D9+g0bWR2cTKPJwRKbmA8AEQDWSPN0idJJVV6+cK2yICdvVWnuKYm+
M3b8Kw9KdQful6+RHpZNW4LPbdNUKW5Unywj8Rwg/OFOiTQlhV4Qu7ooQqG6to7m/Km6sgn9GVS8
h4k4tpyVI8T186VuscQM52E1sQkyN3Q35WMpNo1+5jPJ2Tl1O5e8edoSBaO/XMJVGuWztsYY4QIz
BOZKn0ZUjKt6EHWpyO0n5hXwi575a5HD8gClFaT81qNChf/K54i/ZLrAz6c6owDPHm1XHqTlykjD
visemz1m7tLNv9b9rUEvW2FEVcaXf+cDpQ8lzHt2qwbkqx1aprdklnv/VFnp/LFM9b7Qa0coDVVN
p2J5B7/dtdmvf2UDGxSL1RXYFjFWdo3cX0xX+ohxEIu6wqifrlJnf5DkLa28OYMX//RPEVysjuBg
B7ReRBDEmZGQI7lGr0biUaNzEmW4jfepGyUYx0NHAnvhZZejxdwTsvR5L8jYO/ppGDBAJfmb7tWA
EvFW/ToMP1RdQxMV796deIJ+s6+fVEmqRgGrWOya7RPnmdCujKU6zTUnmOl9Hf1TazEDL/LNcT7E
2pyEbcXxNeVDo4S11OiQvya9IzZUOs70wWB9IyH9YWweamKF9dJh/0USlT7JWU44jrWrAA9YKoPT
BsnDdUMvPUYthx7T0q52WA0EiR/0pRsyx/DTMgm2EBOmYh5JgNXg97/AkPTUDwY3kPskN3XJYAct
f60RyNAEwdc+JFyNv28YKA28AXyqXZ1hfIEByaI2LrSK9GA5lUTweAL7l8aUkYLxjvUtiDluFdsx
dWHXNi4lAnSGMAVWLQIPb9KKRmv45ANmuKuXXdyXyhyOqooYYYykxj1cuPg4uXRwmjZhrI+OMg+7
+u4QIREa7JLK3TmU7ImJgzLgUqCh1VhiREJdlG1Bp5lb6nI0Zx3LZNsQvFTRmLbonZkLCUv+wSco
JsH5g28XTEJzg7Web+qq7jKNNs4BcXMCfyieR6+Io3QMGsOl6JLimXZ0wfDAX6aRXOGE+1gI9oL+
PTfuS3N5DoGYP1vUTC07u89BwYj9ZsQm+DCQ8J7fb509OZMf5TPiobJGhI+XzQRSzQY6m7z/1icD
e/jFSeOcV/zrEdApbOlmQCgcAl4HX/s5VbJFkfHcAqrwF0AU7H+vZ3M7/m9mxj1AlM2sxbPkOVFA
LHGXhZ7edAAb9wSaz8SJaAZE5Z8m0F1SEJeLVSQkMwMN/LyZZkgGEoMG9dZoBUZliJ1dpfpN9XW+
n5KBaSnwBtkPq2qHnVbPI2CvUgWWtrMurf91emZ+6Gm6gYcrMTWDeLy/DTQ75RsB8CxmDy4pd6Uq
CwaiRPRODT6GQ0m4nSaJy4JlzaZA61gXbRp1IslhjX5e9nlwfDNlzazmCiNLuyB8y7SQjsZrGCTM
evx5r5iCYHrQGTDaa1nFd8/dUXz2xQVIwNUqfNklNkpkJOyEB6/c3P6e7/bdWi3YHRyLlTqSrAKt
PBzjZAb9kuT7YCjP1HIDqBk0O/znqe+rYm9WRXf1htk71Ed1SThndHhxWV9FK/VIx31FCcCS5ykG
PXeGBxdfXXatUyoJ7whTW+vfyzEgDxAEi5hfSg7BOiobxFJAOE16pzrDtyJlliMQYnzzes046BD0
uvVoH9vmPUiexZ7XrRz1gmmbV2wh+aqo/bzLKL6cWU3zRFZxBg3eH9ZTYf6j48Ev6edktUUHT/nB
TAGjmc/jewlETv31STRf2E5iCohVlPMaB0/qqUqfey7MQ3i1uM2OL8wVFJvY2vxLl+7BJJD3y7/v
/MEs7i3jsVw3QBH8k15JFB1HvKHRpZy5TdUXkfB/cR3Y0nCgmrCVmwoaSLvquCuICditABngb4JV
0VXBdt0+R2nRfgZqgv7aF9fCVlw7j/6f2X95awme1bc2B4Xf561OchsxFTWq4OH6476Q6t1qypAr
W7tgo4+W7joD+GdGkiTJGa5lXeXn7C4fdOc6cETP6pYIMIUJt9q+iJQ6KC5mC1bVUBbSU2bFK2ue
eyv+Bo/+pj6ClfHZciqOQ1HRG3FQ1zQwsqqDztUzX+fMwMA7LizZ5esy75y6TikVycd3EicfpdyN
lhlTahhztnW11FCPLp75pcascByiPBFP3K172jw3faCy5E7SPrD1hA12htTKlYqDc6A7UTjuwY8D
V0jhaFGnUDHEI0Do7yDrxe3gAjH4IKcsohz47jXcRMooc+01M0SZUHdAZK954xrLidumFFkDVXVB
Y9Ajut2Y5goT6j+5dwFTTaio7gIRI/ZC00QwJsw1oiu4IgSQEJ8djtxlH5QX0n76kRFOiCAS3KtP
dAEFgD5+t/DJskmAAfm8aM9pxsZJbwCro+g+VID+fY96SAUv6yc1gD/CDujMalMx187z3ndr+4wa
xVdHBDXRGu3H8dixu0eoVCJAtQsCMDEnZIXSuOggX1z3dI/L0TEa26imX7k5s/prDnIZ1gmbvI8V
W5e8brrq1/HC3GA1YE3QMHaimDKeDaLBbtlVVQ0v2rNf1AW7zIGfT+8kZ4J2+MDm/KYD1F6CY/v8
lpvm1uTy8ZU7dLZk+02d4OOoW7n/DcTS4BnTq3Kw1SjLswAAimLOBgLxAmVCaY3wfVIkdRjJmTMg
0K3d2r/VNuv9qf9OtChfSzts/voI6iRg7kUICD7S/BqxU+jBim5XwEUr/tU3TAAXmIBJLy8uiDTs
iNXnSd/KMVyLYEhU1H9mTgnusYivUW+7tOOlVyCKy90J9ecAJnG25Fz2bZQZ22smzZKlJWKVy6g5
3dw9Q0n7fszdtlMshmGWtsSk2+FEqT26iuFOOu0AQqtRS9B/paEiY6IOTqkkBOzKdCbXrGRSbmOW
VZklYAt8l0sEu4izyTZwxmDC8/eVvaL1GGHKjk3xse/nkWaJT76nAJpzOAsjpCEmmVx+m6JM8Ud/
5lZ+dN/i3ixvfSHNCGUksGv+liej7g/1y1ux1QCC+KZz9HfRCAEDgAhmEunbmbHeoETuCsHnCuYl
mS8hNcV8p86rZufls3S1TL7f3ncon2UMQZXK+YXpsTZFtM7FpI5Ab8rDbfAD2xnjwWVXrnHQzSLA
NN2fqqZo/hsWoSr3qJ4EIFrbKfn67NFauMd7OKB6Ip2sqpeLxV0D3lHsD0jeq7A2dFgM/QBnXh4e
g71sAx4KwquNb3Qv2NVWhoi1C+NRZ2u1iBTnCRlfAk9cuvvU1SCkUqcGEw09uzIi3haIZf3R103Y
q2edu2BtUe0H31BvdjXLqrQg3SzGqrQxK8L4bcn6IkxEVILaIA4dsEl8qUgOdin02A6wwLRprBNl
VEPXaAPKWjVDn+SEp9hFo/7j3G8MocseJRah5xiTWLr34dKkR1YMelscGlsHMIBPmOIBcmOrOjtY
fFgCnlvVfRari4NoqQtjgaTcBJXrd6sSyDLu8XDUugq48Yqj3ELFdLsGiB63wZ/oQwgm9wqcs/Nl
JTOEaeQYDOe+bqIfc5NGaiQbFMpS351yENlwxfhRBmd5l7ug67j28oFyrnbXVWKMd1vZ6Xoriuo5
9Groyc9n/Stomawm2ra6v2IpwXUv0l7lAWSL7P4oi7vWr0xjwJaMAVzK0ofziQ7T98Ob7PwJzc+v
vETijbvZheWWUcZ6DcA/gkNS2m5Qqw6Sm3tTXFlaDHlrsXOuF+X2TH2BCMDN/Wd+kYzpDLPmETNw
Ss+ixYTA9kmFg7UcUKNgfx1Y5b9J8nPH12dqDJcKQrYjNZAHRkxev65rq0vVRtSeNhFX6XLEhvpC
pp1/FSiKvo9JicfJIlikEmmAE+ySjZ6QauuA3vKeZK0z/Ql5RFFbHkASJIAzKQlvGtTZxHJUeDUz
uj4ZEhRGjc/GUvWCBoY5CB8ckv9kLew9qC0pXrI5zvJL7OtG9wGt8RJdmFo7+lIptaw1xq4VmQhq
2xO0dbc76Vz1WYMqoTspw28O3XgYBQW5G8TsmnMgaf7LMJa1RBNJBeVD40Ko/383q5eM5BuAIKZw
/q5E6FqvqSYu1RTwMMekjLx+9QvdJGOYrAuLptzKi/9FQPbxhUoeS7F0yILB7NNrCpMiYC0NY9LI
FPmB7PuOq0eEdsMw18P4uFU4VcoarwrvZlilOhIL3TdPsrOoo+IEb069oIzx0ctnP0ZfrM4v7ak2
av6PsnbAftU59Tt2m8hz5XWJrljRkWKeZlhZW38CzweA9YW+3vcujdTfHDvoelve713vIp/KPQSn
gj14Yp6Jku69RMQwomBW4O5VXpO33QvNaqvGbbcopqfK4sjxXr3dakbcgShtEbDl24NVzA3iCJ3+
bCU4P61M7zHcaBB32zdxcDlei8lWArq1QTX9ZhXiCaLvM+NueSNBhvBY+UJmhPkweorWmqAFvtSx
euBuFfpJsNXBq6TZIEAXkfOaV5dVH8tV/MfS4bIwxGWdV6bvxflRGJ9V5RWaSlLWWgtiDRhRfHXf
ASfEXaLhcWU/z/km8UqfP6zjzZw4Hbfb7NWweu60YdZ8G5Y3HNPKVjNnb1ItTxcVl2dYRIGr3jWg
y64/Rur2mCxO4gfFZCLLio99fe5pqQOfIq8ZLCgKBEWzUGe1hEt6gfuTdltqGofsyLgQFDrg5apm
ov9Va/5KPexheK1Nb11Jn7soyiRUOQjGEtQwiNv3vdBHoElsUabCiIhy6eQv6Rw+breocmyPQQwe
0eF/wVDZgt0LBdtPik7RdHPsu8uj+FP2q7T7LUtR/DHvvpToLtzrzCrx+j+HA+Txdu9ofVtjfmkP
1BxlyPaEmiDV6l4rxEkJ3iyTSxyvwuz0eAlGgU+ubVsfdkfX3iQxV/WTBSnPhXwJF93HHnO2HO+t
uegdEOeZpjlbmMW2qIkmPCQJquYUFM+DBOFv2oQNAZ5VbfoHm9lHx+JnFfBjVWmYKqXFWNFcmhAG
4GBoNep2adGoi0pzsxDtgnMGZxGdfQW4OD2qriygHZ5Qw3Ygcy3o/fB01sToefeUeksD3+KGh8LG
S2yILfu5dZ1iIFjJAFlgaeuPqjPYCaZ0KNCaD5tLacoyBWLnzIK/w88brqXC4vATdAfyqPKyHY5P
sF9EKz+v+kXeRCXZ9VtP/gnQqJTNTOJZX5M9+vmdo2PYXUMrR3kOqjfxQuI0bHOs5dQQwLEycE4/
4ujQMHYYJ/f5SHCFzRlHepZSkhe6G2lPgMQ2LxIF6FkwvTsNOz1Rk8G/ZiCqSQQQIC+H52Da5qJK
TFdm0lOxoVYL5DrmB3eZtjOiQSIV8CrLJdaBBBAfGewJ0tt6L517flOjeu2GdXaOSrXeKHPbz10N
Hh7Nk5T6pJ+hjJ7N/eRs0eV0SRz7BVQui2ylp9IVYkolV6EPZGaQTyKr2qpdgAHjk9sfhqTtlqc+
eYSleB/rScUKmhUIvBNG3q6Iu511pq61BwZ7DIlloTLmedOXy+d0jEgBidkMN5iUeZmmzdajsMuP
5eFyH8rEArSgEVVYYc2C+sz6zJZ7RJ7SOIAgPR+f42HJ8qKohPnB9w00dgK1xs0B0EajVNB++ntw
E0raLY8UVw2GKnEEzTGFZn+JsIdx52nxhzxhXeHqnuDQfqqCneQMJi0EMqrLQOoOR1gmBzkWCVCh
BHlJcJA4yjwhmqe5FA1K5wCrsWFdwWBkKhhOnUr2D9qPNZIu08rOSR6yn4uW4z8kILT9xe30HA8X
58sskfHtjz8Kw7Pkswpp325ND7fkNZwXQKqZfzxBiMSKsSTW8tY66F7+/5UTUhytH8rqYgmkFsNF
/l8DnI+ZMHuLdpID45zhOQLbxBzxIlb1q5DdvvZ5QywfkO9vAckvdIndC3bJuOESfscZp7AdA6Fs
MgXm1KoLlqeI+YreeR7zC05oA4mxqFveKzNIoHdkcfi6ufypBtkMo572Od95gg7hLXt64SPVGsQ+
kz2FG+sRrohS0boZpjEl/CdzrTcencHvoYvDkBIEbRTzl1ByqgV+SsulohQ3RP2U9j8xPrTFNixW
MC0Arz0Jv4pfkY8Px0QK6JZX/FrLYbzHbYI/bj6k6vFV9jJ55vBjDaQKAG6bcMzECjjkuoSqwLR/
3gqOCHDWGIIchSpDsVi48l0sL3+uBrJLPVpYSc8hyvYjUCXX64apTUNnBkvtX37Acp323hwtt3RR
v3keo0mPEHjSpkPPfMyUQ+vS9xhbzyoQxWf1/QdPGT+EcvZcH2lHIRjV6mbv1QHa/H7YL1jEO6tY
6WBX/Wbe9H24pOa0UeBZ34Gxqf+a16OKrlkv1Ku51dVlOxI9ghGwbZufXe61MdsMx5/UwGSxyCVb
jF4K6tGs/3CVaWca/NQ43fVaJ8FVKSEuCAxRJtozTQIEZ/aw8pX+5ZR8cDdIfeP5X1DoUblEST1Y
N/jEX6COhj0IB8flrwRL87DeSmBlRVXnY1kpP/ydu1kkoT4VG6i5mItLO23iDyx5hHzZFTTjUqWY
w/2bNLuXQvStOfW40IprEhgspb6U+DnrgVrMDyuCZl6YnyQHXm1nRpYwm08mlGyvC6SSNAlLI97c
j9gUT+ErV3PZmMU1DEPCdKrYXKt5zSxOB4Yko1+xVox9iXONmsV9z7u71ZqzTZOVQOJ07x61ygiC
LrLQ28/ZgphsapcO7upxgrmMpqFlG1YeMK3tQYR4z2g120qrO+EWrqRG2DDnk4fxtS0GnkVcNxup
o+wOiwtTx48MRukP45+5mgqNe9MOL19PieIGLw+MxJHe0USQMVDYLPzlUvf/CNyP/+8Xf5wfr+rX
W4Bcwd1zhIV0c3kA+GdX94psNvVX8giDOKh4liDllwfQLiz3SHVgW0X6usT6LMfUysvfdOxafMOu
s/AfjlINVSxjnPjAPj3/Zx4yDznKFaphzDq/MV3UrtsVgyBjr8aWJkhx+BNxFOm8jMr0x7QqM7Px
h08W/fwsi2pTE5E2zZqVqSKqD8Pyvu93bjq/8KlP7ZnKN/rwD3i1A83YmPnYMgprO7G0hVR8zrHF
7xkzZOivstapUkYbVvwL1Gy/nF52NnrC+qZhvNVQRrHQo82kFaYkbzBw7Kn4WXAxcZ0Nvt2THIqS
IhyYGB9n7TElQb7aR3MMp85+VU9MlsNtsmeJaqsrxdVISCRmDcRXS7bg+ylc5yiBIVXKzoM+nfyc
Q4QOXP6ibkqvsX6jztTQLS+yjW0Bzp17hCkjsfCTWm8kRi3Vfe6YZm4nsg3Z0FUj08PEJGkel+DG
1IvZlCVVmxVwmMO4rfNxqend/q58p+iVDA6jhQyQs+zcsY7sLeBdi3rilzVsFdxtgAIbPCB7z049
qxnmg+jV+1uhGiiR4epF5e46fHKF8a10E2CTa5o2UnC920XSWP4Y4jHXsZBz3mcbtI19Z5/rCU7M
nJMfRCdfsSxVmxl3i4Les9P6uDc2/Jg4fYu4zDeILlXMI/g8rFayDszcWP5+ygmCS2EhVmZRhRvN
CWJKGFUg4YksD6yYrLHPnHYTswV1jKJCGFijTLYFgzfFEJeXMsDVvBICrk3nbULnS8oWcTFEKD/k
I1Z395pAQrr54xjut+qWnPO8wnbE2CsqOxkmu8DV4D+nTW9YL00SP3tCFUkdBkvarneDNkuFX5m4
VHCI5u6yXBmlISmDKmgejTB9u5tG4MnqEdizlu8Xa4iSs7qPZkHgvhOd5yeehLotzbrvw1rPoPY/
uALB2SA3PwcSOStn5AKZ+8KUk+kbgn0GgUXrEg74LcQncRMwYTmXXPvj7QVijl6UKBfwXiCjF17w
9GgaWyqbi0/1Asi4qy0Qmt7w6hR0IRPEGfifRCLR/Fu3PpIH4yeWo8D01lfE25io2HznHujCSSmf
1NAEgwCtPTHu1On5wpCgb+zQOaAUq3dWRRMJ5Z4puEmHPXv7wF0sg5UVw2DEzqNypOfMt2jknzDG
ivK4ubfcX4QZfDwJE4CAzOBe50JDXIi8mYF1DnDcd9vqlHynqlMeoueHJ0NuUU0nTtvnGC2DOpqt
ewyvS3Ai8PGF+frXDd3qQKq5jpshzGZ3rpxpVXyjGGgx82MoklgMq+8sF8JW4x+mCJCvNIJQ8aKE
9DmETmcz5OUXOvI2KwGV8FBAHsaQpdDTZipQDSlCFXtVXQO1NcFCcPnnMGDP5zleVdjqCXFFoJPT
S1xaGXgJodJEirp47gxr6z33D9lCTQpCCkHTljJ39aaDcCwTkkwshUlr3EI65n1qDLov4Saq5v08
afE2FspSqXTXwY3iPGh2wOGqYHUCWUNGkg7qMJUCddefxLFKFQVmLyVIsVdUUbyr3uCu5kz2YV9n
5R/B2wy1oZaOD0TBYxPjgN5dqXrvHKLRxIJ5gD8PLTxKo1yFXPPPGIwY83i91mjanHAP5Kj8hfPQ
mrmPdNxaVToe183ztLoj0Pn2YmcmmqMPAm5NBI0m1BCSMBMNjFMM5aN8oc9c4BT7tbP6CTXc0yVN
qF7sIweQ4I4+iAzari/PGaISVFxp8cy3xUAqXyhRWRrWKROrZ9JsQpe17CzZqVhWcSwzz/Fe26h5
aj8zybX+rpkjde7wQ59odKoskmBnG2GqPsochI8Rc/adFKUYDx+WCB2YZUzlDte0ubM5yVHR6501
ygoUxmlvlD+g0f8PWzrKo2p03sT2RDXUKAUYnYhVKO3HfxZjv2vKu/pI+YpFHtjhfO47CIin37D7
GA0ZhUv0NwlUtYBvN0h/7n1u81gnp6+cKPbLPVcbXKi5m4Db3gFQ0IfU9DS/17HxqKxLisEp70B6
80XZj9abz2skPyUBglCxzWc/cMcXT5CZq8Pgsuq4667azd61XJbyI6713sJeAKVIm+NZBu2xJbLA
7ZEbf3wcXo9D1lfI509wNz0tsMEXx1TlABi1ApIsS7VUsFrHztmqkStxAuSDjp8k+lwfO/IgZi3A
iLTHr1VOEXXRvii2fF/VtXxiK2mIGjw0ACRJ7eiXuXcKnhsxm7cmADgcKYCE1K6TdcQLFvuF/Qdk
jvrD/pp5PS5LEGOBDfiXJoszHvGvNTiIGhZauIXI3WZj60h8br+VGYZ0zwm4G+dxuQXwelP/VBES
KC+lKiunzGvDRZXt0ZOtWTHxpYutECB3TMr69Z94t1+LEwnYeJl3D9J25cCRH2C59hJLJW61vYRl
kRvMOO8Onu3Kzwy4JDA3YRvMZtSiIJ52amOisdEWIjonkwskEtLvuMBIMuVthizzDM4E75PlTbDK
NNVB/QuHZO9qrBY+DUS5t0zBrhe+mfvM+sn59a2pyMJHjerML2/OEb1rPilSqi1rrmQnFTbZN1yA
XukMvmgkcaIkSqDUnyIum6SLIumq2qJVbqZIFXmFUaeRZY26x7Yk5yTIDsvD/8pWUVvIAcKw7ARO
b/Fg6JkBilasu9sLrGgbKw6JhnNql551LPxyeYwx/SSDbjMpi1mSgu6+Mp8rEpHOlIYtFopRfb6Q
8xfYRBLiTnYfP7ZIfalAa6r3MLh2PFNMzg03ZmJKlXF2Qm9ox3wArl/XPxhFoC5c+ti9psYZbBsB
/tD8d7oKqQobQmfcx1UDLHhwOdky/8KB16o5LtItOnNLD32bJv/vVbKBIRK5Vitr4I9J+HWYKBfw
i5kLRASaqN02sCR+Y3geh2Y30Sb6qEm99d6fZVp/+JMIEmzYgBSaDHERtB65z+sxaW4jqDAhNIae
JbVa2Zpiw/i82MNSKXeLGWuZHbReCY/cRAA0GYyzvgyrc3C6BFEvsucB3MXy00wCYHzMUBEk2tzd
h8svMkn7G1i33G76NJ5hN8BFlKQl4uz/bIkS8cVAtaSYxVTrZkLUqBTFXeSxRGp7NPWOeoeE5k+R
xJjXTdpmdZ1WVpXNNGczKuvzNDTsaLbIc3UO/Yme2PL9x1pnx4ESXXFLkWsImz48ZKgYJLM+e8qE
Jcuo6luY16OTYV8CGcRLCzAolGW/osXAKH3SpTeuYpUUzNBEfOSku42cgKLUKKZKf5NREW27s8FS
ncq9jvntQQPthhx4thvLyIO1+7KkHfDOfXABhuKTKw5uzBnnlHYmCC6Y6TIYSxz9unhiouvIZlnF
SffTZNBt2h/ok1V9ssvEWCTNB9K8fnN0Y7vxvyTAWhXRxA/KLTKkKb5WlhB521xwg/rybgvIE1Bs
UfEmsLXCLkDBTljYZ6Zh0PAibwGSZkw/4JVr9HFSxKjMNQyRut1KDPomTlOXN6Z85p7WgQm8iGxm
+b/yQSHSn2zSgWQSDPNzqNHq5zRtucFQLGuG/U8Tp9S7TRlqT15eKIse7qEU9M1r55bqfLwTRLmR
eO5sm4t4zvTtB6zWY7enXRAWOhpsOOg9li5BF2ZeBvtHKiTHynmItaHsWCCidLJYUXk81+d9S1yN
Y2T5ypZ9JxU4PTpLJuCfbJI7sAmcAXKX5hxfS3kUlKmrp2ZQTqrL70lakB7depYZxXHrTPxjZUvj
xS9sndFpzXi9PBdpy86jafdgOfDhO4X5RQChEsCAUxlK5EyZV90MNzMQS6lPBYh1//Zj78ZqfXg6
FJPr0bglpTF+MEd/AJBIOjADXv1vcDB8RqtLlWnbR+AF4WCdMCCpEIq5kcNyAEmDMUWghdx9VP+k
tYWD+fMzkm6Ohe905ZndZuUwdB65nA1/EjSTlDsPl2yml0cYPjEVLgYx5UdGtiqdBqv8Gbrx/aZc
1crYxRPxlfxzBhSmWPtzi6Cbc2yCf3SUddaBVQKcmP4xuop+0NyYlYqLARfhQIJESNNEoTNxkgyy
BFBGtQN27wEi1ryNE1enEVIRM7r7dvboQO5GxL+3tmaDHbCioHHglEPxVc8zoWWnzYs5DjQlWeEz
rX1t8e9GjIFM50DVDvyJfsYHRBxDUl5JYvm0xVNmwb4+4QFsl1B6Tgh/F8iLlyzuGUVO7QnZyXxp
ZpjE6bd3HksPLXDfzalmwRHniAdNWf8KMYLdFZJUs17SF7A28wfctdVY07+SLvKqZPpCiYlnTjrp
Zsd1oNwiYnmHa733oiSm2AocDPUdUnetAfO+8hS+eKKPD5GrHvpNLQUFugK9KOxLhIuoL71WUgq4
pxZmNp7FHj4MsTnrf2Lk0jNGOjgxlVM0hSfMAdiybkupMhvoYEB9YROKamX/MWWw4SbatDDuykGD
IEYhOH1cYbe3YPwl0nsBTsT1xWtk6QWaQiL33FRHWf9mXzMqVZjLSZWfwL4v1j8rbYS84UQhV1zW
rMZsHoa7PI2yxhbxKRupLwnv69JzklPiIg1z4ABigeSrbocwsakvyrdezvnPQkZrIYwnqafxLMSw
zKqHDVIqsH2yOIm6zw8ttY1yeGXFSNg+ovW+5doSRvd/PEDomeXl342v0l05H1ZqElu4kzpi8Vrn
FTIEBy8GAC25y2nwMoiMC2QyiuYSmkYjKQF0vFuh1Tpky7xg5sBOLYmP17FU50+rWFkf3p+cLhtq
ue5f757CTuMTGsb/VhXR9IO40CmoxugII7zfwwu/GyLKCm6uIj4iv1hA5L1tjXfKOvgSjro42Jit
qIHo2sRg4u6XDMyHKNV7pFYoaNAK7iZN1Tga9+SVBD0l0c7JotDFprY7odtd8Xw3HHO2TcJageKY
s2yWlCh4/dqfbYLNx+1/dGq/Cpji2vl54fN4Pi45/PHueD0mn4+Cd3im24iQ4SFiDw0bjbYevJ25
EuSmEd3Kh5GxKkFB30dV8H/sM2CeqIK0lxjkA/hZR/VO3gXeh+3M6NSf2QTeDANI3YdaKMWUisJ9
SWm90cMysFPsiZ5y+W2nHznjRXHg2dOdhHztSJBYNzGiDNbn1bKOhA74W5fgApc/FSJ5ydAsZ9dR
ZVJ8ikmcki3cMAp6fC05sy6giyCE9mREbnYl5GZNlt9u1uOnSApz3WNkjWQgg7ktedbeGIaXoh3o
CIORX+7xRDK6c5iByylAcAbVjiuuion5UMhZrpVsJ7eLjf4TgwgyoB7OuOPEAUl1I++bLBpymNK9
YSiyXCDKLSxEXkgCP/Bow2ofyaInlEgHAeN4C5MnD1/QBhqCvUHphAKe5gkR0IKdmSiwI69r/Ugx
zr13v9FFikwQbbZAG9ee9hhdc+No13EeeL/BHRqG3MEK55aiBtXbhJTMFXbyjhvA3IIMgbKtAMUT
FNpFM//5NkRzO93G+nsufCDShs5p0o0MROUFzx3zCD7T2cT6zpwVqPTM7mwmNqkUypIo4KSHXl4w
A6zXbU2pcEY4rClNIaEMFlabGxJbwGrJvE1rEV8nwchOesAw/IRLvyhEyMRzd43KuFzGxPKFQO99
SywG3/4SO/7/akFEZ0R5DdbElfdIr6o25iBbFxcR6m1CxAxs2mn3hb7aCR4lxyED2MSWJ0oUY4q3
tSWQ8uX73HzMh8LkN4BgTETfH4qXx3oh8mrmc2jxAcG4A0yajVEwGfQvfAbpvtI3SB8J5u/b5sdC
zrh5w6qKM/hXtesggrN7fSUsQUdG3BDOajgfyomdzdvfL3WJkt/w2k9nBhO8hTQ5CmsnUB73OrV+
/oRYGSaaH/rPUEeehnczjfVqW9l/DK68Cikuafym4H9hPtRR296p29zU64rr5jUMII2wUpu6wu9M
f784Q+noSzhs7Anni3SprKmB4OnBJhvNPXZ9TCiNtG68Tn1EyiNVPXj+ACO/ibr1KIveqQOVZ+K4
mH3VLezYwJHYQYlAqF08Sh6Eo04eUc7C9dxYurHhlQM5JsfM62ybVUAMFhJLiP7C6VVOlMriwcJg
PEz3TwVQVDW8wtHFjXUDeyU8QNrskYfUzDT0unly3ih8hXcknRZp6IHC1FfwGsgX86BzcQJdzZOj
eCk0Nh9bwwIgaLjvu8x/C36e0yTjpPWA5uz9VVobbaR9N/1JGrG1Igwx5UoV3F8952VUTIn1ZXK1
7qJLwbxMgpzkabdUDBMLZbFY6gcZRyEC8U34qs2Cpby3kvSlpRxxyZxxvnsaO+mjEXX+5Yu0eZx6
fSsP4URy3+3cb1XUGhCKeeUMukC0xF3dY4lanHcxosLK1X21l4yMjONUSdquf7wkvWA19UNMAwkl
pIWOWqRoLK+0lza5u4DDYM/WUezUOCx6KMSGYZ2Dnrx7AeCZAr1RoiTR2y+xyvHPwpE5L6mCqIwl
5P34VUaMleC1WIns9W7pcvVZa1/tUT0V4ptP9iDdwbVwFkFHsum87VNfL7lQd5tanfGmULNWrX4q
9buQ6zK5/PbmNZFMSDAB7ioTw+mkpVuGk+ssMsG7TzGsKvS8Q7P2LnfYEyKH+AkQqmqh6al6iWg8
GPUO7iIt/Ub6kbhratY7W5rsI0UfgwmGbhDtks/Pn75x+hiAPEUCMITGHFBZKQjvPa7RTu3Vrp2L
tvcM0nHGdfYijt2vzcXRhx4MqQt49mJRl4pBM7qn/KbqzZeRh5as3CKard0l8eG7MGEyzdfV7P0b
b+ER1nISdLAxXgIbbF6/sxGTk6WwHnx5tcnkgFbJYhyPq2JuDH3aGF89VA9hD2hGwY0RF3E1Pchk
H0R/3ex0j6nViozG3yTs4qf9KZxTEdB2tvHveR/avMxxiWr4E9uE1LL8RLXybhPWz75TnffZH24z
cJTITfR6VleloWIgvvBH5R+UMNUOXM8W0v5W2rb5d/va04HLNqvw4IEjTQiolVhJLnbUrX/EOKG4
eEQ7MJFibHUBmJd3MIxgNvjKCB01KcuREePtYVouArETnDcPF2jKPCiy65yhqbXDKJmqSoK/VIqh
xmcYRqoG8+yQeBqIM4mHo/NQKsp6FP89c3HiWJj5lmPHxmTFZN6xrD0Gj/u2/w3dO2Qr77KcZApV
UZSXZ3sqJ/yBy1U23jdKFgOUnqdtscOD9CvzwLMGNaA2pj87LrtFiPGho47sfoSpb/BqC7H3aFRp
K3gj8JCQjxpF2d22EjdOSrYpTWwN0Gd4rJe/asY2Ffw/X4Pm/9XBGdtvvDOPV+jq5CL+ln/HHEfc
vEvX5N0/Xh19uPtlxIDLje+qaaUgsoskYhIunaSwyLvvHoMwDQMC+4QtchVtGJV/Y57a33GOkm9g
tdnr9oKWKPNOmv54SGxW3FwpdyF6yaYBR2JFIeY8H0cf/YuQzC1D/f4OAaLzCMXmoLWG4+s7ITTK
QV3/9XZP3JaZYaRP/dTHhhAuYiCVanz1Pf2AXf8v24Ux1BNbfG4dqztGPDoxXPv2AKzfsZ+wawlt
0rKvIfwD4iq2j725PftKNdtgpLYB+ASJX3VqgG9wgK9tPhIwRSP3uzJGil6XnB0EcmDVUg9bpcD1
1X5bqtSEQEg5nvFzLI/PHE/SYNhHRTPKAO2Msn4gXGgZbothKTVTDH1aqrk20ZMIbtgTI5Ss29oK
wcyFxt50X02CoyeZqybUfydyOHN+EUTPJX8+Rn+GuPX7J//le6SpNBsVaunIhduiFKuIUP5lKZKX
wDLrYXoxKuF/eArguFsB3I6VrrzVEErpXSgFYpB46H21Smz07TJ+bBOuE4x9PU3W+ixUGRw+0hG7
I29a11M0TXuWCZkglYhHp7iKjBtBkvm0QrcJbqwmGuWdGRHSPzIJMnuB/0T3NEafDmeNdJdAhKuj
tCPpo7fyIB4kOA5x1EI5550/Pr063lHhFgZFgV5pzuPDYxEBxabRF6B7TMty2aEOFQqf3soC6Gt6
Bnen1V5hQkrLxZDFx5cI7Lw1iulLDTylifFM0R5wrrP4mJ0c/GXmAbYkthvDdeUnDtvHzl8g5cNM
oqfIMQLYh6LFTcCott2eLli9Jf/Tn9PYJeXkwNdLI+xGKhyHoYkeBOCjiPvZFRRmwKVEYIX9L79X
NkNuuvKruywd/Mw/3toIHyNVq/ZdGdsffqAPeEsJqdOJrxDM2B8PIVvEcJuZwLtJ3GfUXTYBHp4j
YjRrrj1Zl1kPzPHCJ/qnHGDMfXc/sQoJT72KmF/Aq2ZZGsJlfEu7Oy444uMwrV7xYS+kY5rc0Csy
f8qmqSqj2d+dooWLsME42XX/7g0zebnTKPb3ApXfkPXxv/v+jciSI75XMHIiNJwl9p0JWd47zi5o
t2CNUsURAttqCbac/d8M7SmlMkZKn/U4lyU18zALXgOMe9oHw8ATW0SqLAOGL9niBdXk9wWIgKJJ
4+22x8fBGZDA58BCiJIdvkWjBDfneDmSRAfP51BxoCrctYFxucMdL0RwupwmiVeGRTJeB0twbj3S
tyRpP+z82Wuky4pGB1wXkFCCJLh+5HcFrlaVrXFYs4WsrxgfuPwQFTtq1pYmpyOm8KdGFvBc7dO/
xvlja5TglIGVBCw5RwBiZBaw+gkz8eegVIr1VGUj67FltUWfaPS9Vdq+huPr9BjD5HBHfI8083zr
x58LHkKogKz0BVteVhelVVHGPoDlETxl98NyIcicoWLJYcBE2o/k94ziGQLHB0Q9qF3j8iGss25K
FxQiSe6i6xhdzcmOktZCtDrDvWhmHwlvYtilAMQKHSvqW/1yC+T25uyjZgON3ySgAbX6kTWil0UT
f2cEevB8tk6GJEo75of7KXPFvjrEr2UJGFwEScQuN+5PUjqG40IbAFdVkhf8ebJzjejhyx7ignUL
N0pMJy6IQQ+oZh+sH9hN4GBSmshRZ4BAO1sJ9PybRMmHBlPTIriIWBhsQ6VwhUALlRc16jDh0Q3t
xCk+EJdysvO6djusXZJjDkXXt6dgrORu9eqH9NFNipgHkaAMkp0+RQZQm74x7zGLaFXuAU0vZoTh
ht6iKhpkX/aYtshXcUM9p5vpYbpgRTbY5oiSsDw7upS8Wqa59whBU5ofk5+zSAVLu+Y3y5nLPJXx
C2fTyWGcB7PWDMN/zFQeSE2aSGIYm9lRYxmste5qO+eVwCc0dLf2xWi+i3CIBi9Sp36CjuqOZTP3
0g+qALXQbIMMNi0AyavBseXcYp6YjVBMfQsfnqZ/9BXjgHQDuyloufUn7RbfhrmmRiRWgyxW+sJw
eM1e5YT3QInItF0tYpGfiMximmNqAjgvab7PJ+VEMe+9ndvLmuaso+hHbtY4c2FgVD3CEZTTwJII
U0Vnb4uo7+cm+HiJOLmNUvQIvw7ajNSgTbAthi4sI6G+ryt9vi7almGD7QcuaowiSodQdV2Tty/U
g35i6MRacsSN9Xy58u1BTLhD4uoY+RRBVpLs258uithOR8qFWye7AbalSPCNG8HBXVHLJL6IZ7tS
c8INA81x81loiv66RSvMPrfvtndG6Flg39Mgl2dtHRxo0P1Nq2/DIZ3q+kq2ccFQplRLqrn1wZFG
YC+e8pGROuLwNJ/9KdQi/7YDZOrONU1Kcwr9L8YLdXC3rFeSE/c4HSWfTjQq37ewfkMgrio438lV
etv2/Iys7M0WSdu0TV7cxxXhq+msdr7/tmZoKImmq3E/YPiINutZWfNwWDwQ6t3PNzrTDbTHoG2d
sbgQ4cSHpj99gWlc+Yi6ayopldnueBu0IwDY/sP8K20Wmt+6gJPXA7dNOele955reK7XMNjNZXGq
lMUvfPovmc1tHc4bREkC7U0UiVAGJ4RMKgRlS1lwbXDSw9h5rbywM086l+oCt0RInuEgunsTAjNF
jdVbcSWfjDIflhBgsGCeMZ28EbwWnqz0GPQZ27flL2/EfX0OeCxZKNPwF8perDhJypgpL7rqKBhN
0JDZ93PdXhEKSHCwHqCq1DD4uQbEFu3KcLEfbS3LTn0rvEBbqsJpoRZGgIvl/EQWEc3H26zLmXaj
7mbf0k+helNc2HXuWdeg4i2gIBPCIOuxsAwMMEuA+AuBm10ZL/383f4+r9cRVNFCATUKgAZ1Vak4
lTEDV6oh/3lX7zWvigd7j1l+KNmU5JsZulj81oWVRD9w7yQxl843/ku+n9MSImJyVeYd1upuMqN+
1+mPBr9Soq3KWLwyzewH5E5DV3+3brQ9MS5Wgs/K47B4lbjnz2AcHX3DB4CSe30XBdrza72PdIPd
bkmldHcwymb/kuJvAWQ/J3cl6AtE+Iq2iYK7NxulWu3Ml2m/SVyx/W3LaY6WLbBmQ1St6ykSrPmu
PTnuZtDr49Bc3qVVi4fsajlJtP+Y2SJPEWB4GPE9t2FwDDUn+OYSVVdDigfJCsawmwL5ffQ68GCK
YPw/9ZxUklidwEuog2PtPFsA2sqkWV/5cvHmcGz6ciM3de9zCaYvQs65DT4dI4BUGQ05V/M6TDJ9
Ab6xsaxegE5lZM0M5wmVBzYMsRSQp4Sa6wEF6XYzBaxc8x1i8syCjdjbtdyRCAZNaVqNH+4sMS+a
QnN7OJMaq1rXpSmfNdQtEUebBeCc6yjeH8OWm9tK+PyQw+NYhkgN7uyZ4I5r5rOVhQxDU8ZAbnun
j5yHbe/HcXz6CeouK1tEDKHASAxEyNjE86PXEXUvWu5Nmfo+A8qfQmj9ge2v7kzZesJkM1NEHJhc
aSA5NwcV3dKEF74FnQ9VSfQjeBTkZvTUNI39v5e+lPnL7grPDWc2tnnHIqZps95uMinKks9av4IW
75lXZCicp6g8XOOgrokOYKjka5yr+xtSc4q1Icg8iG8/Rwy4nN1Yb1UZoZCwHh6veb6B6HMz5Rie
6BKZgr/+zK1svoJvMtg/5FPmTWf5bQByvIfUyFmxj/tTF1FhDaJzrzBkl4GyI5DtOewjfP647dXn
64Mu1ilH9m7whjv+txn3+AHkqS6rOdZ5MTHENUkcPHv8SplKBJ3mCp+DIxsLZCGovcY1KMeb5O42
byIb6vwj5LBaJd0p0DE8xEgvzJbASnstaSvT5OK3IyeOuA6fYGJtgcW4q6L26UpXr1D5W6NGH2XD
yXJ+ikJcFRotJBA4lCaR0amEGr7RBX4I3wHjf86nHUL00X+NB5+7A2s09e/lxeMhsEDJjnMuOXac
7gW6O+yWsVpEN6fk8HJDmmaxXRy7NNb907/nsOmNQa9QgD5ogC1Zi3Tf1f8dujx82p8+nIzoBWHo
nMFIF+w29beJRyvZeYikHsg6zlnpWV6BBixFicKQHdzOaLwrypAFqdRUzseGzwhZAOyg5hwLgLo4
ci90IYFhjys1/ulHu0oSw6/+QXf0i9YW9UFl8gO0mIsqB8xcLC9jpV9Dt7TdZsft3EAEbJJyzCgt
Fa0q8RKa1PaCmN0uu2LRUtlDjkw98XERhrAB0iKOZD5zhu4rPG1uBHSMQtqfvdvSSm9oCx69GTnh
QsrlBeiIV6h++afXSUidQa+UC+4i3mbXnrc96BaF6XOoy6cw0CiRBWR9z7mFZOUDVlfi4I5Fnn9W
Oc6KFfKQDfDIAV3/cDTvWOL16kPg8ibtF57vTg0weOdjlp+RqjYI/Jqu1rFStkmQfU6/PGHhU7iB
ETy1PABwwJYhseCU1U2zKgCaWQaXJhImSIO9sioqp2/tvcZP5MJAQ08TE3aH9+BdYi18aZHMCtTz
8uZkqg4E4C0JUQBVA8SYBTzmyXDa/EmFSHFJIglpLkR1c7XYkYtCGeZNqWdZ5b1tw4xIuU3ldSXf
Ll61lm71vQqkV7ZOVieNavwse5/MKXcxzLSXtMRLkkVwkJfZKJ5EADUNZ5SZzh6XzIsYAX9CmLXK
r2em6wUI866k8MMSgMLtsKtXXyloS2gYRGHRJvqkfI7SBEv0LBjlMv/2Q71CBpYZqj7JiXBJ78os
3PPZpuOkqsXTw5qukn6NaPo05TQJ9s1aLvsCfrg2WQD1EHRCuP6yiRX9w+ivNRYxVByERSYBn/Bu
/qHK1npHo1Q9RYMaI5N4Iuk9w8f7bU+TTTEYdEtMFlO4mAKWsDOgVyZBLKubSl3+Kn2bDmk1u/mb
f2C/pyCbujrLSIAkFA2LRjwJJbRGAxM6JeZfEblyJNes6wE20Ar+hCs9yZ9I1k/BMk46FyzL4EwB
fqi/KcU5er+nFobpKlCSBuoi7Ra5A/FA81TqhdLDwBobQJYAZR3+gnfaxphgSPpy/0ijszcS0+Tv
6RFy3uYMN6BYgmS323BWO0w4/fPfg7InfeNX8Zo5jmRgcnPcNq6seGIkFy+UNrB/PoG9PNF8rZhk
r6B5zu8vQIR9oVH4GCgORNFd85T3AGi2OmsyFbGY4W4/U8S6Zmp0vCC1zBOvZ2uAiuP5duzDLpRr
FPIjeCELKma3VyrQJwhykZopfLEzM4TywPNZrym3O2RzUjDWdglED52npb/Gd6Zl1N2yIhsseMYp
9KKutsquUoerFs/V2dmc8mLj1I9sMXgEDPW9kfqdz8YZcZvE6bhzmsJxZnwol2WVDYyf20mMlB/2
AJQeFCDtfGhDzh00k1YADkXb7YvP652WnumbOSvNQaeVQgutpli63eDebn6hEfUtbDwaYQLzC5Hg
Ys6/VaEGMsKrennHz5dpg+dRmg/l5LCEykSVKvzHChg22N5GVqvKhnO++xmXOJZTPyf+02XfuNcJ
EDT0TGm6DZ2qjGauEhHPn87i8LF8rwglboI4SkVJaFi2n1pUMu1OgHSsGcTWhM/IhGlVNFs1NN/F
BwPMX8W7oIXVbvqxvMFiFwkXiRjRwqU4Er3JPLXCPh7c89/qpZG2ZcSg+io/MAdqc6BJgVVHVYop
A+ZjAyaZEiU7BFC/55uTgHlBd3bYoO4Zk8Y9ouT/+v7eNCInTkfF07gobU4aJFAT/6uXPc0qpvVg
E1lObXQCqej1HjXsoG5efZgAJasstJvGiCt3KPVFpHoND/+b8aEPSmSha1qXcUZQc0yZiSTL3Ae8
NSpIviBh9tH5lyslYRK2Y20gQmROKDfv6WFEe2/DkpVFxcBBYe1Ql21UDP6e2Pz5nGBIeXYCGr5d
vZUnVUTvAUp/rvSmK9M07U0MN2mN7ZNIq4QdgBnSiLTLWsTj06BzJaARq2hfjBh9pDhYYq3XmLRT
85th+5h5kisWSJeku/IRjA7OQbQoucNJX0bdeTSFqQWkRYru5QXr6zHeLi38t3cwzeaeBLqCzh9l
clOoSTYPCMsVLqPTPaf5yHV5TR1LUyoFigdcUPnqn7uz4yvhIMnTo27N+SpQBSEITrzcNWOYQY6y
bvWXB5PTEBXQJhIDK4SvohbBpEFDzNrkB4PxGRFPzoMdfsv9IPxwAs9Ct682kAewJMwlAXCskCRz
O+rBxHArwov5KRFFGLfzzs5Actu/bNH6pHgXf8wAxMhm1PUss3wMoazND3zfM8VkX48GQQ0zIFYJ
nzBskbFen1yVC+8EueCRBesV4MqYy3Uo4z/9G8WsGANyv73FMmL/Qo+//HdkgSiDtc7knMY1373s
+7SKKkmvgKFaMFC9LrLONb16/0Oy9S09RpcxT35qVXHTUP5Tgqj9/Co2uuZO/q+CqbvyCBmJUNXO
hZnkPHD+zm6fr88fGDFgrtjAlzia6UAOhKIZD4B9p2Cc8Q2yEi/fTjpXCY8NuPP40MRCvOXJaW23
N7ADcdpK7cgb2rV/1VbUvd7Xx88U1UztBAYQOzmsrUHvmr5ska6uSTzaO7amNojG0jj3aZnmakGx
VYt/QwVqr9HQKuIs17jN4HzcNF8KZ/8onHvDTGxiszVnBNi1pATh6aXrZ/0OvNTEtX33uzJX/qR7
YJesk7p0arBY721GI1XuKdEz2OqiAmUlrACS2Ul4y7K0RQAzF0xVgtnHKtcsygzGScmxr0F9gr+n
MXzG6dKVSygJ0HGW0FEycdmGcFbYnloXiOPHGgkWTnRqtD2SV5wwio7L3BmkZRPUnwJ1j37xxDsI
VHizOggBFBSXRXDUiXU/z2QUqBouDl5Ma51UhMExkYTVrgbw6DNyCG/Z0dcaXcSsppl0ABRzFYH+
+LP5b6z5QiFwWfqRPuQkMHA9LU56mO/amiQmo7QXtgGX2VUhjuEDC9Xk8Tp0atsbH5LL9Nt5sylY
YwlKB+LT9xtw8h3QQVbH/It6Hqk2f1+9poOnlXLtYiNuIzSgiV94Ob+si5zc+wxrGOxiKN1RJC3y
LfW3Akm+0kqiUypMqy3Q3DcfC4zs+tnOpHZ7W6XNkTH3MGy1DYGmLwM3V8BKrCa0WIEGzWqGql0G
BcANjG4bT8IXFxjpF1Z6wquAXZ0adGCdxoNBM3YPZFTtPRq6g+BDOBcsB8nD/bDNjTTVfJB5Rt0k
Gk8cHOJbwrwfnhSjgqhXR09+fGJHComaNarfz6GFn1Fy6ciCop1jKcx4f2m/3/jfbmm11sxE4p/O
zRD6+euyD94ltNolfD/U/4xfTNfm9nDYQdxqHn7lHtqkP7y0rEu3WZ3dYfQKAAigzi55G2TT21/r
v/88+HAhRF4lfV41SK8JvPLU00NCLSJ8AtTHwp12TWeyZuUmkArOKejJfdjHa3ZNnji89mfLYKbd
Vn9XwESfS2U7M4Xr1JrRKisg78WXPJT30KLj//uLTMIV4x/tLsroRUkdG/iE9M+P9QCEzqgTrWba
Mrt9OUVpUm7Tvg92BVwDRa8s6xiiw60vBZmIYNYeHlzht6pWx8DMGatyfbG66AjjqL3kJovrLc+U
XxZp3d4mKaN474lwI9Fsr/3ThMPepUYfv29UPR21O5S5he9Yw8OVyvwlmgyZzeKem3NRRz69aEJi
zZJuy9UGFV3UjhIYjV29z1A83v8w+1SDEuY2pWE6AHyWQ+/Bke6g26+IR8Lq3TP9g4d+g36wMWjl
Rk58NbODBqJOQrCin2ApZa4fmE1FavP8St2h2gfw7kqOBerF6tHb27k9hK1TCHDXE/le0EclX8/J
+4kNFYjBu1yrL5tuZXSYIABmdYNpv2IaoZne7wgOgVbqhOfVX/R/4oDpKtqeOY2rj+xmrJvU8Es/
c55wbjme+ZGneB7dbaq+jjzwf/w06LYtEDUheJ8m9ZBWYwx6mVO1KSSX7wU3g5LRUOXcX4D8vm6Y
SfizMIEb64JYq8f7XJYKXPCGMWKjjtDUtifSynLlmURTcyhC0k5AsKqf7twf8/vXrhnw2wFuFKvw
Nt5F7Wmfp2eO+IDJcfkJuwrK3+cz1hQ9zDVZViBBd36KrgBB6a+vMhgNdVgD0efo5SmYx07irOAD
sd6rhaQcGyVTBc22SKZm7UiuArL3M8IBK2+BdrYlfk9e2iQlMFpav+QWiRanjy6eD2Jxir2Ryxx/
tG+ED95Vt4wP4H284waD4Mh2MaMFs/u8TvJC1SUZHa0reRP1bCDfFutx2PmR5++BqpoyGnjhD7lk
CAq2hwdgsX37+m8Mm2g7H+jzPzLbZn4OQAgedekB49zygK/EWJmg9i11Z1teeM4SlWLz23PxPMiB
k9UXdhJrJo8HloEHdi5xWueesmxWM9MSjwgzb+Z0iYInyFzmdMg26MPnZSIfJt6nHoVWjMFmOs21
k4kwlp0c/wegEuZV4dQzi/6QszbDlMxa1fu+wUaLvd1GPmSdVIZxa5U0RJo1PhbzjGtZcFSQ7c2n
pNhOz/4Bl402xiUENirgREizH2j6NTWhGviSaKhnl9a+3q0AOLXQZ2on/6+E1uktU9UdGXIqmfVf
QbywT1NWt7g0MT9+EeSZDSI5ntnmH8QwI0GrDCLquO8hKoo3+yBPE1k9GQpFb2P5iyJeWJ9ObDFr
FN9SS0TDgmptoAELN+bSi/AmDDxgSItnkKsow3AeMx1ErGVshJInTwz0iriLrQL3XZiSnPoCKHpP
g9PE869FPUE2XE/lsYxhM0Q1zQnG1ARYySywkw40HgVzHzzCgWMkF+AfJ1qTXgizmG98w8rrBZgS
rSeJB2kSw42iCLEH4AjdO8wtQ2CZLSV+5UecjnWvI4jJNOCqj1uSYDr7buoe+qNTx+/5jnz95/VW
rcKd6ZVweCJAn2iEIa2RHbzv3fOFgc430Rn53T0XK7SszJzCXhKnTW5EqKXrko8EhOBIz68xMcwq
35T5s0vpfjY2CfvIY2JyjRheumzMXGtnMbqqlMcePKcvM1LvxEZrb2oMUYI97hiLdrmV9Sm9+0y6
oi0+hE6fU8yTbxLQNSEPL3/ZhARVD+DIqL84aMXNbapW79PYZVdUMlcRF3s4iP/NdWShSDsuZfEd
utPovpJ2vQ77l1SNIHGSLw2lwsHPxJexJylaiWC2itYVuTSFkSbQ3HdhA6kvRt9iVyTOlsH3Kxqy
++Xo5qCsp9MBqnQpe1XsE4ol7maOG0/lbdiPeCD1D5EMXAwJlZT6CXVQrLf28930W3XaKJICvSot
cM3xGqoubz4H/8v8cxSqHaBuIL4WCa56jMifBY03oGje6CDoZIqU6g78MGVyIrnuDB6i6LPUhORE
ml7v+hq/b4R6334Ts5k0y1HTdtqpPHGUeTxIuPKamW8EyHNYZZQKwl6qlVG3eRdS+iajmTEfQoyg
SMLl8h4oUbDk9NlBvOY91MsCJK3vEQ+7N+qQPES1dN8qrP2m6Amly/PfxS/YXkXoArtC8Rub2acc
K5Hwq6zj9yqkj8/6o9A4MiUsM4oQhZg6vS40+1FDRk3igbhBLuIMna9VyLYtXenUHdccy0r4Ee/9
DxUhVzODPDD/cZnmHgzkuSwOs0v5+o0sW5cSCeu+sBd49oRjTyldi3WfioWTfpnpfMW6Hkb7/zvf
0IJhG4ktg6K0+cqAYk6u8RiXsXrG1ELZCf78FWKbXl+Rr65bun8w3fyAdSJV7OECWEYVa18YFFvl
KZu9J/S/LK9HGUhc/lJzHSOpmhctb65pVKyA1SEcUXkz859pGAaioHf671b1YI7XYVxL85jvuPzO
M0VXehm/7N55I/IbDlHPa6x51hFmHZ6TiRoQ7Us/idlYuTpEnusEHJuV6ehR4C+YFL1SfdP5qe2v
mPqNLmc/rWsECETUVCseOnQpivASJm1gYDHb/QQUUhHKOkS9eqzUY5fK/m5+JFYf+mmUUiKpwuyT
jyWrcydy7vIEc0/UHCOJKJ80BFFUUzkoCa/3YxH4tXCAdqqfDiDM5SJ6F5gMYpuDd0UEalr+UKIv
Ryn9LWZYgCp4orv3axAmwQGcQjQ1NAwqoH1YWCRrun4d1Js7me+Wk5VnxZvqC7KEfjNRDCJgxQkp
VYwnK1gDsU6h+jtatogD9CUhQZwC9rHnJpi2Z/5Y3vXaxnkUrUqnLpP5nVG4uwOWMkw/0bgkgcvy
ewQKx1rCJC60Amnh9avY1Fqd78eLAxoHOI2kq27MG4hw+ohOFCP2bpe53mul5klx3a7zvu1Rszc9
ZIyVszDD3IitcwYeWEOy5fhRBjJ92zDd7H0c27Q2vhH+KhiBceHffVYcTA1mHp16aFBMXWsJF49a
6prnKxsk7cUwmzHYv7yJxW1O49PqK4A4GrEYFafKZRzos5pOe3jFHUj0xZ7NKjPFZ7TtycPa+3JI
R2oOS52Cbsry7RHj1Yw3eXnYmnRvEud1gCeih2rYmyp0buWuTf8AIYKOKY8omtzvHh0XkGx2eZxk
pSbS4ExVZ5ZdRgMcyNqcTPowOMsF0/srPWbWLbWElWpgGWMXfbtFOnUgEhGst5NNa22BuP4mMs3C
jWlb+Jb11lED/nvGBr+zZZCqmXTegyXkn8g084omrY06NT49FIrYIRkJZHhIzVAtGTxoPs74Ah/L
B4/BbFOaWvEF//56g5kGyEgAMWN35aXQlFFEzUObW3lwpNxbyrIDFmwOUPrgmZgNuSoxCUSfrrVQ
Hd0zjW9bUfTxx6O/a2KTVawIuAAdrAfrqeDGCmCNHQmkc2KVoD05TL2YhJnMCPhHzTxrzkJPRaB7
n8pnqAluLyxZRFm2+/maRMAex1UGC6WQIZ8+oCtUm/Ebbn1pzNR70+XO5Lpy6Z6OlCWjyR135bAG
yh+pa50Y74vgeC8/wr6YzqgbUdN6hTGsytPqyZxE+D3mQNJSZPbyai3vRWCTYz15fFp27r9BmOz4
INdZrzQRccwoKIXfvKbmcOp9gAzhjPP+hHybhYrpaHe5L6cc4p2Rv/h9pyaoqfULDneE8QCObMzz
6SpQFDhYBckLh0JKUDXCDG6s8SAGMNMj2Vi75E+vecCGfPgETNMo+wEXijm4r2xoBIhICty/F5O7
KWnUmIXevr2tyK1TEPfteGofqKeYePx1Fr2uOfN5wscEvINwnz52PVYC+pm0sKAsk3584FEKca4n
QXlYPCEXZFrs5Ho+BYWzXIh+dWUiJIQcS2reDl40CP7DB6gzXXmNEZFmEUjuhYKTr921B4RE8Wnp
qO9a9BOzc6LjkVi/dZYzq0R+isuekcKGygqBA+v3gATxQh9nknHRdWRu4o+GsL+EINsd9/zv0Dxa
wfGz5rGSqXYvm7bSk87YiL4c/GbMXOiG0Of+9TG5H0hrNr1iKA8yLRwIJp4u2Xl6cEOb0SistF/j
LMkMzdkUwU9oRjQZXA+f6Y2Dfkth0v4nCKjFEaEl1QHOH+f21bFR8AQaPq3UCx4CIOuGhwzVlWML
h2yaIdQOgs2EI8h1T6F6uFeIhoJTDPtKKPvUHFij8/7Ik9QF2CpnYoyqKjCXBkEgyYiM/aIcQL31
Sfs/iwIv43jhBcZdD/jmx8LNw/GdU7MnSL0OM3TvDeCD5ed7WAVznKjlppdmnG8ugrPScPBx58Zj
BHdL9v4pFOM2uy4vdOqpLwUHxmEprtwCCGYnNTpeMTyQf8aN3T/LdTFz8SihDHQbwQZqonYIs/Bs
2rOfG/Zga3oOTJ4OzsBTn+ZfHqyyBlOHZc5mLUHVloISG+0+zDySdwJQAQa7vaEddG4xomnwTOX9
e2rLCqGiu3QbH8x1oS6I29y1kxWQFJTDefm79DEAzHOSxjPoTfJP1dOkT1hLkSUQk4c5NZdXUJmi
bMrqRu1JPpazXCL0dKCKutz82yQAAFivFjzwuDzY+ks7zlwC+xF3MDt7RkPXvLicxmRf8tq9ylpB
NLdiCe71eECz7wDZVA6bl1bAPuKAbp5YnTqPEo9MbVewkJOH1kTAjCJBw5XFCsX+Klhm7a8oHyhY
F0KYNW6+kNrWa6UeX2BFHyE0LWUd7J5uvhIwkXokxJBpx6Xvm9+7OPrefmAzuVlGq3o2XNB8MmQN
cEqd7pnl79Z8QY3bbGIqv2BVzLhVmVotRmbRygaeynS4lEH03eDcJR9QnY+UNS49QAfQb6MbzFf5
MxgEtTyLyKBlMA354CwhrzJW6v2iVta4mCZLm3YT9LfQPEieRc3FaEROJutTYSbrqfRt/xmguSH5
sU+nzsN6ezC0+g+EKA171RG6w+kVst1wSUBzEa8eh4IwRmZwPnzsD4ce6ePdRbYML3+NLzhDmaUy
F2MP1tVaKTpHs7v9RyAIQnH25UunUlMWSZ4CZYciDEOeSaQDucVqttwFr36tV0+67cKOztEoSNTh
VMGeJYYOAIHnbi5nHUQBM2W6PgYM5g/NOuivlXIPNKDxMmP534c6yCPvq5f9eOnTL/+2MIop7PMR
1fzj6SzltfDIBsgNmtHWSZP8DaDxnvyUfvfafx+pFbyfHyTq1h5sqwimXJ8fGL47bLj/UZFHN6K6
sb7eAy10oV402RGW9sFbty0XR1HTMeKRSjbaISvhyAmnoA7Nw6/DTvEPol9Y8y89zkA61wMbmPmU
eWgAT7Yh2BblHIU+ygJuk+3EBiyNvhAhkSB/ZtDe27q6s99oGtVya8j4fe03yn4vG74ytGriKGDZ
fFmaYQZDIyWiq4itzdnVp1lfy6S8gTz8I/yKH5RxpITnAl77LWBk0jAkWUcBr5J1st5ClMZ4oBRY
xB/WFdXMs4M2MCdnU+Z7Q9ee8dXv64USk6NoN9O+ip8rWHmhXWCkKDUlD8KcO7JVoWetWcEAVtO9
7pdvZHR2+BygFf8HaNa5XrzdXrAgZ6GEYqe3t0pODhnuskGpvew25eufashdTgX4CSqTG83jUcDL
RF9DDUulKt3Ho0f7PxeGffPROTDOsQGnuleQju5+XYm5L4Hg5iximXJ2DbIEVTZGtcW5DCn1tHs8
6owOMpP5Htaa/hZYLAjkKtSW3zoj29CmJGxs57bseqjP6xLvKCd2MpC1LnuuCO3NkfJIHojNbcRD
qn9cEHdiwALPlR2SAbAUpe9OIIv6qFAOlsVop8SeMotjRPqP9UrOtIWqVFy2D68SQFDBG3/elkrM
yDrKERhOhl8nFmWRgcR0JNctmdTC+y0YjItWeZ63RMtwRHrNHs5H0ArZEHQWowSwYdH9KcNBmSof
b/b63YcidXGQn/V7lXQBOFLr9yIP+8XnfoImMQZmuCNDg/i3lWh5qw4H5iSGVk6Nu4uzb5OThiz1
VcNwDCBlt2LkGQkuSNKbhLl4okj2UztQ8yBDlrZ23dhDeWgh73HJXVlkNFRfgky7EMRm9ERHrbdo
W2j95Z4LpNgxrbJUT1VNQswHqFUGjZIRKIdbX8igNXCIBsIF6tBeMsYOjBNSNuo8RH30WhsVKDHI
0c/VMs7hS1dlMh6R6rbtlfVcZD5P8PAnK8LhWfICekXtc/3JqYomWn2eaMqVKQvWTrlCwRcfMlQK
APub7SFXJjFjI+FcsWNG4y/tDVAzrC4woo1a8nWaozWkQ4/csI9gHtUZFZaQ4Dgo3U7TBm0wil1n
5F05u2oi9rd0FfU+zBQIfFl93iqXKauOlZk0h5inN34YF/R8QiceSFQZiLwhM6l5VmvSZ4munLLc
nT1gdnVK1/e2T6qjmHOOxG6bwNmTdkmp3w2hkhjwxtG01k/fmUW8e7CNsW3T9UJo4BGB9uPrF3j4
asCTxtQL67NIUqxm9NoJPfdaS2xLP/i4JHmf+rB/q9DH/roSOgQb7RGguh4RNRxa+Zdr4ZCclj+3
FLgNF3IrgMO+VXMGLow9Oczn+9FwRsoERE13zZwfW0yRgrTkS4F73Ti2RhXcaWSVm2HN8h2nuVqm
L4wOG5QLtsDz+8DF6LaUUYH3SyCZjFwAOjpaiB6SaIQout4A0CzC0OGAScP43VS4a28wFq7Uiyff
kKq7CRK6O9y4tTGYDoP+8DWVvmSH/E+ktYyjm1U4kCDX/cKSshRn+ox54gpZ5pCmIRuOo8Un+pb0
vNvx0aCsGNM74v9H9wI0Az3NlDu0zw5EMyORfYQD0OkYFRdZJIrm1Dw83GCLWNiEDf9HwbMs0B1c
aXieP6Ma7JKo46BhNZ2vauneEp9MY+Zaym3wGfLoAYIDFK1sVGvHD+dMeXIx4qUAf/OFfo/S33na
kb/497oGYsE39KzvkJvtLv3N4QSTTqmQTxBa+RxyxkJB7Ak2INk2gCWCW27eXJgiT38ocMERIA5z
C/p2eYpLENoRqBBDakxK7FuAv7nY3dj5yUzQohpEo5Ysrp9g3xhjsj8LIYGPRWWJX4RmfJSzcZ94
bnTEEMwbdXQjV0iewsR96KUqlrVIMB5QMlGj40Afj7udW9FR4FU5LIdMgY2/8Au3y8ya7rUOwHcv
SJDNYB7s0tcf51blEDXiOjWT73loZAJ4TS3fEuUSwl69qIHIvHBZGlJrujTOb8fDxgbHeZPYraTs
jWThbYZr5kB8OgknldQBh3kyegUANz4lTGCpQvqCbcXHZaiU429PtgJdfZTBG1UdydN2xurdqpaJ
acu0B92Dd5O91wSy6ZEoDhAYLnioWn/w1xXBaVU77BzEUgL+wYqO4EZ2Dr2uVMHWiie3hiB7Bgbs
wEmzVR7XZbtL1GwlVRb0Ln1nDJJW41E+OwUSSIdIHfEQMfRl+G1pJdpxC3ow3jTAj8O6Cf1nQ18O
GK0wpOQtXvWyMQ+kFgIT3t9IJK+cP2rFF84qab2c3TwVGlGnj5HBHwcpPEIZj0j9rs54xFhFLH3r
VXEiSNgIUmwQBxFdw1Npyf49PX+4l6o8ezdvHUgl+DocdxebM5muQuPq8gUbJr+HqlbTgSLwmLwO
Wn1uID/5s3nNBg+qXbZuLVmajrSii0N9msc9BnvbEwzyqZUlfJdrnPTsk884DIAr9Y1+cO7R3HW3
Lv7pqKFl/2l7ZP0QUCy3eU/XXqoONqFk7RB1WzE3KzZE0W/42DFL+xPxqlD+tcEfedBUjtPLm1gz
OM3NMMepDO4CUIFTe3uUIb/F9WOz/kvCYhtn6H6Ov2qib/Qk8ChCRRQW3ODa8nmHYFj8jPdk90B4
90YgZUMSMzcHqtgTgi7UXyWITZWOjdjbdQLKQrb1YfNnG/Y5d6BNcfrm2Fb/dr5JMQNdiA7DUxf/
irjwqLtY2YSQO70NmNgQBGHrofQEioE/qCwNNX0Fmv9JwUcZmpQYpmpXJEe6BB/T0Ol/ECI+bh5o
qw5VsXdZ1jWH7bpvzj+BX4jU+CazSbz+VZrQH1aL2Ftd7dJiWEWNV0f8ueSR6VMpDeGj1DJv+oJm
Y5evwVBy9d6p2i8iIl1zprAa/aF9UxNK/nxWePXRlQyLm9BMETIFJxStUzswlyZUuPf0wvtUuTBE
LD3wqbac8YLpuhLPQ0OKWmZnsUE2dSkycXDAvfUTSwMuoLW55YmpPwSenTPzeV66J8JU3vBIqkh+
2K80cnbcYOE46MHzLXcAj0emLDn0UfVdh1PCISh7exlQZAQ+SLM+He9ihSwatJzWiO4MdJ6Du1GS
APKGzsCHxW1LE7U9FvFHpoua72Lj1EOk6H4N6xGZJ9D+fEKZaXgCfI4aD+O+PWfFXB7Uo6AK2VVT
zcHF3wXwl2b+I1HIH1+yjoZNyVTWekj8kkZL3TIBVq3uuHyGXuNS1dCb+1epEz1nETgD01OqEPnK
LcM5V9DwS1Dv/3VMeZQIkjz178iuVUztcilizaoE0Vre4cUkgdEYcPoWVRRIQnNiv/6gTYgxUbgw
pSi5im6Nx/QGKy0g6evx+LYUBEpDkMPKqv73lNb2SRc1+bwjlZeB3Mvu2zqs/2J8iRK25+7HXbKM
Mz0HFu0W9BHDlqI2uZtrJ2CYc0obixY+gVAhiWCfXOU/wKRZlLbodgEl12anWVy3a/mhNj8gz8rd
PBvtwttjT6HHO01PuUal3doRSHZersnJqvm1Fk2i0c/GImQqpdZNiNTEUb2XMLfERXMuKhSKCkUv
M6kJk5dcKYPPYACGMEpMDz8U/yREE4QuSYpnlh21UD3hH0qdksunrmFwIO2KvvNihsz1Xgt9hxNJ
lca5FxaC801VhSWYd8ASdfSjSgQuOHLU5bqT71nKGAZz2xd2KiQ//ZDEPu9BX/UhBlVzCiwKBz0q
7yLQ/8x6kxCe4ndv6HNQfDlwAZ57BbhkKJRZI+tlNzPvJe4rh+jkZoEkgFpPe0v+U4pqFk/XPdgn
LZWwr0bPFBsG5zabSpexr7ZruflyFUjEH7MtcZdoRVCZ6xYLJQVjphu41bB+KP570LXaXvglcflK
hlnqMY82izNI03Sejxyn5dwqfhXIuqdqwVaUTPYrF0CRd4/dDWVOkQeGY7QtyjpAMsTDe0kbqTWJ
xIsg7l4pDxrPGojFns8kwKSQWMJayTqUILnEmQr/tdU6Gh5hqa29YNecFCQAcNUldz/H+9Mvwejv
9nmsEGb50m8REniRPFtyQ3KlvuGgBcnx5C1Y77EkmxX2osll4HGOhdPyB8L/nBZlZlLjvVT1uS4N
9fqpMQt1CioHCgzGsWZ5SU8nMfQ2SC6DRVm6XlQVifjZQ8nzYK7LOYrmctZrMod9JFWxkQpygp8M
siceCBIauiq0IX8/QfmdVuTQ3niM778NW7iEZFrnK7Qty0kfowil7lejb/Kv+tbniFiLpDBmmPEb
QrhSKpKaGXr40f5e0LewT95Y6cIVDrxcNd2qU66kKfGcABM813DAijHv99GY+l4FZMXFZWEaM6b0
E2RXjX5ESxllFz9NN5lfFRW8wqKxrDIrh8cZm4iMo3NTCtt+FV8RivOrXBTgkBbf6fzBkvH3goXg
ldMgc/iEoUlwaxtqfrTVKH29MN5uLscg1IVXzFkjZ1G/Q8bTA0m6sarp3cfp/UoW5f7oi3R8sobq
rmEFUuqZSiUFEzHvjg7JDXttpbbkgBwqtN7SdYPLJVTRiOiu0rELmUwVbvC6Op86rsIOuY0xdnTf
q451KEUm+w1oS1D2stToJuee6wfnbtBtuDXs7EMef0e882oVUykn2pBKwhVWZXCtbPxxEGhj9QGN
DYiFILQu76Hy4ti4k33AoObqIdFZF9Vf4/abGfpiJZWRgEoeIl0K/BW1zxrN0sLaFzbAq4ULcszk
xXxyuCleTuFz9LKfjGux+WuJLfkeQG4GdYEWBkLNAEGEaLqA/Ff0SQXO5DsSL6UWfeLJy21d5MbQ
hHg8SG4yFCedtQNx6n+4rHt9Gw0LlurLqfeQYMi/p8s6O3LsN0smbZ2DKhAxY2QyPSNTjFNTs9se
+bq1NUfiwlmfXUje+s16HzUORO5863r0acFbMlhF9ENFgWadh8/UYeQ2aJaT8xmiVFBvPa8ugyY0
6Co1U1Q/gBXC/EKG2Tg/rC3OpsVMNPWGaMfeWg8+vND5D0DsAluGl5pqDWfAgrFNh3HKmz6jVWgj
IitRbrrFPJ7Nr7I4ox5OE+/lzEJUYbY9mXZM3cCgqroMiRLmK3YErzrU8MLbrqgHOc9MdYLTMvCL
nqohqE6xZzP+ZIUUTccY6A574asUqW/xGKYRxouJh5Y/zp+x1vDsPBN9hCtwulvlCZz4NRyW8Bay
o2LyX5uVJOSHBIItj5j9YoKrkkM31MtcgbYHnii60Rp1nO6cYUsELzlBTYbg7BNzzha24q5botez
YlNuFYsk/yTSnDZJIlSZeyUlK5jjqb3ZPF8wWe//OswHk1ok9LOvZk8tVjWxuhzeqAauoU3En2s7
7kCOkvaOhcyqFrOKHOzIt8Mveg034ltx0dxHzQJ6wibsTDSF2jcNLWBat5ucC4FcmVIPZINzSSnd
d09fSA5wqc+uDTPl3lIbAJMLrvIFRk1ZZGR6qlx63fAWyJUH/tDnctXFTwv1uO3mjBrOm1aw/yzX
HtAcRxl8awpj2oIEbYENNxiqVjAcMATqMfd5D4tk3UXLqT7cg1m4BW6Le3tGyXjh79IY4FXLw00w
ICJK93CDzhCzXtkM/dVIhPBDEGzP4Ahs4ZV+EFJRZi9LDVHMEZ42+ChyOzZf/qJBWwnli3cyXr12
meOV1XnzpT4ySHDpukZp5OUNcoFrbjymDxgfFoSFrONrSFPwT3deD2TwcMK5hFTz+0hAvh8vlW4G
ZAihBHcmNAyytHik3WjKkaevIVH1DVbSTA5tcIMS9JsOAoXi67h2TSFa5Rf2rxJq9/94VU1oQ7yT
sDUmpnCOoP+KAfQ8TA0eWzUcNxXfcqlE92JRSCmAKt5bVQHfnaCQ9oQNxsFFhmvtNVi9zNRwxm49
BSRaXtnymRfCAoMVQhehvSFYrGCvMPpOYBBH9xZTJyps/eb1b96nktDXuCeKB/4W6xAk+GBEA3Aq
MDlv1q7uvrjzRf7cQ9DfkzX/tP0ThJweKSKDqKs29j7b2HKpbcYjEuHUkN64otFXENhSMZaQOQ9u
JSG95D0VHsDTPM5m2qssy8r+pQ488eSJRVsSabyZlPOUVYpL/sjXF7/dNpngeuxtbAE6gxi47Ik3
H4/Ambwv3B6HbFGc9YILftjfXzRxyLxf5oSvIUcVxgBiE5KixShaf3TurY/0utuIl3IPxAXKtXZW
RZ1gt+WGBW3VRXZxDp10HMe6QE/3cfkavk8bCYtILaNLDDGpH9SoLlO+PFHBzEnNWFcHbTfirh1n
CbwMLsaaLHTnkPq82YZp95xBVyFjSU5ylFCfQVzNmcDzqlO6nDGgj3vkiM0DnhPtoO/5qSXzEUfM
RjlN7j++FqS2dvsjqW07GvtYdtnErDLxvWOUBM/UyuCa3yZFRgw1Uq2KIl2cT66Ek+2hOct4QIDI
xx8jwojuJpH2KlCxtVkR5Prw+PfyzM4ec4F+rCRsVDo5ZTsUg9yLoUzcE6BV0hTZ1NKwWKZKOh/g
HsVpxRHzz4vtJ7E+qtQ6QxfVD3Sth3QLgJDzaHBwbVYeDrQ8jiDUChWk0AeuYGoqVMoKd/cAmom0
vlE+h77l9lxOgpHz6n/vtH0Dki1Vhrm7TGikdY0f1R8cO/h1SCJ4Aw2wA29Sp727U6WrJE2pLvvY
hP7aZpyKBvwHz5DDrKzapX6x6RJQhUpPK0uljsEyC1VUKXf2Hj71B7XPe4kfzgu0HDxTKFnDU7Oa
kP3E6ajtDVlI1UopRieC42aw4gfyM+/Edx11dgETraVATRDetJrVeI25R6IRQiD+q1MaSH5ebbpt
Xkxlv0zrD6FGVqtlfFzI/mBCuQ5NqBH0a1laEqxndWBuPbwI2pYQuRcNMv2tect72e/nm512fXSi
mu622myGFw64UPLr8h5MDJ/x58dLVHSdaL2AN+MuhsAirUcxqYYsde4v5PXpjWVK4pYeXNPLsyTR
NYc0S/wJiBUnK1SxuoBZjsApaoWgZ8CiTgaez1XXT1WvJn2OqXHzBPbe52UyCC9t1qrcT1oxrtto
BEM76F5Jj2A9jCPK8sX7vu90wN5c0ptjpzlLytAKTX3WLYdeaBWXNAPhCkAYS7/YKB5YiNKudemH
GD0RPnkRF5XfCGBLsskUc3EPZ8jnBN5h+KdELEv0nraet4xI8f5RvuR63GM7plbkLNdwiGQ7fJsp
gUB1BHUOGHGMkbHbm3VS6DkyQPPj0x/ImRzB1w81gyaduW1dqahRB+NjwHSoEXc9eo/Gwu5Bt93c
+6+ijgNoFeXDeXqD4sAqCCCwCFKfI3eI0zQ6+mvhB2QyuG3CvBFSUnsxCC5vJ3fV6nNZ3PWT+a3b
HpIUFQ3hep8m/KHLtzwL0XcauqSjanFSsZDA+EDs0lfinxTuei6gp/sjc1mMYrKrGv+tqV8nJwi0
yHYoFaCiCUvXJq9f59F3UlGemRSEH8cvaHlmtzQ7dQnLo6ztSfH3eZfkMuKo1ENXY8Vd0TR4g7Q6
67MkDiQ0VkTO4vSqdVYGZIybIP3vHKVimbFW/Wde6aqj8wvddkKaggd/x6uq+brUeFrPy9qne90/
BRj+uHBtD/3DEWAXsu9/e1e9ClkyKNLU+mVLX9Knoix8N1vEdz0tLVl+djD9g7A9aO9sHK1rCp67
9dOXNpSXknXay21orsVGN97JL6aNEz8xmjK4qhyVfzsYyULj2K5VnQETPsaw9nWRqJau4zUzx8vz
tRazyDuzb0ZqCYbCFkK1HuOdjzlQopbb9/RL6m2S2t9dcmgLPr4ySIx2LnDX93Ed1NfURWuiZkfC
P1P8G4jfp9mDYEe2U6BSnUzGPcHNfTmIS+uCfang1WO9/wUot+QMZFqZF3klHbu31esdufsO9HVd
A3opF15H/Pe9EeBz6tfbGIDGmEf/3xwra+R0thGsj0W0/gzhyxsbqEFG2p3AWFPgBxeAwuKZoz/y
KOsd12v1j8Spdi06hMOs/BC1P9C8bGbSrxYzv58HLipNw8rT73dEZZ+oeUElC4LDGbezGf807UJ5
leW100p1e201PW1HjO7akH13yGWdBT41/LCgudyzrG1LGCUDPPzew4eajBQZv1uPB5h4K0ygn5WD
/KiX80s7Vvvd7RHgIXUaZbJ4xnMIywNd378zNkRFbyUZg/186TmgW4knZy+JtEr0O0eGmtRqVmS+
H3Ba4smf+baIHISrsnLTVE+74UW3GpdkTibkZ3pK3thx8l+b/azcHvgTdg6hh1xCMUC2Vdrfjllv
BpeuuP12rk3nAscGnZCLXeVNUUX6LkgDeS92vDA6P4yQHh9Y3yV/8EmnWRzniZknpfGHn9+c4zW9
w0jZDpzSsbzGdjaniR0U4E6bSxbQfR2VhPpuJ0w5ycU5tk76pqSgCQ9GcMztsfdV6z3edChIOnqx
Ck20c/sg5EtWTfoR4Ib3udtEiOG+FByNQi/0Sa2hGUDzDH6efURi2d0pglC7r6al6VtCRB3ntSe4
b6f4rmIdwv1It5wcMbMW9Bt0RySGXj7n8h7oXKsfVONZIJTqU+hLpdUudLo9DBrxOlAXnli+RMXZ
y8cnhiz70AafQXCgiN6kcrPUsm5tO0lRlE7zsYGs1Xk01DbYF9/jROmG5jhy/VjVVTmB5klkbAsK
hvjME4g0J8F7NxEYSUPolr76JABrNEBSUz56dH1RZ/U5lXuWT7rjsf9nbq1p8hekJf+P3f6ToSwz
D0lL10nPYUkKMk+1+y8hv2nSqFC5jAK1IuPiIdH1vfV/Dp4iPkkjio9Ite/nYMsGNIDPvPGJaYJf
lYDjly1j5MDzGJmlWBfpw9jqvtIj2HTaxnnr/d3V+MlG/sGeY33f3RriKk0V+HYRCzEbifQBce0h
4n4vGxGlNWqYVbzT/QTTrGpFcWuO/IBnyJyHd9J0ouMiEny9FLH66fTEjS5voSiWwYiJ6IqfgM9n
4q+pHIqB3Kfn7uuQQyd9e0eSuFpgHslDEMVY3yXOdAaXLrJHUg1IZM1sP29lIi0l8m8LoVb+nxDx
feTxhx5Ko2kNJI8RU2HAbNhevkrj+jWEZCwlpLtZHPX0yuBDnft8yHN9tEpChzUH8sj9LDn7Skyy
osf3uI3JFS2l3fachDTQxWYvCOswkvSAwH6RsTDiswzdYZfdJYLCNHIM9Eg7rywXrWu66gSKSLeL
3QqIHg7aMaBRLB+yTYAKpN5Nm7Cp9i1eXt0AcV1ikgAkkHMh2BjbTMxDugd4sgkIoNJdDdaqMfPz
+HGDoYnxbtCZjXQ9fHHsjgCFdbW7lnhcNglleUFWf3fPnc/nseTQeeVLvFFdMA7s4nMXmXtL4on3
OZgIiW20OVWa33P4fkv4GH8CyLF7YZdPluVEf3HcNg8KzVLF6I9/o1FB/xAkXH/keWBsJPtkgI6H
ikA/ztPFbarqDcmowSx5/gzMEkx9zDRdTnMg5uiBfRyKbtX7m6LPwqrE3s0JvCN4YSgNuZEh+tdC
DqEPd9rIG3aisaKc9yjbJc5r4BIPdMndRYrF9d/qCOf3Pi917b8n2OLDKJUXflcPRuKXYSvfX6/V
ifmTFcsw+YVL46yVocJxHAwhPHF3w8rKnYmgU+CwraSwIRVDArYcff7q23RI+UcRYb1VHiGTjOAX
q+dTyhxXfvGNfNzUFNbDTaD6exkOm1g0NakfZg9BR6BM62Wva/LPM5n/VaQunrEtct0J+lUb9IWJ
MSHjm9l8o3FOOLoK+Niolq+XgC2/NWCVCWqBOHjmqxXxZHZ7hBUeLU1DDDk8u23oW40yPef+5CME
o/kv2njxpp/pNBXajO0PARNV0gQCC0pTrrei+zprYCIlrU0DR5CtJEyXJ0EDZGme1KsQrnUUmEd8
gpM/LSaBFSJGtRDa2tVaOfRh7CdUSk/pWI+3NWiGVskXWXOAeBryEyl6PO+LzrGxGE0Jo/dNenSW
EI0qdPQNv/XQ4vIhnk8Hk1tpNb1pEcHexrZkxZp3wAwARW18JRJgg9DDO80N+Ep1b6JXrtldWAXh
QgMW35WOE+XyFRplO4Z1sfpCrkFqC91y6PQWHnczJxuS7gjmADj4bmiELDqMZIH68z43kMAgc+XK
ZLe6auRyH91AIsbsr4k9PQs3NJtGeOy99QyJi+4jFiSOELsXLtouDgM3UX13T84QeNU9pvhSZzG7
8kOFPBReUUj9EWqkAf+x+/yjTa5CW2kNlhukSJE4kBttIk4PMqTXjYeAC0idxYEC6pJcbu/ZPB2s
0aAalOMloWiDungc0BSfsjroWYuDQOzhDuZ2U1lTFiSbAJHFqwe/ihWdXhFjvOZeGv09h13eRHXD
hm815feQLm76QE/yOCPQU7Z2hlUJk/p1ibaz31OdAjcbIE+wFpFKTs0rJfWkG/rIG3l3JLJlTJDn
Cq37sIWnRQn8qtjiN9M+nAuSWEkqA/g/ApPt/Bfh0t6NviA61YaRzKg61KhDf13rsKLnJwzcVYZb
gRZ2WeSX8K4JQjM6E6NGklzqJ8lU8YxblcfZIARLSRlYjVUFOY6SOa1d2hOdRrbkIu3Z+fVLmlFq
QZq5iP8hOC08RxIqdTsVwiOXFTSaxkAJdsBZP8wvQLFi/kxAdOl2j5XhyvFgDD9f/QmYNeH+EPwW
+ubwQBV1Wxzp+woNr+ZU8I4zvM3JtV+FLs5eotLImNVZmfqh5CUMHja/VNrtZWNVDRcod0zv6R1t
ustFoS+XWi2CmsBrscD+YCb3smF84iFiOFjnOR7vbQb3YJ4JmZZ0Ao/xkwnEW4Gqldw33t0Lcr55
0R7o3vrM+RT2Xy8EbBKDkhHAArdo7IslmHzFG66R24dCzRykPHhViBWtmdP96IuDVqcOZcJVyEkw
z9EaYDO2bxDkMCYori2KHI7CCIj9OAIjRa1KdtQniEWAzxvwBmTzdlssnAz+AAkQTPuSJcyP6M5R
pV3Wwb9UMw60pv3ZxdspqqHgE2KuDmxlqUsAw0OrD161T8IFi9TgEJaxaYJnHZCfpbOV86ZV1wj4
Q/KRMBwhJvCnZ8t+7VSH1q7pKq49o8JaBP7Prbsfv74W0Om604c4HELiBkru6U2ttKdrGBeMP2At
Axz8Z40cj7TGpoPbyafEnk8jNUSOCmVI/STDKgxCYqVCVcwfRmPN3dY+by3f6y0zaBZ8iE4yn/sU
3TqR26XTJknrw5sNqKOuqMbkPizgz44/VtPTGhl71MZ08dcvg78y0va5ViCm35PvoDY5ivGgVD57
oioIPg9G2/UBAqRZSTP+aqebuFzG6xslMu9YTUa+FW5t8/2OGnMKrGS5O2vKzVoSH+0Ykv2Z7xpO
V/8Zt7b2w2NO9J03ky29kuPWWp7n6bAQUahv1MUhRwzHxdWBK/RXd2flKehhIRrcVi7DjDO3pz68
p3sqOZRd3JJ63E8n1R1LYCIr7B6NF76bot4X9OfNy00nxNVycNoo1YAalS1cMElnMZ+l6UYbfve9
6SwC3nuoDv6eCf49r/m8+LhNooh4+FYC37Y+G6QIEeA2GkHNYr/q72SWTxjB/pvHb4XQXAtQQdpC
b/NjuExO0GVLKY93GCGrNqFBqW8mAS1FfULIg92sb8E28mP7q+GjBhcxSevcbou0lGDWj7767ViS
uytvX0UQy4ZEyRCQYm5xcY5G6TWZU6LdM2XEUZdi6/SEBuX12kWZg+N85u7uErXnj/nbIg9iRjCX
NTSjjnVElEhS3vk+UK0k2Ui0T/KAP1urvOZIf+MuN0kooMV5id0Zz3sDAusQtLNMwkhlnCaBqwx+
Tj1mP1OFIuou/NaseAbalWD10TwAu+FjA4atKIthhaOH7jc7egQX6DoniGBXyNudTSyKDNbk67ZZ
O1olp3dYSnGR6v4O7iJl5X1UP3Xk/Hg5fDtVH48Q4rDkxulsXQRXA26srikHOGwc/eoqwe7udY2q
NOgbASvitBYiY+JB5JNYY74y/bI0kAtdYf4oOeWnnRNb/zacKEpGqSg7LGfXVhzZSwQp/yv6TWsZ
0HpK9RQC44nF2Alrj8CQ+MpbD4J2REa7tWT08cTt5tydqjK2FdsENCKSs7LcI/aXT6IL6l1JcHl0
sgUHgJ/DDCbpMJomJZOJ2r0KF2q3FsL3FvZgPWUmj9f6SI31/7DnZzQK7rR6Zy2kaoZKr1Mva/GU
Xg3Gj0R61G0peTAlRsJbGzIv9jceglyBNuIBojjAB8hDXvd4j35C7YoZaR/pFzEO4GRMWC2IzqJk
7J8Z7yRmXLTXHaUHkovnZ2HVAXuVfDqVBbZjd+3y2qWTkpdLPrXAqVV13cMDOEA/vJQaZ/+5i3h8
cKPlVEwHtx999w+58pSx9Pm82NEQLeZ7bpNJ8HOWgE8V+AdJcBbMgASBJ84SDTzmIZYFClZ2HJmV
mQGNoGrGWdvtLTGnGCZ0spIoArf4Mt2MFX3s0csAxKbdPCrFwclSvoaegK82uRAjvXQOHH5B94wy
re2p+9ad9ldgJadY1+c7QBhUN3ssqdwY7V8+9ic2KIrg0j07W+Iy8pjQS4Vo3nAu9k6W1GQIdUqS
XYGgT6y2MhBU9ZR6LMtoX0icVp32gmjg8IqkgmIDGlIRGod17xUGEuaGX8TJICg9qJQ6IG0Wck3H
W5N7eS/eT/lHPzZrsl6wSbowdL40JJCPHCtGhvfql2xexB5yngKRYEWEzVWrSMo6SbfY8MLOZ8ZM
KzsIo5E/OPPkgEXmjYFwg8mcRD03HWHrTbn200UaYoRK+fIYHjNzkE5yqSzaROsCiF/ROIp7Wlf6
0nKMA3I4APp3hDZ6KSJfcb/p0R8WDHgf9bnF2xoisRr06jK6NLTj71s1JVVNL9IeXv3IOhdVTjHf
6u+sRqAmkzA8+T2M2JppOR/aern7r2/18N0Ddu4lCzm6WO6qPpzVF56HFXEUq4e0tu2m7C8H6NK1
0qQIhBPyi9QE3GzkndInz8nno7Vd/0lGoMdWbZ4aOv04L+PhoqiAQKGb4s0vRKQCdHJ1OJY1gCbh
1mnuYNVwPdBJXpVyzgtW0Oieu+CnBO1rPunddUbNdH1LYZwTAtIvqE2p8oPmKg+Qnbu4EDR77VQ8
UeqLvfuayWsRJByQzp12wPPxFvlpdk8aff3i0p8SucWqFBxJilSG+dJoy4B6posavsVln3+xQ4Lb
g5wVI1SkJ5wcXYtPm69ZkcwXMalarCqfvdMnATDMVoUy63MgYxCs9u9UcRsYcuSJmoohFTMmGWS8
cJSbRgKoeyeDZqp7aNmko8F7HyoWl1rdX4A8GqFHBV1lz8fmctveL7NcrLIycwY0BqN8UL9HTLc6
PmxjunfgICilicT3iSWKvyb4/dwy291FbyyyrKiclpDnI6Zy58CRXvVTwjCwGK7XIsYZrXH6ULGW
nD5ENnGpdZi7utkwQOTnhQ389xsRh9bv7DuIL9iLMhHff/+77XWiSXX9S6vixIw2dguoiTeVYZYu
09UvwjJJ6FeRmJx6gDjjHZaIy6JaJTeynJHsRjVkFX0fNtTcwvGJO6DKsip5wUpDNq3eXS77oQRm
9m9G81FccQ5YnEMuekO4kPE49RE5hLLiYs9cbcoF4TCA9TaTFxTNTI5N9Izoo0HB4W3h+qJ5nwda
rmgiKJwveBqVnMJXhoMbUBNkqu2ko66OKcqffJO5rx/dUkfTFv5PD6KJMNmuYLsobXCFMj+niO9M
UvDNI3ep4+cEq2buL5l8MKIT1YQS730NvGMWDiOrgzdeujby6XSkm41OfP5VVCVxv7JJwxqZnrOH
MZBp6HUj6zdBz8kl//fLmOoUackZ6Jro/k/aOVnFcKhk8FboxYi2f6E6tFwUYlkdwOiDc0smwGb8
L6r/QNd9erR95PN4Z18v1cIenWSUFcCfpsZG8sBMZZNQS66L7hhSLmsQVh2CLlFtKMii4IUpTw5G
ps9p7L8lKSEEAUNIuV3/SvZOEicIVIwy55QHp+JyyIzhQkMWptEUlMb0lC1jbrMdhhdwQQxFHI1B
mA02K4uTy59LB32gsjj4/ZIYZ3E/yDX7l8MXUuMcNjDNmCVoe8CtUvHj+0qPRYdudED56wdtYIQV
5IOxzU/b+52GVF8g7R5y4teQT0xI51JAwyo7EjStuPz0qpqMwmGZONCh3GAXejs2d5Y7k2lUivfM
7w1/ovhmTr9UsYuzS6FrVOh1PDNdBT282wDqvoPKZgCbbCjH/Sm5eWj+Fsp5isLHdviFF4CUgrR5
HDd4NMZIEM/7n7inXzHf+Csv1nov8wk+j89XLMrT9ISsCJVoqVlOQc2FODwzSwHaFwisCqGG7hwL
mNr48Ov6xHMGXaKrAf0pUBAlFND+UazelapdSlbEFmNkaXANhCYKXRTHsm6srA52q+R0MLpXZXTS
5YP60Wxn5FXMb9PW58t/akndiQp/c6rcQ6NnM7Z37+Ks3vuRSvdPfd2Fs2+X7ocUxo2IBaDTjE06
ShAwTrcfxgYSM0LrJ3fLwrW7mHFlpog9lhFUN5iqnqenlvhAMguLC1EKIhZWIBQpd+S6ddKgjNK9
I+a03/mF1W+I33uwqtHVdLhSYgLgnQNBJtVJU9pK9GKS1wHXj1TvTFbC44DfpJlZmOw48yn3WQ5k
Wijv+qsUfF9SDk0t4WsgS+zKxSe8CdeVTWSym8hedVRJtgOTmEBUNffAWlLll58Pg7wVvn0muD2l
/Gsk9EbxTzmi+NCTqVj/qABtfM/aXBtzJf7n8yqFVUdZBpaBJwT9b5cAa2MI474ByNL6C3kuIyRZ
1wIRE6A+ztSeO6InwZfht+TqsHJcPCYORH2o1bquoVwVcW7UUCkvvBFsHUGehV2foZQkSd43I8cJ
6LanWOrq78j+ix/EsZEM57netkoAgM9wCuHS+21UdsG2S6x8ot6ULjV+mFb2m/be8mTVw49bkDW6
ke+Om5855vcQO/yYti/69jVIK9b+i2SHeT6tdFBj6C5uHQBn6LHUAs+RAfhTt7Xy9mExdoWrvlqZ
UMr0JcqICW1G0jZWldSu8HrFA0DnGIiaTZx829wEHdk7zGesHxbkaOE1a2dbWDpYNF8JUSzNInwn
8GEovuteOKkZymAh1EaZwaVrWNYVIanvWEUu1j7ZXmOUl3+SnuI6QHujceZNejx3XsVTkqFDsz4t
MQGnU2uhTcjaPaICw5V3Y1qpy0394VqfBAKFYZBb00SrOuIgFDW0YQvN7DvJflHZ/ikgnuXCKjhB
N4hwRIkXujFYzaGhYc/dfuk1HUDfMy+z9b1Ss7a9guIRJWpWdeu4Xy3M/fgSmDXfgUphgWo12dXN
d5NbuOhViVydFKkFvimW0A2KOsnbKY2jHbrn7dDXk3FuS6DI1AWODMk58/xRb3GiAzWZGAGiX3d7
m9rQoE2AyhlR09AMAGf9FbnY12lA3K5Mj2cbed2wAjsRJzLRdA26x7iWVbkh/IUk1bX6bxjoeV8c
j4OYbPBFrRSPUP+eFHg90DWng0pqOK4NH40nikCWs7wIEv++7EyDuZBp7VD8KpsgdkFWzmsiqYhC
xq+RyGDAY3BI5AI3RqriHSOqMql4Z6jkgeLp5duRlufvGeYWD9y9RyBLIrdlumXrritTFo0MuLQQ
BfQ26CIjkrwz/73jOASt1qHBrhS72SbJ+Vh6vDizXf+DD7lqGrAk1JS96KejwXpThZtV6fL0Nnyy
iIarhGuP1fcOASOkJTa00+io1+C2oy15v16fIg4klOAUTWZMAzW9+foC23TCJkiq/fMjBP0m4a/w
v3YYILtR8CzUz7ySeOEmQQodIrVMaOSjIll8cG/CAcq9dFuH9enF9CYQhlV9OXicvuS3Byjoo1bO
o9TckrmMnOF4N0QIMDzbv21xTsivzuxGl9UeZMXmYNKaZXf95k0E1m5LaBxSgqDU0AxfCdvTtMHY
0Lw22dhOt4Dne23XJA7FE4phJVmIDRc6EG5eaEj5MsOQbBGg22RoibgxOet0tVe6kSUkOuB8T1rl
nUnWcDB/terZND4X8y3IQgexGzl9sB9ObQ55QFVQMg7GtHrK0zZ7zlaAmzxwbtA7ajFbk37+k5O9
D1IhzpZpDgKz4ps7sHAtV9ymB631BfpeWDtpdcnS46y2RiSFbNkshDNhKbIXvrw5DCHV9UgpMg8e
5NoMAPfKyhq4psTwQwiPa15oG8rJH+fa3MXaPvGH74iGQPJqJpcjEzRVMBGhadJxGIZYxzkKOAvQ
BqoqT84pSJlokWDEF2+YPmcQN51PxkcAoOkiPsvASMw8aleO7in1VrNn02wjRBZRSiFPyYjkqXo0
gIwQx0DfyDJuYM9Sph5Gy0vJ0fowOCXn/2i4HOpdyxG6MQBaXzHMRs415/4nVZHLe0KJsnLz8kNS
kdW2JDUAWLWz0QiB61gm324M+y/6Gy9eH9r0hjtr4bwwMhsfilT/hoMb9Xb5F3UwiPe2oAJWoIbS
814wuYpyao04QAMUKtVIf/CcZj/70UMlUmeaKuQLDTBTvqC4smqBm+3yhqpGb6kqL/vlor5p+wuT
ZILiPNDUbTMLGovs6bNd4ds71nY6ObJAmGlpxDCy17PDiRfa3fNvSLH7HbOMDz8nkhIQkf93ylU6
GpXHIRE9uSnQMpTgUEcIjO6tPOLpJuryX0e0W5cp3/5k1oJANrk1tFErb2XCKhioFRwkkZy3xFh0
VyzuUEe4+wx4iRYQJpv84mdiCiCJ935Sq4DJUas5VgwtUy4AchYF5TnFibJLNVO2rtYlLmFnGhgZ
5DIMQNXzKuCGnK/doFMRCnqpwULzgr79tycBFAnDujmzQpYD96SVb69Kcv1Ym8gNc+l+4qkaPo99
Fozpq7kwN1lmwYmKKIQCqaWNwXbEu7+s3hFsPr2TB0vZ3dPtI+MlgHT/8j+l/MyvYsUJEwl+2EkY
5szWNjTEPc3a6tXdsPHfPtD2D3f0T7khd8KjWSVTIKhd+uFSekIiCKN3zpJu7eIhkYW3PuNqZwdR
jnhSat5Y5ftKxeXS1mexlQ60x/pUVeo/VD9sWv7TmzAYCesZC5iHnlTJKA9xwfynY5TyCe7OuS5g
zVr7Z6ynE0irJ2rXqk5u7SciGAIoetYysawVLUsCcbqM756d5JzX6joG4OGe5uiLTheFTGFZYjrn
GoPbETRnuWTMsEN/1L+uPJI17tbbtPzTDjD3Wu+cOFPzUOol2FVMaxUsLKk/6cJ+I7ByQpgm+uoa
jxXvgkbpe9Woo4JliKNmsX1DGmVvsGF4q5YidqQYRX9gPCTnDYCo8kQtRM7VMb/zGh2w3H3FbXxO
JP7BAb6zXiptG2D6Zot7KO0MIt8LCQb3MymihjTkPmpil7K4HwkB/714XeJqdtPkG3GaYPhZo2xu
xO+o9YiIgRvU4KUoYPnKIDHaOKEUKq12xNq/mHbso0h8oc4iJoz4pkaOHeNxeMimgKccgiuZjXou
D1BxTlCJaHwososviLrPIANybq+uYloLdwJZX3Pvyzo8wbCOZwpRtE10S5RtzCMZ6xUe6Jdcb6d0
AaExWqDcDNcfe/24zVUQoOlTciOq2ZQ59yi0mq8NtghPyPJwODPtVkHQ2eYWgUlh28PFrsG6Z8vy
VG8t8hAAxkDPbliTKGOU245GArQTuPadAtWYVW3zo0mYNUXUr45YeR8v4gJvFowx0g0576yOxFTb
4VIZuhaTb7sND2MqDnSuUG8XKuwx1w/sRWiZj03YgySr/FXCPbFpzO28+Auwa/ErUcbZjpXgSDCB
w8dGVSf9fDRlSB7HlCAxcfaEvVXC0FZZgqlCEl3fV9fRtqJUdB0clQQf9zhCwpLMOa0nkdTjMEif
L91anyZYBehW2QcqdKd/8j7oRv/T+aG1N0QidUVOsdAaG0iioZvzBEDKeCGPX7dv/zZvMYNYGp2E
cH4ysirqNP392UooXZtBx0iwLNXNdquswQc5vcpU4S+rd2NK5scu1GyWOCHUfASbp2LTn27VSGae
Av/YI1hlzCJz6S28MZlmjh3NX/GnuH50ROmJ+WL7b7EaF4ttUjeNlmSR1NifrFUgMlZazZ/yA2Uc
4VRatfwSEyXiFPm+TV5ISlefOzN4RbTGgVR0i1I2LOHEKXtEleISZD3XIhsY5xLs4SJUFH5d219F
EFR4XsD/cIAZns3e5JOLQ1447n6xsU4udAb2AJZm9zI8XH9p3Z9aeAEkxacU8XZthup+yR1e2CP5
COunOTbkvqpIXM5t9kYfd6FIj4CIK2lD5O9AyRTgYDBH3LiCcjVUPDK6A9L4sLzSgkTb7Q702X0k
YYx2ijlP3BINtCK9+CvCSza4haU6/fG0Dd3V2BL3mzZs+8gzLF3IkJ9uT3wZK+iKgWCdLsE2GoRr
yrTqZvn6PcGvVvtsS/mSUpZMW6uEV6ER6kjPbLcEugT5Do8UIXuT62sEa3C7tTvfB0Wjzyww6FJF
I8vs8fjXxBLrRHYWjs3v4UyJH1hRtThnVFOPKWuclMj9zogqY760GY7Y8qwuFwb/Bn39KUDbaFzC
KWnMprIRYpXcirbc1EyweXIYEazpdXnTElYPTzKex2TZMpdqpUy7BlpyRFfoDuU1nnidlWh+V6kA
soO0Lif9MHjcJMGCNluAr7ViQX+SYqy6dvjc03xQkCsa5DkTWbHF+bh0OM6YTbNAOaX0M/6NE5RJ
QsacLH2prNA+/JRwWSebPMKOvcrnJtL1jPhd4ppjjeNrUiBoxacMgwohkbpQcZvcEql7qGa9ejAn
4GGloChkPxNKfRhe29luUIRAQ72ZZgke8dfbZZ3bSnYEufOJ+U664wn9P9Fm+rtczrRPaENqXQ22
Gwl5Gc/VnFSHeYxy0ED+gbkoHMr6Te3hU+yuzLorW8Y8d3a5HJJM9vbX78Pu3GOw9UDlA0S/NKGR
f6vCy9AH9UJOb0Rm+k8eQ8BnYGY4h3wGHO7p/yaqZLsxbL3Ziu0+LaZhHOT9dmcq5yEJXgxs8EMX
LCLajwwPHxkqjpqyHw4T/Ig49SHEIrIg9gex4WUANwT8rWw4lxS5/t6U4ovk2n10cSvzAqA1jMdh
M8Ft3afy9SH/a3SEOe/SklkiWy1RIgtsqf4BuXwbNmWlAm7r93vEpnCQ7lNCH1GQlccnw89rPQOV
FqAi0HJfyK8VPM0dpk6GCOs2neqWNeQoJE24QY/4nPJ0u6v0mI/jloMhap29giHblI4b6yTZ2zd5
L7Fbr2hVut03OoCN731+RIMmOFLSCPCwD59+Bopr0Xx/YIwy33D061MTc4OozCkK9b0DQ68zxFEm
d2evn0vgvZpgqZaG11aLWOkWMLef6q/nmUjHlblpGzop3RT7o5joyJZBKKZxzmkKUTkDvJnEtICh
aLrzwsw6c0TZfklXT/B5oezP0PRWy8kwX9FY/Wb3kFOAJbkZ0EGGhQbTTrUeV/JmdJGSwyjwpw63
Hf7iba70FUvhX5QnJrXX8qdfXAVpjtzZMDdexpVYU2RYHvpRZluTxF5cCTwQEiqSnlR07XHw2yQq
uMSGlwwRLo4V0yMf/gwl8UxRnanOqXID+U7/GrJ9hxfAK0T6hcp2ZGLYkcW1I8PrJPac6C9KSNH4
BpsyyhZvvToDrzBBuhVOrgfLXlXUWLyOQdwT+Lri6CM1j/wA+rkh70+eTo69VTy9bElHMlfltpSO
6yg+LM1Hvlsd/e0zu9CBAY/rJNeqjRbCKFFZG7t1SiKlxEkyuDoRJahcIyWvAaWmej4zWf7Zsr7H
KqTxdzCoCYL+Ddd3ORThDnAddxFzauomKQWNTWt7MVVbEq7KZUtrHtfhcooIF8rTZD+ujSJ5tve3
O+krjViFEate9UFqCcoJuLekofRYm5oqhvnyVCHuwHtjKIANj27ivfo6H5JofqYa9Br4dR5phA9y
JG0O7oPlQlMLHXG8ce7KzumHF80mvOMvp1RW1llEgozWRIG7xjdSi68Xs7kv3A1W6rxnJg9QrG+o
FWkizH46bmQHRDOCoM5IbIA9hvRhnz3nEd+HN6Ud3t0HMl0inPxD+Yx/vCW/7mTrb5LDBJyxIDyN
a1rp7c1DwAnfapVhI8bJrHTSVQAFT6JXvhoZ/8lp0x0d45p7XqwoJTzh/ezTa7dG5jQbJjPxXZBB
zSB5Z0jZ2niepl8ca78Z9FrwV7HBMLqHlC6ysAo/EUiUsX2USzXeXFqLk1rkShiKkZ2BNcfS6eIu
TocZz3eyAv5nQmUjQcal+ZVQH6bQb8TYXSJwQjfOUBjMDU83oMydqgTq9nQyQ9hQU6HBFXYNPbMT
5wF9KkxWI7IRsNiDX9w4w9wJ7SDiv+r4XDXWawtMLKtl+6TqROgvDkdgdcBPV+EAuQ3kqklHdvXf
Z+7xg/r6JOhlYGAfcaize61GlwQESgLp83nyIPSjfGjilZF7JZ858aEDA/ORfTqxSCBrC2EmXyry
s9SEgjs35plJBW+vELbkmzxG16OGdmzKtkGM+3DNNiXsxNELvxbznEOHYexb0Jv8STlIoOsDD5IE
TChZ22z0JrNTyPz2/k/p4O9b5gB6Et3gBU3oEy3eZi3pO+f+D7PdsaaWwSoVR1gzgMo0iFJtkONp
POQTpi3Zq5fAdwFQE7BB7UmQhZRVBbvKh1NnM4zOzB1wK5Fp7HfjVddZZFg91rxKvd9kU0Gjiph/
2ChUp18xSsWh+hjedUTggT8+Ut+Ohr/8gJSkE/qTXt5kR+bdQyGcnUHR+gtKF93+2Pz6yZSBnaEE
apSTKd5jXO3zqtT+Sx+5m9ezSPz4uPoMICygDUp+M7S0hKHG06vmTtaPDLNSWkg83pR6p+9CrSjM
92tCJMRUDIlU2amvNe/EktoFLQpvpa7CFZR1+a0DNbA+eSu2Y5waxJFciRgVv7zIoYvOqmAMpVBi
XLtwbqzYsu9Ej4za24HAYHvm/uOs9zK+JwKAVcPqO7TEy38JYVrGdMzsp+re8aoPvOfChaZqZlQi
tbQ7Y/2VqVBR6uYU6WHrqgiKtGufIV0gS7TsEkQQZ4BD4cn+1yum0i6MbrTzpoIO1O32RhcUo1DM
eMrpY64esOG1ztxQPqJRsp6L2vJywLyJ0AuMPDysnVWiUgqBEgitA7jlkbNonptlgCGgAK6UfX9E
Yc21E+AqOAWSMJLaaBVaDHxWUsQMG1PvynmHcyD6RuOjhQ86RZclP3/yJxrUqX57rQh7xE8axrOh
5WYMM975B31haXF/stVMXrKkPkbdx7Bvk07JlnEn89WUM06iFuPnmNc/g2QGoI4RgxfblOTAOuTx
FulbBu3heLTqdeRBben7N10AfpmgjgEu0act85IILRSF0nwE7IL3el/xhu5xHJD64+6vvEosG/HG
XaNwxbWYf+fsxtTM3sIbLi6hCEFzHKNIjJoh0lXAfmxWjw+24WEUn2LTpR0o+Gvdl4pSOcCasyhk
baQDoyujM8YeIhp5Y2BpDAfW1YIj/VUF9y0g3mxBVps41gmzwImb7sQv0y5CCg6EfbS48fgidWXy
CpdBYKDyR4NunkeKRaYkUPp6ru/M9uzPfhPPVXFQVWtRij8Q0pUreEKsRsp+P2gbzZdJUvhuBju5
/d88nXRlCWf5g2ZgrQlEWQaJH2U7W4ChtHfzIw8NR/szuN6ApOgZTzT3DffQ1n9p8WQlk1DhdIMR
m1EsOQuPkDee6/L+wxU3NPHPz9omE4FxCf7Igp3VVyrjRi7bTKTU8V3SaYUCtcYWVEYSxb/fdU/U
sUj0igHc3DWjeCdvtEtUJK2djDhqqnUxUmdDJ1Da5QwXpNQIHyFfgKv/VU1ED5UNNyd6ico7UvOB
zTIQ3qnoxDyyTHdaaNkbFiSdAQIbG3UQlArRTdm/ARHttLM1yEZOrPFv32NkHwMb7fu8Epg8vNnP
z3mq3vatHcvO36bJhoYvcVcRCoDTVHGoDcJ9+RKZr6tDGB2sheLQI+mcSgXlMsRdKwxNdgJV96m8
5zj0A2GFGpFjdvdDRmvsbUp3vW2wyu+jkujwK2PHmxqYCOeUthcIdBqMxUsf1bgDeqHm1oITxZXL
OsDS9Q+J+NI0U7sjso7dfnI+zWcOT1o9L+pI264M0wKr2mMxFa+BdMatx0YGJkxx48Bs5U1zFYh2
iVqdoYqMZDZKXcfW3RFpcjpgloLkanfjjU6i+/wJKUNkFVPFmXqtQ7jEvovFYEycsl3/GADprlBm
8JQTiELbRS66bkLcnQVSl7Zf7JfK/M+2BXEdrFGNTWX7iYBEYk8Oa6oza8GOEDLJCwEq7ZOAm6jm
AhzFKKDUyvaG7dSagKWTUBOWMXLvbApM8r9AB2IrxguMaHVXgi2J3gw+xqFHgevA+iYFPkwSEb9W
0RTbhEXMwqXHW1jiCT40eSFB0ckDDlxxrPtJnnDq7tnL8NIzdTWiY3WQGfx1JhqbMGwy7nzQXR36
gH0Flm7m8k3SDVaD42TlhaCXZGrngXdPf/pdyi/mi1O5UXnbbAylgynWwIFSGY/uIqKav2BshRuK
uFEgRbXREonXLlwPbtKDKB6wwpx5cCv84MlwJTinwqhEyJGVs1i0Quez7JRNs8PVxuzlDI1QIz6Z
tNw/If3uzYS209IDXzM+9aWArA77LCZ2rf5sh+Mho9EY5zrR3554Wy3NV9Pau/K8LnGVgbg+UTBh
uURnVN96ZWoxop/vXpbB5+uolTjJgt62k23hRMsCOLgWjD+XFPOtwq3CVFF68A6uQv6TVS6qSZmu
KZewVxjATw5Ydfip3hLOEjLUZRdhm7aFGYhWlYtm0xZFYnbwsgf/CqcFcxTV3gzgSHrvinyc+1qb
7W4y3OEJgtjyQMOs2pkgRN6QC/pPibdaHSt+0s/rK4k47aHGQevVtIte3C/OQq6Cl2Y4j+yR/g/a
hvVOLhhkmdhHZu9MAiVYwY/HODtki6eVjUNQ95LIQAFkZR1M2SpXtrgyQjenD3dakEtZUUk3nfdp
R5HyY7MLD5p1fA4pn7bg4lkFuk/jx+MKs8EMyMBHZsmFAhTSnMjX7h7xrRohigP3cBjG5zdAmKVT
ZPE9UDZ6boTY0JiRzIP4Ttf7AWaubuoAbzyic+JlyUSscKCTRMKl7DCW/fFOQkomAN2/Lntc5+x8
abRB38Lga4kGkNAnwKrGau34P58vMZ/sqrCyy5QYyuDa2F5tCBU7AwtH0RrtXrwbBkoTtCmiFF9Y
zIiE72j/8kVqgLV9tqkUWkhkFX3XNeZ2pIcbjRSH1CylSSMTUqJl6TehFuGS62Eb3ATRlU2HlA5J
QQXF9/12MjZpaDFFAWaD7YxaBLv4j2vrszLdSoFLhxC1S1ygE4P9ocfucEoYDMY/oh4B33arTRBG
lGnddyG7rxE7SC6mwUvqohRH7KDxXUYJwH4P2Sm3/Ar51NY/LjJ8Xc+vU+rAyqbXf+ceN4A8ksql
znB9pNqjPJDtPvBZAh+c1BBj1MKdLk0ecxUrWaPep8U931ifft9800OTITVU7fAY8O12RlGqeT5W
uGT2YPQBIYDmOT33PcZyWO8Ff93sNsEI7NCT8URhowIXlPJy0odDpBQk6sK3N+T5cMmSjDwkZwfq
M2pvyap6oeRDZv3uaDaXrqElR4NrJvVK9T3YveTopiwHU1V1V01jR8mf/LW8EMPE2ki5AcfqoEr7
xG92B3D4aQaC/3sqnRXg3PY0iiYzbSteKtQvDPbbQzicHbiflt49LPiJ3Rao7hzX/jX7WeKc2XCy
7emLOj1Stu+1L9nWUu2zuEZx5f3H13JogIeY83Bh3wdSdzC4pTgpooojBwHzt0190lCGnPSY6bmM
izwQL+VmOhIYdnPkVD3YZdMDt/kqE7LpaEQ1Jl2GKRiOK6LZV4mDnB7us4G24CJPXvFGji9HDPZV
uinRdtKsT/lueOCw//5wi4mlkr5jVa7SJg64qzr0KffykUtWyz5+ijiv87Uxy1W0b8zOzf4GlGCY
W6m0yLUWlxxN5G5iROpDM64OEKSvAeyBE3hL3GB3WjDSaQ1/IqXnIr0vjAND1oVl0IWosTL8gqS2
T9FEu6L7/hv0Sgk5gxvETvCWbyxSxeOWIes2zO0tgUGgH5WAgICBNYrMFQX47P8labIzhWKFzms9
ijejeHf/ecQVcwYQcoIRzqiNYuicKDCMP7Vobyi0CZth/Vo1t1jCV+VLOqzHc01oPcfWkGYFLzAv
KE6d+FzBKTeHFqG+IUYBevuus039Fo74BO8eCsUIgDXJ0sJiW6DRM1p20QOIHYfZ48z5Dan0uF2K
i2PasHqm7SBlD/U0vnSy752aifgz2tFalqHSKQw3VykTIAYwKWC8/1TLJhpUCk98KvDpgCHxKfP/
PxONYOR2+p34Aeu8fSb5WXBCvpCh4wLQUM3p7N3d/3vTEQrh5U64uq/y/3TjKyXB1JdZJhQ7OtP2
8DuMS9AiUt6OlXstaMz1pSfG+Fowuw7i2cibIv4OAAMDix8h3SjZItZURXt+IIK372tNDr4srQ5b
7qaBjjCPi41WyqY4l8BN+KlkNVhgoU/cNLo7aM/ocgCw/5t3v39T/FsnELPu1fPU2crHUptHXA+3
kzYVK/UdDJwe3D6+as8kJaqM3rJGhq17smAZiFCS/D8XEPBQxW22AOh0ema4ZsgGkofStLWNtNAB
BTkIUnbGO5bCyXE/+S4DFU4HtL8e9fKMFWKcPSXRAtBltPYfWDhVXOh7xh4E7oPxxNthuZ7p2jK6
TUb3qFPhsC8qO9m253VXIbIT5byT69kjAVqVHDgH9YLeBMg0Iy0WS4HAISKpV9n6wZbAk3yrUP8b
kBjm70xotwhueM+KutABvY9ZodjMQEhUsYkosHA4EwQTY0lFQpUa/xUy95baMmYT87FWm+aVKTXe
wKqgnQlsVouk3aMQHcAOmMTb8uCORjihr0fIvOuWuGOOgYrEjkOK3Q+yC3Jq4WioBnhHfo/qg0AS
HBIdn6YiM9nErJI888SQ5xiZlS1roD0v6PJ6EP+mhjFWb8jtTI16EpTpe3J15tmWfQ9XDrRhPmdR
ubTDefUldsXU7F2bGzYiWLXqvsZOuaBLWKEVxhq7FFgJ0fkti3Onb8RxR2bZPIUm366ILADItuV/
NoNrL6mik02IAcOOWR3/D8S4bcWfWX+OE6c0428NLrpLyBQ7Y+ugov6x+J0L+IACYSpq69HPt2vs
TdJUufKlekydvb1uy6rkR3Hqh8p4DYtPXX/Jl6DLINZ/owNgSYqcHwGDJ0Zjdf6FXf6RQsJqO159
mytLqUGmR0XR9jrru/5QN6PL/ZOxjEN9KkwKPR3VIG4dDogUf7kmI85r/vhcqwd900QvpcV/620i
NVozu3A0VbECt3Z1eO4UI0ZCdbmHVNfjGl/b/tBhGCVglwuiTr/LJAQDn94GkEjElUwsX3eT5vjL
1mr4unPA+y/0+jttcLl3t2IvvwB8mEyuZh0LYtKKY0DdgwHIvfQMxn/U1PS6K5PD7FJf+QPwYpPD
ueVm4qmASL2xRiYLjj9hOB7WQLKp/8ATJuNZkGra3fCY5kRPhEkKhmodNlX8Ol3Y8wyeHnryr4mv
O9fkURshNWgaKg9A6NhMfm00vVCmFGfvO0OiEdnFZ4ONOOYd55ZF5hfZdPePDyxTauTiG4WafRwi
DYHNjd1XHxitJYt6qs7QTScxR1efwXBaqB7zUHXUCbQGo/M9RrYvTHIMcQdfai5EkUqORc3bXDBP
ZvTs9+lXSLhPX4FI8qkbhgD6X+JDKrrrbWfNTaM7ZToya/j8gQtc6mnocUOTSRGbkLi0lRfcnJul
t3dD2Kjzq6virhY0+taXyDnhTkeXU1AHhKCmudpSng8+CYJm8vkTT66nQ5ZLIPTxhkImfpiWvStZ
rszAbQb4UTwJOvszwg7INdmZK40OdIxD9yiStvblOaN+6yWfisTk/tyOzhUCEYcAgqEMSLhVrHJb
PTi8axH0HoLK0QkiAiBAL7Sug1kxH1Mc605Jyc6v7kHi2yxE/fBrLE4ExkcYDmeHGmi055LoV3oK
GD3M+oCn080a6yZoupqme6eqUBhz3+TYPiZxTe4HpINo24eCJNqVtB7IDazjkl3nSkhYI6b9FCSd
Kl4xth+b5sAeG3ZzEVVOSphKn/pkeRF3eF2oqh+bqdv/ujQNcwEy/8UROM4aceo7lgvcwjhjehHk
rgVByY22mHYC/Qub6Be0sLYShNkWZ/uAmm9j0DJpNNncMHsoWqgzU5bxqEDmt3CkSrQWzPobYcA9
+Ana2YaIbs6A291msshVLOlA9LQw0KLf59GskxvjoZ9bx7RWFnOdahGW7MBtk3EpSWP3wQWXYbi1
ojuovPMbTlSlEEbHpFPl459LTET4WMWlkN9v4VE1sk/3WRLLrTEIFrF5AI2qkHTEN4LJ4KSY1huf
OyOPFsTpb2VC22kVNJLd+KGAYWpdV1LFQriMRinDO57Wv6YWjdEAX3Z9R5IRpcICBpP4iovQDOwX
YWKehO7csi8E/n+C88WuwzV39EbgoufxfmIqvmYMj28KUWGUL0NRODGs5QWqbZG24Y62AFSeEBNy
/NTVtcpyrkSKvhlqp7x2FF7ZA5f9q5EI5ADGx8IVJi8CYCJDuow+YnHWOT38jVcz9x3/KCrMxbRp
FiMywYqDrrBKzGOptBhRcBgC+TgHiciw4BcFh25wKWSyOPeYHumw1BtTehij2gapK771IPTyiEgA
MmRq0IENoEH1yPpahhAxYGxC1sRg8FTj0vtDYFbU7MQt1N2jWyDavu2UOX5HUxj9PgEr9yTUYDgP
ASunPSQdgzlE872VJkZmNgpvMJCWR5hrCgvEd9E78vocK/P4FqfsFIdcGqVx9O7KgkZQr2TxBrRa
B8EeCmoh6zrJp6MzLNp/oaDCCf7sXcnUxSukP4NppyfDKWlYhVr0WzC/1RkLHImBCDYug7W+L99Y
3cXcB8DX2UOzWeqFtC+KIjSDYFPouSwmzaYVMILlzslPdjia0Ha4xHgJk7VhHOMBnxvTRWfvsU+G
Wdeetzhy/alrDLXxOFoZOuwk8mOelbCWVNZD5c/a7dC7ALW6kC1Pv/GXvq8ME1fdIWQldUcc+MxE
o9BMTTxQGH4/RFp3XH1NNooHft3NdvY92eNX6XaYtPPriTFub5kvatKUpvj6nBlfilKBgbh9auGU
Nhh08zr86Bb/wKtyDdMlYo0EwbT2LYDJbvJ+v5hIYRl0qhdTMi7gCFJNwE7hMa4XbfolMW0jadFu
ZX/UaFy1wy7X2BItNUa3bmV6ExIDEgY7BAU224GCQKN81ZjvVRPJJxBHkqA2jvGbsgzgsrSeYngU
3TgoIUSjgL8WpcJIMtSuisIhbGPk+DrQ7qckHkWttoW/RKof28Hctmnh2U8pv9FnBeTaef4yZQ+v
SetfdfIlmKGv5fbV+veMXpBW/hyJgDny3B0vsAvusFgQenWOE6NKsACrhVHYSsdH/ElUk/WkLOX9
09/vV7yGhLRfDTvQYWSbSTOtc38CgGbreloeaGuEhzt2QPRPf483Ry5C0HcRig/gQNNqSGWKmsic
ZQNUT+qSyYFhFhvcyE83WytzPIjPKVM4RFLpmV/A/stZU0zqLAsKbfHejKXsLdQRNRewPuITD3G7
rHmpNOP5o2ALPOs9OAMxYsh1k7VZNJhoBQKKEQSZ87i4ULoR15jhhv2fz8/8UVZuXLQX5Ml7CY4L
56HQea4usDKIE58+9DGN+CFRFllUalaZIfitzHgh3rZNS3Y0eyjmG28rzTAvj/QHvlIDKd9RgbrG
VIYARybRFbWxTDv7z2uBmeVW1lNThaNKLGmj6v/CU18cbYOD/Ew398OJ1oHBZH3M3bZ8HKpXY+Yo
xu6XbhOX2xpw+NF54DGcSkVcUcaLcODtgDPFDDrsN4ebpzCq2ITDYZO7owxzk2BkXuD4llTBP72S
ThP9yddF7Rs7bCQG/HMsPMRwTOzqd5Nmdnvd/8FZ78N5pAxaNtm+iIY27IpY6Q6luYkq4QmnhQJu
2cy/C9mFNMqUQD2GZyAot/l1ZI3zVtW5VfIkNbwftTthP8MWwdzgzl1duOlzm/vaRwMUJRR+WGQj
yYqawW8p4hjG8ffobAgE/+rezGJIHNwWP2AKzcflE8SbUUQPaNQ9UJBSg1zJD5ACZYxiUp/JqgGX
ceW5ufj2kcXaNzBLx21tUHLHUrvAqCYlJl/ZiaToN3IzXJoOkGgpxxVdt5m2ux7LAT8v8H9SgBmw
N+3YcUWKsQQBhg+18jnNkIwE4vmg77jt5zKA+gOPC30c/BpITgU6sLKbH+1tds+EXZOpy/WZek3L
yvTIdOzy0mJ0DNTJa0pTF+Q+MO8AvuGGQRHPGSrJTDf1whuiH149g1d0j9qRXKKzRqCSjeyN53mm
w9hQ9K42miAgkNrx71HUaRMjnJCfQqsY3m29kN5OVdf3pTVkPwQMxZzCQ+xHioW+44EgqzR2dPVR
aO6i/y9cmBRt1s85xk5f85ravLPOqHCORWnlbNb9x6QUl1CVMe6eH5N8NNqoRJdyJpp9ml5xjh3S
XsuZZSKDL0S+skZJrnZfsPR1ku9w04j9yDdIEnxWFE+A4UsL/Bg2d9ZxPnXTtyRKtbQr9X9Jhk1k
Lo8F6DwY6G3MKeexrHoTz3jezA/0nsKo34+IDXb3CpipgcXHQHt1dmIGpZfdsD8leY8mdYE5cc9w
b7dEGof628AtphfSAxos/tg1Nvnu8SKFM62Fg2zdVB17UY9yB0hi/JN2p/BYUxYek5JUYsndIDyQ
S7NJ0qVzRfyXO4RXFs4P4VDhTnGMdx6/t1yXEwa+eQhikXlF5NA5jZsfqaJ+RfrOk9VLnIWlE4iJ
GgE1Yjn8uQk8yr7C5FJzHWgzRLZoPbV4aIGWXF7OXxq/ACmwNhXRfNGoWzyV8Ng3dY7iQ98kN82+
hLovae0/HGgejmBxIqkFyqReLp3MyJMoiCRuMMrShO68bsKbLQNIfiuNnYobYZRgQ+7qzTvhgJ6c
Bdnk4P1cSlBF3nl3/nVoIIRW0AbFMXKZOA2M699lNV06rtpOsy/ZE3vYYCT+sAGWJWDGInTJSEHT
pkNhNYqciSfJX0bRar2EsPTkMsd2lWZGdUurtpluRhqJOXwZqDpRy8LS05ZjOxP6gZlzijYvijsF
iKZtj3HOWtuj/TQpMnPGF36KxjHZd/Bbh+0WJomBLUOBNlh0+Tkeq9UfJEiB6gP7XElRVO6aqV5L
ob+kboYxl2Px0ej24jhmhtDc2LGzSFPJkzVRXyI8rKEZ5cfXoNVwYvUBIqrd2zp9rlfEhd9Iwgcf
0AbC+zrrzJd+qSp8+B+t7f6p2p8of/jQVF5yj5wCMQMJ/9L+eP5oZISOBGXwFJQb1ul1QSMe4S3H
V+kn2+DCintQmlJth67pZj/9l4NjpH/+lxblksbyWk+9S7Xb6olba54DkxwAd+xESuonk/tYqVsV
a1JbSD+RXUH1jufFIvrsb6YSaupg5KTWtCi892/ugs9gp5LXDM3j+6RDzy2prpvvDGOS7bQWyLPd
4ABBldjH4WUUfzGrH8/Nff9yo8jICLpjpOicEbYq7qKB57MBzr1EMoNIw2Z7np0wh1pOBIqUwsmM
zLfSfaKei1I/JYS0509CcKedPdhD2EeqXe5uCGYNm7Ui+/AxPIzzExbsA6XaEI661yIEBK8l891/
zExsJfUD9g9G03NUzeLYcYNgYXoo5VTRdLqly5JlcZsU9z22VQvRuwPMedh75RQ8qfgpks9umi8h
nF4Pwg6Wqqv9ZAWnw+fgXMMISmYjrRl2cjEDhbQBTSJp20Wt8cXVqcBl47TwJ1IaTjWVNkmfCf8F
letfLG9p+GBRuX+hXFcgfUg7RJfLHBhTgp1IR/Gt/T1TCdMWF29ASv1mjhuJd7pnvj81hLKjl3Bu
Ka4HnFVKR0Jk32pK0+G+96V9oP4ikWZlBbo+4fbFknBwhuxHTrDixapkjPfIN09aoOrGvutHWUoq
sRDkBW9HX2sXAP3p64n1kJnlJ6aioRc/Fnphcu0mtCeOWvPtIiVqGrCRXLffoFNGgdGsjUc748Ws
kzZoRmYcrTykCox8V+yDFhSSDLMQ6fYUa4n8ipcLYwzJwd9WKc1rLhfjL7SGjMQA3DqB7zhAx99a
+uW8sj8lMyf00HHrJoj3CF+cq8a6S63SeRrhH1ytgKs3hgTSr9l/zPaFVzcFIP+DE/e3x5ZXFmm2
8yX863axx7p6wpRFyeDa+TwHASNCGwRtv7AnpjtG/Z2ASywrCjlFhL3+nZp1f/HPh0MkzQTgTb8a
FejyqnAkLsPl/LH1HjYp0QjZM2TdsdPwPMHx4VeiYuk5nJUmqDEn7UHIHQnyirzbY9d6LvNttRKA
ThUr7/AlsupwT7CeKZz4pSoUYpce5Ii7BX4DoksXjXaNA2ydTduHZYaHmc8V6fYcPGStCGnKOWqm
E/0a+S4JUeLbuzE+wAjG2pdxbikTr7P/00Qccrn0HJqPBVVIvX9Q2/f6YjBYD6agBHYMxSPYsIRW
5RegupyF4JiJd7+kSUAKkmUu7AzNa7yUaEsUgEyA4UVaDTt5I3/was+9qTOwlLt6rAvcMTLz3YW6
9d6iZj6NqBgsZ4yp1I9PHiRpcq3cOjYUWApGGqifWyy4k4dmLOQ3Ln7I9GVHubjDVGBLAoDRa6RG
dy4zDQtdIcly8/MrREPoZ2hXp0xWuaNMXv5jQTwF2ZGTp7V2bIezcOc7hZ6rIrCwbivuEBhZfhs4
YZ105PIV/pZk2czIg8bgRRYes6idstRJk5nt1raXxsl2D7N/D16SIxSlW0JYzXlIfFpdkhDiDhkP
GRYX3T+o5u06PTxEv79u5W0hc76qxjdIBwEgLzs8VwFqyLfZUpqjWyIlULdgIz1Wl8bU/OHDImIO
dk1qC9wTMTOKh4njMi651WUh9IplbL8uDhu2lUaV4THMY8snvBYDTIn8SGvall4ZzfUZJQGl7tin
/2BZbnWeHzHRCRg4cXHmJ5xYRg0iYjWtO3zY2FJJNde9R6Gc/XHyw5oe3dvsOy0H9aAVIkn8CQzX
N1Oe6Mx9KJB07TCYDaRmqxiJTQhxsaacFyXutM4PlvzG+AUAc9LbfiE6q7GqEb17+8RaLRleuULA
jaYA99MC3LlcY5TW46P4a3pcQwkasnozbjMRft91TfqiIq4YRGr6U4WkzVeHKTAcWoBK8X+E1DlE
v6m1I6CfHhxN+gH7dvIt4nYbz/Uyjv+x/aO/l3SwkKW39c6lr8m7q4ytt5d/X0CBoqawTrEy8HRE
+0DvN9IhqEm51wJJoJhIL/1XEBWwJsGi3ISS/TSPRsG9E5XtRlEi3dUjBFl26JinO5r7ly+Q5qjg
ky18KdCksKHJis3HlcGb3RBoX3uu5o0epLv2leEX9u6mRuvI8/+zE+neXvVAvGBV7gJ85hEPksKg
kVquY7JVfeieMLK8/L5bhqalX9FUOL0NEQnbWFO+85fPIgrfOkLKxpX40GT+z9c2KjUvR70W0Hl5
Ej73WlWtERMf+ZzpoPSz+NkH//vhgQPbfkbkHY9q5+qIuIOF+BbcD5NB61EgRvoj/N485twyocDr
o88lsXk+jVSO/gvw07jdmXCWJdAJ+7/99fEfITWBo0AZatovh25VC4cRtzeMmQDGnKcdCDyz5YLB
FERqY5JawxbYj2OY7PffvgPfMMZgSZMKv9aIhILDJsRQzJO/BntUItU/QhPhvYMtSx6TtwcAHeGb
el8tgm54NJ/5vhAqTlQpNgKEDFjHlXGGkh8T26cnB6mTFuD4Hdl70schttxMdRsTepqkneiQbW+o
G1MPLaUxwoZkHYLcZvc9g/h7TPs+k9rlSjsIHB6Ze7tcF5tHN77agIUB3+krjSrMZ6ZJ2QcpUC+8
HHM1lAhGIj22Q4MI2f85xTtR5ZYYj5eTLaq0t0Hwj0q+1FNwxU/O/Zm1k3BdDpxDCSKxllXBYbTl
YH5XEPcFhYg2WB37DIqYKU0OanZwgdrbaOZrQFbmxqd0RlXkYRABPR2ezXl2Un6FC7TwqhMOp2jf
dVVhQGTEXfkyVxmRrZKafZ8/c8jN6Scd4C7QJR2TWbcLa6LIn4T8puS7LGJCSTDl4XbB/QdVrZB3
7xpP8f0cNFDQMIp521Cdtnq1UaBhDgCwwrs5lKB6QYy7zIxADQTEh2Pe2klmvTZj1aHXRtBOPoJt
I5SngxZmiQi5vMmlZqF+iYWG6tJID1Q/oX9SdgHfxLZ9aigibbHaV3uRnwZ9yicxjVPEwxVCU8h3
uTT8R9zPDWBxsf4OHvlvirLaxM9tZzpUgslX8lvqnYeqwEwSGtfimXwl0V0GDpHOO6IBIDQ1gSzC
JLD2WI6/qzrwSOpUTqkOF35lroK/Dq1mlvFGJkOsbgRMYXlbJ2SvBHnE1jmrWnsPnbfNTVpSipvM
byCdlZOOV3uw9NGcWHZoOj2lBJqfCXSZ/iayuu7tH8DQRStkf88KhvXd2NFxisUMfRSAfP4dJ1F1
+ObtLIxRKMd6crGT4L441mI9pcyuFLuaRD96i+4PmPls+Rh2dfAocxF1irTTojJ55C6ozOjEH63B
VZwz9s4vfMXGbQqj0iPGI4nUHg3SsCZ0c9CT6RqSRUNeL6cHuVnS+hYhmyi6L6BBoZh9avbCo4E7
fCJl4J9GqscbZdASLWfRYnS7ka21w6Ot9D9RlpVmhC1w2V47OUUE0DBkbPL1D5t4p+FDO8UYUI60
VsdQ4OFFdtXVPujdM1EsVXwteOWBPiQpuvcq2cZd+r65MUWSZ5sPiNo5ykBuABFTidYPOVZhl7h5
sM2XjSloDe7ijJjkrwzkzPnYD4mJGDOrHKYc7PPd176y+20eZPSPZchdmE0wyUrXo23cf6WJoSBb
+TzFqv9IZSmjYdkOlECn6kpVcCm5tqBMcYLCClrdYwYaVVmAZMC5dum87P+AvRXvyVZSXWn7lBb7
aAEcnhJyTRdoHyjVUT4qwz7eAPW7kqO30dTEm1Mo8bCGLe93cW0up1mFWy4gvOtJGl1b+dCBRJPu
0zS1bKuLsfBfSETF9DgIOXltBvfoFt34AOByyLy7XDYOn24VBtriidsgV4PgRtOS930mMQOBDLxT
+OWBX00ntirk6S0m3vu+3p2C6HdGFotA2enySOIQpbL1Izu6OyDD5WuiJbFU1Kq7ArPOzqJXEL+2
0v3sr/B5eyB7mYunQysNf1tOj1kbdVcTSKgu2vgshgw51aGUsObFLIigHEYw4BvwsM0hj6x04By6
DWNl5h5fGHX58TF2xodZcQXCkiR8HCiDFmrKJfroFJf9T3gaRIfkSpGARVR5AcvBA8LFVVBmQwIm
SXZk82uZNn1YfXalEw4yNTBKNa19KU4BAoUG1GLFpG2b0NYMqSMaM0DYj+EGaADX/jA9YDJ5ehYS
Kk++wjYbSw7TFqkFrJil4QmLGg5fZSyuVblyqp8YTropAxn6f1XTfLIvGZzVrhfHLrmBzyFqigqm
DDgIBVjc1ucrH14dORkfp+35w2yfHNjuULRjIrVajkEMv7UsNv70QMoNT55yweilJAUsj6WF9+rX
MH5EjllgPABP9j2vsSUIV+LwWE+UlNEe0VPlB00OYocNxNdJjiikLSo3GFbHBLxR1xpUnvxm0rIH
ZsFmdxdf9RWkIq/ufAi90kGgCBQULhjKl7ZjeOTaqafgoYTIB7cDTlLRO+SwXRQcgeduasbE98MH
C1NjtEidthKF4DafMgA6XEqnngPFVMjpk+NyXTmkH46ez9Mp8B1YibA2U+bFCRuJl6C9QGY/9UtZ
J1pkSWZGrxZuFSlwUPwzJdqaNfWEL9TLrXdOxL5mww26oLXN+vHmQJX3WccbwIOXE8MpqMVJnEQz
uN990OtQnI2elP6F1mFA1w5Bm5L6CHw5/rP+CSNqstY49mGgK3u+xt3yat2gF67pqxeBUNXli+Ah
GcZfjlIZRsrWx7rdG2VVuQ1m/PUpL7ZN4dwCD73jOXiT0IctCb0xDACdab1Wpd3DsJKjUDbuqwWE
ErftU70ZsR8neevCKzhK05dTJ9mtU45xJ3sBvGsh+830bc3uefOdKleJOC8y6JKWcfWPkkIiDVKP
XOl03hxPVaKcTcNHDGHmZ9GBoxtMf+Lrce6sQcdj702ldXole/MxsZANcw4VeN+aVkILIy/Ue+pM
8AP6Rr+VM6oT4ZJQZyl8/2RM1aqbQVtXnAJZ5r1wazYAldcjX7PQC1JtIz0ZFdS5CHtctEIvxPIE
h2v9jy2eguxj+t0eflz19WT7Kd5I4bJ5SPiUeMDba7dSw8xvgumP78BpkxtxVH/Xe6/MQnYHYWcV
pBvadDSYkOWy5sc2Fqf/Q6CxE9KDiDvts0omEuJ8HwhTAyGbyTugm+uyI4Jc3f7r5mBKbFOEq/Cv
a2e6pZFHiZhTgN9MIlUfxurYextrgVHtym/DsR3OpbXkq/mKiU3NktIdgL9G/ae/dcLeBB0G9Zq+
pVPhwooiFJcNaTmtxzZlmwcy7sXR8J8Dy2oK/jCK7BJXRAsH2QCFNV4c7Digk9iiI+yDgRacScXD
KwwanLSzoSFVSlPWLsUD1+gYE4hrjtn+xHgquGsI5/rrmV5TzLeH/jQqR9CM4rq7Aw4tm2FxZ0ww
U3K5mQbveP786AJSZFF/I3HYxiZoLljek1w71kZuoH6dZ+VpeAhM4Go/vjS9RRiN+pWm9FjRkifp
BHqehYd/j1H8jwE1bW5+nlHRS6WG8TunoyOlzO2aUUVQaroquPh8je0vTc86BmQo6LuLt4Kc/i7+
PBirH+LSZhyZUz3NPKzXH7naBMcTwPe38FeB2RFelLX8JojAwlLPx9lNdllnymAbJ137ExC8yvTg
40V/iL5eSCpQsy0Zgz/wzJajYtq8TxYV9Vab910pBN4OhZsPIjKgvcVKClgVcsDZO8DdSUwmxU7G
LbWFUCrCapMWOo66mI9gmXR+gJfI6nmnBYey3XfgLmdJTQCwQlfMTgEFV4sr5Ukw9K1KdZdyNEfs
PpnH8ZUDx1mNgYAbq0AK0J3xxFs0dGSxzdfqr/70XI97NgRtUS1dtSWz/+9/6sazc4HaJtWAuhef
AtoD65XXTRD5GxIaVrS+XerAIRMRjcmHBG0VkM/8ArRplPO1qNnijGfz1kFL8xDQpRjMZKJWXqh1
/X9c6R7MiLvTq+giuEz00HcFzZXu2ZmBKz5ELYDpMChahRQVTc16W6dG7DrsRdaPqdYGD0wUbnkH
vXAMyIAZxdiY6sVDKGLKOnnoIdJAzYObg//vyjpEkpEB9BhFJ4S4DdwOBHeRyioam1cCIE5nOB5s
cDxcwmvm9+vrmb2zfgq74NHt+APEwMMq6ooFKTSJ0jcJbrAExLW8pWWPA2kK3ULKpuKJQh9ahjtB
ZFNwaCBdA+AOurWf+0Iz6wLkE59QpfiTBXQH4yMpHi5d72++vgyrycA5SIWyMqdMTQwt6amwOa37
IRkWuQeA/keYHue4KnoQgMdtK9pfMq3J7IfgatcPF0sDf6c/L205BkcasmpYVVls6dYGEIJD//c/
PYmFXjbCw818cjRVGK57FhTvl8AYR4yNhGilSKifTmgs5UcU0BKov/YRya4diDUDyr20lSlicKmk
uDXBvA+nj6zQLT2mAvyMi6ET7K4sh/AYV4w+aDmxPc1CDpkWTFHsWpyddCBqNALBcL0qinMFUQkI
bFU14jXmaAUM4Mg/zemL2KLVDzCWvmivWzaqR+W+q6BTPV4ShpPMZNiqOHth8Yc8pEMTuc3J1sCv
Y42s4ZxnFfMuLW8jOjYC/BRbGwp59nJ9qVHjmfruusJUspjZo7Y3oOos0dcqG9RE3DnaR6fgpGOY
NuEpSM3l9dYtiyZJtpY72yhnz5bmGBPYvBqSvILD03okWXDcWSfoi9iG5R9WhQJtVVLU7WgsMWCj
yMs5jso+WeYaYY+nbUpv2rWVl1nklzQXFUOT/MHS3kOaT9yHhs+WrSp57QNrX1fjUXhXi5pEe1YD
MYl2R7sqG+eIMHc4OOh9nrNA4Ep12Yww5pAlnLRqkDiSjOGS9jyrSnHXJpCRWrq4UrNCOyyMSlhN
++p/tTu6zUI2lLXxS2D/dgeQB3r+XIWD5JRmFK1dlIXNGhuPak1jUy0GszhJ17VcrJK1gqMlP9FJ
9WATcZ6O/F2YjoRRA/yduBco+jQJQtY6d3H4fNwRp3qPDJEfmM1K4BCc2tTN7GhxnbHXAjeMrMNV
kaBdUbtlzff54ShRmq7XgZPGFfirsM5XL2bDxeXO7kBVOcOE80DFrBbHlTrEgxJqPSojh/YX1/Ab
ox3Ylal62W6tt0kBjJGanjTBDOQ00pIBYkzl4fbcXX4wIfmqrxIcHglyCiWvVxofk098ef41WDpn
exJupCQfDYDD9WSca8g8vpckGo9Czmy+1gK9nysizQsWmO1mHzkp7f731nBBi8PGenDVvj334XJt
Z2Mikx6r1mK/mH6m7/sVwqIo5tzBG9okHTxzotOGSj/QAS4Nrv10/3JqTkmAYB/99RcThB/HlFF9
bLe1EJcFLkAjC7Z+vTtFlR06spKono8bvAmhlFq35Pc0p3ED42xuAIx/tESiQ6aFbv/XQiBT0qhM
UT9pKSenW/aUQ7iLtSzHodQA+8Fh8Hop7GUPKpgvlbVJQ96y+MqUjdj1eB7wf0JkN+E8JeX1AmmB
g0NOcAWvgtcGF/NJRogO3wqclQCbTNV6XQGezVJ1MMT1c8rikxg7WrceMWPTfK3PWyD3deO4n9H4
Z3C4vOVYT7GIUMw5DJqoQiCs3jE2i2SbY1pnoSplDieNVXS4G6wxCqxziWQmoOFyoFSfVuk+XBK9
l9IeS9l52Wv/26CQ/WCe35l7V9NHjBrjWfg0LqXNVWqif3dJ1B0Iab59lmjYJm/N0KLkyW5uYyK9
vNFK/jwXjZHJvpPSEy4oqvnanvzm+SZQQDDQMd6VeO38YOrjs9uq7CJIOUcPPKR9EJ4RWZVAQ+VM
twztR8Z46uDOWGFDmH/HPhYtwmdT/nAVqCwLkau7t3T0RsWNFGCVOVf7CkjpOeOx2m4hnS2s3N03
GYoH38g2G7hTF5EbevV7vPOLJNG7EzfQhd2iLpPMd6YUtDg6/OK9ScMxMT5t+mPcLVZKEIKIiZHd
3bjT/O6xmtUu9zdL5jD1rnfJ6khfj+igrmqrpNK+7iXPL/a7WiXNGlmJ+xlScWiJbgXKgM6cF2Ka
8JzoBYIc4AtqGd1lM9wvlO4UwIL5nAs00cEK1WI4/pQ3k+yPr2z45B7n4iv5jNSiQQp9Pi+Rn1wf
q0ap4lAe1H/jAbaLt1b+Ztxs/HYIeDWTZJ5UlCH2AoecK3eWZ4bD22rGG8VgPy41MHIK33wb26fR
0ONoEsX0mvortOoqaaWwujgRB6mzTatY8AEbUEvZ/TGXPnyCOIs22QJXL96RyvpFnYJLjtDsCgW3
Q+DpE+Ka/xmAUZauM9pPZ4I6CSgyXSAQwjHqblQXQSjeoNPxAyiH5lnSPB3JHLcIbHtQF8IrLWYA
8LBqgToEgswVtmETJHM5iT6aScLAxhcrQnbqQGziXqNCg3aACWRMk6guxHakSTcP6sviaGF9WZVc
+k8xL9g+SJ5nCu2K1q7PFP+xOVzXEs8kMTbRsDQF6D5mD+/ADiOtu3gyCz+/LGUWa4tcQV9j5i8U
pes22AVrgs+oxZLjXJ+gMYdGlJnT2X2+rrhGz1bXvTfXwvknpyQ1ZqKlimPOtNA1DnkWJcnyp3nZ
lU+HazspBKLLkBTAyAQ4LJmwlScQo3Cc9i3JWsaIWZn9tVXoJjC5QacPhmkd8UigjAUH1sSOvzhE
Mmv+j98aA/5Uw6OB7jOjrapaEqxbIYr/5qNUQbYG6v/+5vtjHo5BJeX0mwo4f67aoJR6UUDoZszZ
rV0nzrp56tZUk7WkIx+DmD1boGWxO66t1oFhZap1u+DptmpUbM7+D/IrnDmOVXxubdYRE3EpRz1L
qEZH7TucAJEkV21nII4yDLAPsZukxcMUli/7Ghmd25UB//OhZ+pOUhvcmRepoIOJVN3j6/3s5gsn
3/vT0ijQ/T4IM/mfgRbl8WmEoJylQWbVb8a/dTngq4xu3G7UI/GhkSJFfwp6LJTDN4RSeWN9WpK4
nxPYumXtw3BlxIKqi7VeOrUFlj3C0+Fz/VMa7h6Q4mUhWnf8q/RoJrLWmYDmz+OyNL866fw1AChT
MwwONWBh0W98Pm1d3nuZUkhGfu0ADHI0U+GU9eAzFfpPN3t1fDixSUi9j9ouLsTNT4ykKcAaK7Hw
ux76RaMbswfQiAiHUYn8wnE6RMZUvlTepMtWPGDvu6CnAMFZolHauuhPuhVe5d401DSrmb3y7eHQ
xyQHNM1yTU5xdFf338v2arASeDYF0zp/VgPEQGWvvMXiO4HSzXaqFtblAA8Y7ADr3LwQlGrrqcIK
JaL0iAgLy9dMPOyo9mR3ed3mxmXQ8ldxR4/3jSHX+eYEFpiFf5d6Bfjk7x2PJ9y6878HG9kfsHsc
k6iBBCbjmUxAq5dHS/Y/r8zl6qDOC3qvyBbpsf2O2cG2wZz2glTM6K7O64b3xyXDfqZj5sskWXpL
JCatkBofzXRoXZZLE2PzLK0JFg9d+Kx4FnfgboZq/MdUid/PWxzGST1E73fK0pGX3dwvefBvbHmn
pBQL66c+W8hT/rZtdrSjlL/jBIJ2FUJwKnPq7mgV3SoBuoA8D966XkpFyd7QdHxk4ihEYxuFlWtZ
TVsiNxJ6bx8qtUjmJU349DWOcEoka45H3vicaKddPcZX9wXUqj5PTrOXN8nFRM031RQyfMrkRkzp
XB2hsjCMJJ1AkpWue3bEbA4LRFft2cZ4Q13bAiCoJU4G37mGw/CAZj+4gCJ79gaNNMw+jzYjnRmD
IyQUKbSBK5BAGzdjo6wQJfG61x7IxfLmJZqVZkz+nb+lJh82EjhEVk1107lJFxeU9DRqAsYoVZ/D
F9p2urRHb4xBLSjYJYVVB+fm2J30LSb/pyv4sQAm96Xfac2wVem1XjI+Cxbbrovyj9rS/WNfQc0k
Pob6NGRVglo2Ntr9vYsrxo4aTSJ7tV+ZzIuG0kHDmE79Kp0zObVZTmuS5jD5JtTrwAAZsbx2uMMF
JVcyfYrDXrrsHQpKBDL+9t7OxaR+2F7Ac84BFcMAqJqqhH6rAU3XRIumepziXbqV7KnqxHKmy35k
9/lo4SKQcet/Ezqv3HflhycYQu3fXnGD7T+4gK3MrH43JQxUlr0Tp53bDS+ECyF4eVSFRF4TjRAe
JkfobaGWeTSjKDr1S35ZYO1bRW0fTQoO79ed3jWXXHFcvy/Uhi8tCIyz5PlMSqErTx0fGqkiTjqP
VaYAiZC5jclYEuA2Z4wvw8FJhlKVx2LEDYulXW1m1fI9pS6zLCL9S/t78eZYfvuUflSRtRlQTA2y
K6F+94KdJmmjkpfBSL6uWtr0tsY1jg083VCnRb1gafBKoyazlZSiT+FlBmDWtxJcsGReyfHjitJl
kcl4NY3wc0le6A3U2vEG0ILtqCP70/ZLoLbY84srq+kancKb0MugpaSpXYhd7oQR2oHeXtffiwk8
EZG9c849nvtve6x713/MsgCxDjdM80i07ozKrTJrJVj/NgrJQVPm5csvDLXiIE+S9EaVtUbZvrpI
FjF4AS6e5/k8twMubjMWx0YLzS0ZPSKSAvvR47oVRi2pNXJ5jv/P3lzPLvnBms5a3TDl8fru1oXx
b8mTy01SngPYuPni4pIVidXOLw4iOaabaQ5aXlz3XCuzoi2hgKcqdnVYPpFEW6wgWrHfSY2hkOc8
C6IRPPhWq6VxGzjtR/lDoZou+tqd/K5R75jkiUgDDaCKSLXyCTEakreNAGkMQDXTo7gO8tv0pNTz
vWtq1MCE5ggYngyRnK81BL7SKb6/LD4PCZrdd4ZCO2j5RI4bj5qyespmmBw2K+bvdqdG4+hVxvXc
uLfUSxXKtWQeIvIkkFD9VJ2hROyhiYBR0ADJR7QGmU9/BO//oA9cql0DzPa/AIpmMU8zYZ1h29Sa
YrId9At2NPuMKEhoTmHnYCKMZ+2c7h7U/tmq3qcYqFM6R5tA+I00VGq4VvCzHqPCyooe/dgE4Uw9
REBMlInn8EumSaRwiy9bjy3xuqPDWUzx6+5dzvJNZnzeDsjzlEh+pCM5SYUptZAd0Zq2ap5nIrDU
I6SC654euMywWLgIvr5xQvtBPh/HVL+jUbi+AJSMUEhBJK+4+uEsnwsg/qoU/4bsKqZCQ8VkVEHe
1FWoQYkHffxaUlY2/11tbXNq9w6ZAj/5408P5ICpx8my1Cu/jOnGAKTaKtejOee0NbDnPBuD+KER
PiZvnvKqblHvKSeYqxOX8LgXIjY2sCpEkIo9tFcxwHfNCv+ppUFFrS/qWXXgRevrepoFFnsE5pZ9
+nSlQjOflmnpk6RQp0P5ujijxRzEyfu1+iFbs4vttmuRGsLFIX4b26e2JdothrGMN0SJgl3ADBUZ
Q+qrEsVYU8BF5nLdyeqnLK2MJhQu1w+DzpWwiSTIpew5mi6baUn+fBHIDsvs+pUy7Ch+EQl+ZWJK
smvEe2796IZtyGSNqi1FI0uvDoMEi16uJSbjRQTq6bFTgRAAVfd9QIiQGzl3VKn18Hau7ZC+PL3e
uCwB3Zb3RZpB5PTQfaH1J4XxPlbnb6Ebhw4jrO+dqNfKVYpGkzWv5N7hpIhUziriaLFtfbxwGTiE
hnvR3afuO+5vMYP0W5FOmOuDv2J5D2uX5BPiWskcTtU5RhVrCAocr3P8+jVEHuw0esxES51IUvSD
cJNDxllIFVP/NbWB7IYqHwQNrpgJ4SYv5/9VOKSAW7Zy5e55vRU6LQPc/3eAhGt12EXwVlFMLENJ
u9jwA/EKXQP17fy5wrcEcQCq0qm96B8jGSnlCZcSzMZOv0a0pmX3mY1tsZ4AUcID5ICsJaiM0AY/
laeF/fJ4G1TZX+NKG8UQVkjyOy55l0ZzdQcIOl3nbIwjeAMTfHKSbfRewD2JBNsMXTEIyUm6yUbC
LKNmurZDNAEcf55bleSgBk1vHiRvxuY2kPqJAVGHjUmDKeur8lGpGpQLhHHqm7ERcKIUFpE7bBDO
5bPBMQ807DP/d5Fp471hNyl1yN54lnyeBeC3vFfcH+VNWOYUz5JYl0nA8QEpq/cEH5Q8o72bPPro
FypsyOYq/6OoHelYkPO79UAveULlDdsf9yMC+3YkEpXVrO/aIG2uVYgHAhRzhrrRsC81vDo/7vst
dVCW5syiVZaLjdj89Laqh/5usGMqCaEPtM/8/i7E79v/IXakjoUVyvK3/mPurrPHimneKpL9JLTx
p1jKEUUI+TFTvMALhgwQHJ6gXFMGfWvRJINBWMkaWlg/+J9abhH61L6wIZmTd1GbNcIp0PKnq2dW
uaCMOK0Y73KyFYmQ7jVnDr+uGKAmF/qrFo/vpvV71hPk/RIvhljPrpYaHpa/ApsOO7qMRL3Ehuv6
vYgFQeEP3dRjxhHej7RKPJpd1Wzs1oDClqivXILuZ5cB9sQM8N6pJ0xQXuiB9rgVJEmzqoHV6A+j
ay5wFXFAT+PgftywANx5TPMWorZt2asAGL6HMfgP0Au3KGV+kEuZzjxmgXtKJ8AV/a8tdcnuDky5
yHSSDUPu3qRUKm6NxDoH3LdKGf8JZ7oaMo6EhxuzcN3G0OB1s4afrl2tEqPP1e4Rc1QD3FVQ7ZrY
uf4MiO5glLrYTZjjmaIl+0/4GTvmrizLG4fxLuk9cPwsN4JsMqLQa5p+HJaD+sYr6T02H7b5tCJ+
n4pkivs200UMeXC+x4DFFpqry7y1WgZlCHgctaKVIpAV632R3G/fe5Z+lc+oZSbrNf9XvkhKzdkC
lBL1nR9WOSyvXDqKMJPu4ZTj+2I1yOLDLTcYpBh8r6TtAxP6IqAFmLacCu6hWoBnvlC1kQRoNJ/X
Y7EPJ3cvwzA0B4k3EplHzEuQQ9FmOLSX5VBVosQ23nQ30yReX1Tj6p/s4yRw59A3Zp60bD7zoJ/m
B3m+qdz/ZNMl0QEx8xm9Qer0hlhNBhy9rViJffgSbaFfEZnrgEabLa1r+/DMJLRzNqd0TyoLFtFd
0PCuy4fl8ADWcI2stjUMnjM9lmpMr9jKqe5JhyuabLwrkkIXU6KRGLsunKiHnmyX0meRLGlxJO+o
gqOcnAWx70G4JImBYlTgxbRLiYIqemzYjF3uEqJ0qt5H91np2Gsdz0sudBVKkUImKi3ODvTZC//i
SQsoMpLV4oCC2U7rMkTvpOD3ptDGU0TtEkhL50blWGQ3t99E5kDLDh+8YpkQ2xOrtuKdj+vRZjSE
AkzEcJMMSrQARY9K8wn2ZYZiIatnSN1wzzvJSpZoLhPgTtf2usFjFof2IjClOpKVTo11jIQIkYjV
zXmJaCL9XvNYX6fNa8YcAI8R+pyrtG8v8AeU4+xfwEfs6F9wcr+k4gLpTmrldcZf5nr8lOpyUxbK
EM/pp0VIJE5rFj25BRcHA/deWP2aytj+MtenQfpOjlSMV2K8AlYWliGWl8fYMC51jhY4KhfMqfND
g44ufKXCwj0C28s9AdYrkEmDQDNFbf0bvLo3RQfxsXymI/5jQwJ/CmEQeSechFRhDDkrRVgwkf8t
tG6fPgsZ9oQ5+uDXuNI9danVlXJBRtps+zH7JO3inQzP3yCc/BKgYOBPiVvWF55tQqJeA39nU6nL
m+oJoj4WZu/AvaoidHiK+QGVpgWhLqhFdUFpMDRu6pRpHYd2MR5D9P1gPDO2X44t1JUHtEFx9un1
cDcBOhh+H++YNYXoEsvTfV/vtVPtTz8gL16dFebf+ti4NMfv0T4SFCmMob1EugSKGks6+SbqSx6G
5qI7ifQ/m82MLORIMp/HPxA13IoNo6fCoQTzKxeMwMtZSEqIW8JLVjwZktsAllvGlr/QsKOxVd3f
bpfc7ft5VRFc0+Iq4PFV0AiFkSUS3FVHDNTmZ5jvF/ZWKhEoDZqxLtDB+nXCh/e8E2nhY9HtjBXe
8yKEgsGceaov1E/QM2AeoQWmkhgPbVT1mMSYoBmbCCoBitlG0qCLtYQlKiT3PdMoPE6zQaawoHko
NNMYTTp/P0O7YtcGTmqxxl0kL8MntQcinDAt1nIeTDATdN9Gu1wMsh1bWMDf3d+nZggKo2RBbt8k
5bDU3YXVXcy3mg+aA75Qq2s9AcYtuSAGRT19nxoFLptmnMGwGnyeYlhdo8jQuiQoq8u4dRIJFESp
Pm0Nzhez+4WKdShsP7/pK+376W0LmwXflIXkPYA8hASFZ4ydyCoDCpfvnd9Q+qnEgYWJ7UQnzMuJ
9VyxjwRpvXfqwllCO7GMI9WHW8UUEOj80HZ6xev4HygkJXb2wI4ywHTIVWpjgvzJe6q+J8bG7IIB
iiI6PljHt2Bt0KJiQxVKf3pje+pLRZ51lLhlaLE2o5APsSqfhisXmJOBSP3jEQH1n7MmVDukAXOT
yAP0TTpz5hd9Ng27jxu9NV9hdov0A9Vp8acGMf+nr2t7spnuX1WUqktbURNnv9fhssN9x4Lvi3Fb
nbq3+P7R5qmp2eWw02/a0GGgYDxCPtj7p3/R69JXab5L3l0+ZDDuaXpppNifCAg5arXFpqnOua3d
8hiFHzZ5X88lacOoWE/rGyx+lLoymFD8BVmF8vAN3mzwv0Fk4AJ8Bz/FLuVSqpFA/Ctl3R2yyc2I
/xOKKFZ+jwmkeFfXgYYgzC6u/LtnaLg5wFSls4rdENWWvhTx7Ga/gwQ3abRXp7tuYSgBkAVJ+Tti
yOqXKAmlFrsLat/ye+HyZ2jiKspPile5QFlw/u/7UzzR1esHwAwqwpKU6SkjcJsI0K0r8jep+xsc
R+g3+Xt4tjN7owBDqPLwDcsCH1u26ULfURACyzjMBca2q5gd0vY5rLVDQEi2cOlYonZqnniDW0u9
06aNym7OcyQiBOW8HC3EFa1Eb66HXhg+B2+ajdBYeIkct+c7G76r4bnoHU/rkz7sA4tsoVXnjOvx
lfQ7qr4jwxzGQEJYyMd0VP9sqnfM589tGJUIuAWiZ56klEXGgIQ2g2DvoAkggqOyCxwsM+u4Y1yP
3+s+nhPVHfJopGRBfyUxGoxtJ7dw43WCR9FqIhwhvCXo/Bv71AysD64jHTbOIdlI1m5bnGGcZf1E
imb6o20K92VyBqUqG9LWJIM866NElPJum8TEl2kbWENbieGWEoB4b0jqHTUS1rQZI7Tg4bYaWM1t
JgkoEvIR/lG7XqO9CVVPUsspmdv7GBrJHttJ3UDgmVAk55J3tdUY0OdM/da+jec6uumXE7SyMfBI
k8RJklTKSHJdXPM52PBSsX4H5ipatsRow4Iw42xTKBaJaFJV3+icVUlVhqy4bViBQGiUyJKOt6qX
MRDo3YMoct+X7142ExoNzjPVjcmrDyIkiMRrqRl1+8EYHkMIWjoQf5EYsEgOq1cP0N6/jst17+nW
uWfCwYNxLUGXePbvo95xqJ8hGD7avRj2Ie5BEcWY5Bxd8eCNKjzWt2l5HRaFsB8fypA/XCFS2RxZ
/OHoFho5hzqDXCO7W42Z7n4OgHFL31O6u4OFScPx0uVaXeeYAkX9ahsZiLTRhL1+r355TjUjsBYv
SyWeEgPZYDLlDDpci34dL0vg4Rb75crQqHBbI8ja4JtXERMg1nl/5zNHrZsOXR3WGahbQyQXrkaz
e+Nrt46jP6hmy6Dvb5U7Nv69OICp1+F/CcEVhRW1DQVYX8TTs7qbfd1XXyZc6BkGR8nAavDk5J7r
7aevOHXA5V0yWlcnmm4ut5ZApvrFhMS88ckuMWrQdW4uHIhIUKLpAIJrx5blBPwqgbK938e1DK/E
+LlKnDLKUE8xK3V3poAzRNmngTq7v42uLyK8CrQVWr9825N2LivjF+UGMtTfKzIjTDSZCccGmv7V
0rPWpQkmuhz5aKSWzD0Yk8d4bOrGSWlrKJlDoslpKcKgXyzwOq/3yVq2FG/dM+t5L5K0GzC6Fa4l
GgNP1Ktf6F650n33mWN3wdbcxDbHWYikdMdbeakQIDZ3fQlQ3jU39dpMO8FJGm4bmG+ZSGD4eVg/
ZjuT8oWzDcQXz/Qb/dWcJgrUHtvcWWnDTUbmTzekB+kuK/42Ba0h1fJzadEddgF8he4eqZIm7ual
lLIrPLg0tK0AomJOIec38o+aPE/cGF1H4PYLc4aSEl2lIJW+BwIuT42tNwN7nNMoEuNL6OffwFfQ
iGUWeC1W6IOHSapAm8LUxVDp+s9EHXoQryPDTEjXIYTGTvUIOsgM2BfUC0yx6OB4P8fTESYjVWwU
2kKvnK6dia0b65vtrCzk92MHZVafzbcF/wF2KWUlBKE77WQZzl2TSnn6LvL4VGjySzAT1AVLeKtG
hZGULgwXP8JqBT7gqyGwaHpekbuJP48lKBCpvOxItXG3yzHxOZeGRuv+YkCNYKVogEcykiH3YeRU
BKV6NdFQ+5IfpoL2FUbHNEy615syEb1/ZBIaBhCOqyOGiagBlR/leoH83E9jcaHRCgMoVQBlK9u2
3BX+UkeVmTWXJG2vf2y3uKiRO6XSlhFKdyOfvY3r3Zbzk+fm6cr7X4/5WFFc/FOEuHqjQ1pcHr/v
CDq5qdQSBk3CJlIMNBsP5I4fwnwUTO21GKnpffXXZxCS1sDaV/fvCVnhj7JBlBC9hPuhM3TYyuLN
sMcnqc4t3cVpS+lXHQUEV39rq/ePi8nPbx523vHwW5qVo8oDxHJ5VDRzJrqd4cex5aAWtMb3QWIu
2eofRN6W5oCuc4q2HQYSHnYgIRXsfxrotAym8DC3LKfo4SozwX2A1yrVa/c8ampcKymeSg9V9fye
mgoVSrEU60uOeFWbSh9EMrjeKZjYIj20PfAVbNXmrUvjJRqvVPyWlgQ2zNSCEgKLxGR5hZ+V5dlK
8RWOxXQNa4BMEhaUEGHhLdxuHc+BIauo3LDqTk3xgYkqj5uBkSEMaB/ZAHqrZHEvG0+KXcqy7jQf
D9hvtmhIe9hl1pA/pJVokFs54sHrY6IhLO75tXq5RFWN8s+6WuH6wSfsw9DwsvFqsUZJblwJnklH
FzQBAFBv3wy4upF3xWrgdWFYpmXvCc8M628EjgshvFcdFYmMq2Dp5dcwMLi2XDgmbI+Dnbdf5oWv
lNOPkbI8MV41MAUBh/IcAcMXBRNr374UQWR6MzYPh2g+ObYChKXpR6goszSSV7kSpjNwn//YFRdK
WlF/1z+Y7KpoKIUj+5/mh6INdZgPVkd4VR88x27duQR3x7dvTNKAQXax/Ew7KlQmsE/habCEJEVd
MBAeuMokhzx5NeOQ4HPlKxqOgvtJdKw2XoWzizaARiHer5rQw7aZ+LfLUVjNgHlpJ7QWC1qNpUKB
ftNj+hyX8pmNigccQAclGp/46QmJJXB7DyuBuB2TNjsX7s4Q10CxRlf3Qa8dq8mR7jS02vy8e9am
T7tR+cJg9UTMRkaM3oeF+8a6UwEoml7+4o4vP9l4xc0W3zd6rbpl6s/xuQA049FRPoQlHzLgn2QP
+Jl6AzsWLmln94TlWHPOf6cJIhYLxzypQGEiikWf4TNhG3zC5ia3ac+YjwGiwQvUs3pYECzIE45y
QldaFxk8I6kqzc3w+QHfBfC2srDnnyqd1bCVpJphNDguWJ7DNc9dm4ps2pmuOUBAO0l7P0Q1VXa5
fK7hS6EjP+lpjWQP6H59Emn5a2m/V7XPp2CWnnyAKdgUHEuzFMQFbiyDvHMZZVYapMr3QJha9ckD
MDaBwujDgCSCLOTfMI4FqsIeUMAPCWK9+VoQSUJ8ln5YDKdVIuCmncFfSFCA+5drfEdF7GiLHc1E
LiOLk8LLM++paTijoZyB+/o9oBf22eoO2rCUn9U4JBKFJoXns7yYdETpLQ6gZyiLeL6a6NeGRUEQ
fFFFYpaacQSVArFCsMn/zZFvOzwMxh8mErBy18ZpOybq0kETynHKAQwUbMVnvf3GbOXi8DAUbrgN
+Opl60GhUhI+HRtVzRl2uSQUn6fNDIMph9slmtbyx6qxNO954NENBk3nUho3KCYkoZn5qDznweQV
3ZF1SD08n8Ng5muvTkZaT2WqzJKKl65MFIDoQpKQOvM/HNWOYJMwaGhaU+m0vcZdkyllJnhsyotB
H+gM7fYZOfvcp+HaVYvPkdgbQlN2F6NFFovNJTKcDPVDIwSDRP458g24oFB4TKNLHO1afN3aurAU
jwYJfAXDXlOFYXvhwsCAOG6F20BYsosIg0jVTIYBYTehlQZ4Qjb8yMT6s9bH3T0jfZyiIUHVowZd
vlJ5DcIADe+wCsaIoeRp4DYTtoKNlRNfZ180sxyl22YMWUd4AgS4XGLSeq0iVXxEChkDpiCN1IZT
4evdj7HmB0ModdE0VGUz5dsBM1VfLYXapCaf7u4+w/zE3z/UB4izh2GZR7r7srn5FhbUOLF4tES0
/h1TlBjlD5TbTlNcQkTvNxn781urhNRKa1gDYKM9+NEX9ClA5FmHhoQP+eWP+y9BZVkBrs3lJ4fN
nxjx4aCNy8S6Q6imEN/AsNARvrrSCyBlrY59DLfg5Q6Be6ZZLaCSWvhPDn+BjblkrdJY735MGpXw
Edvq7A2rnHWhrX4QKTaKkFAGpTG3xpBJBf53y/I6FGJ4B8xTJTADGJV9WGJnLiJHXALjU7Bj692Z
qNThl31EBp538LyciuKY+t0jU+YVIJiAMz9JNfJ6XNhed3x7x8TQJnKup14Balti3Q1D15+wjOK+
nyutJttW49QVGFvXKen+MzYcYqJ18TmzxpKJCfo29d3Ld171XLQRHZXYitolrCFBBYolJZFqqtD8
ypCwiIJU3Bo2Pm1RMd3VAVEJkMYLpqNZjcv1J614U8akadZMEcHcemwO+JyQold7LhWpgbdz/Pbz
/llljFOyiDhMbq2N6dYnt6BshC2SYhEpmGhk8LKAq8vKRlg5lB9ecpIT4iwCgaxLxNe1/SqgtIlu
Ot4b14IOTUJkhhy5fB/rcney3aoYbntA6BvcqSBWoCPb9hmof+fZdkIQ6+LV8umJCCEXNCFoaXGb
ab/IeR5sKPGSzD9qEhvHcbP14DRAU73B/4/7fY4ip8xGJbs9PZO0YRTnXk8UtJNkZ1y2jpswxiyh
lieO5l7Us51EoYV//pRKLaVzCKaHPt3huVJDH9f+nkTm1Kt51+MClI+MxvSg6clDajtHVCjJIH2B
Kt08S10SRi1kQF+tQTfrCjOFl6+2SU4jLiE85eivmp9zpJkYTXXdKmzQ0pGT1GFgQmKM4IXJX4SN
WKWHkitAKmmI/I6rfsgD8tYSMwKW6xYkQhXtmXqQ5hP4CjT5oOSb1uEuESR6e9uovgiv46Nk+2uV
PEUA/LPKet8V3R90b463Hj61KVM0F4EWvemIKYitgLOXITkVr+y+7q7PNAeJxBFVglWOxeIx/ir9
Pau0LWWZIU6lFzljclvXdDiSK4HSiolyfZGOUyVCGRk41LUFZLxCplDf6JJi8wWOXPPZEjlTqtkf
omqGskhB5qi2d/WlgTjv3i8Ua6RTQX0oxIEXkgqQOyOQU94wTWiYBIuJqih0MwZHUV2mq4eiD88m
ooKNra7Nj5gJMU/U2bB694hiCZpy51cM+1Jinb63wCUwCabXJqSsHs8AoDGlij6tCNYRX7mO7HrT
hWDjxkLlvXGOEEtg1Z0tgKwGR5pYSP1wAgZSLhjVRyuNwGSZB7LogXkcVKzejtVgWv5qvgaj5Xsk
IEM/ZXswCwGmEsAltV6yDtrgDK+fCIN5U2FE3/rvQXuT2Aj8QRlVGpMVQSV7aA/Z3wedHbTYk4K8
2HeUbkFaWgCkXpTGThuWnruZc8L/+JXq3SkalMTg2kiiLwdOB9nubJHtlsziVUjEjBk5wb6jqWHh
H9HDRLUOIle6dfirX6JtJzcGpDYQfDUIFMap7ZXa8bhBmOc4DNkgfsCU67p3lJuBhCRoyPBZz6Y5
hZDOAPG8FxoXLKo/dOfjl4QL/iOqr6d5K7kEvSD/shPHnA8LYU/V8HnAJ2ymuYtDu0Vi8VSuxIQ1
GpXr6mZ3qTN2+f4roYAWHIRgnCNSi5NV5n9YkXIDn+OlBOAo4lRRSMM/wdaCl7RossEL/iS+oHLl
KGpn3mkJceRjrlHTumnDcZyeE+UoJ5Gr9fLyuIAt7zQV6k79l8EtVMbq6SE1YDIb111CDICpP+ex
FFTIIQMG32kRSOVYZjLfKDmwmHyc+j6bZAnvgdlpFJ+IQALoYFGpRjpLZfP+krUBN4/zzW2NV+u9
uWvsUn85BbWJuRmIyGW2e2fd6ceHo+WPFIfSNuaKGWZ07wpCbMIpMsx36J+2tVNIIXvXI8kOgeYs
Po+Udd/cGWm4dV6dEJwG3oClG/8t+s4Z+fK3dOA+XLKDXxXNqKSB8UXz48V9nr4/YC8mMfbl3Ayc
jBITNHbc5oT0z/oQQgvbeDPO7cwTfygc2YAlTc/9MnORR98BuMgNQwsR4K4xG/bz05yp0CjdXnpe
zPFZRvIOGvz4O5sfo+jCIE9ZB08uDuOLT2PH2P1DBpXmn9TbMPF9YuurSFKKAK5OqtvcuYCofvwc
dJvJs6Qc6G/JTOdA3ngrRDdkfzYebTCELtyXLK0CHFTWCYaQ4pIhxT/je7/IgY0RpmUevngrEMot
N9jQ8lQ6BwI2nmUMj+rFNY/obiwz4SVG5UOstrOG2o+ja+rAxG5z6NakERq2WXfjVUGOl8NyoI6G
9fQqtus6ApRtXjmRPR35sXXP+Hw8Ltg3CBM9riOR4uqvAIkWRLrD934vdznGe+Sre/off4Tv5lMW
NHzKK1p80VVtAmposrbxqv12jKwSv+u5VAsmKonVRj2AOXv4WSL934M4vs67aIUgxge7HQTf9o1P
uHVkDNdex8/Ax8JIfMvafhFqmWbjoWc4SgClDXGLAbFNUs8ObAngpIrh0Xf8EaSTX/8GW5ZTMlQE
svz9GoJwcANpOWi23QTaHT9lvgDYJAEJqyybStrGQ2M8NOEtzY+Opj+EY29M/kvyYR/5dJY6p4Ka
VRGZZo8ThddIcwbbJuOJ1aZNnRzNos5OfLcMWUL458NavyagteBAWrF189mHOtzDPwuCb5Y4PwuO
iKBOL0WbDATzcwcxtjv0q2lyW3bXyYZnKDZIF5z5MKzTTZnhxSJ5zi2pIL/exSbcwjW3bNAQJbTa
hCSgdIZrdvpWVgGf24C3ENws7bjkjG6rar/+YKdDjJmhUupbpbw3Ug7f+MtDGn4hryHEsWLtcbKI
H8QBswPKXiZSpHMEfkX4Z10UefT0fEEf23dCnvN52fb6VewUCViTKnVDhr4b7aeoFbcoAhmm4ilI
pdwFq4Q7Zfh0OQX+wz5OfTzQAM208w1AFSYXomzCxyauXrsfV+0Il0mAEG04MivR8WEMUioU/17k
BcOEidZv91bxGY+0IoNPR5IvYgiEi3Xwe+QpOD9KFL6UXRwG/StxeT1m3Ol62DcgD2WDXRiJOn8V
qwh7vKQCWjYDT7MYNpNesRjs3UAdCxsUytZAfOijXAitMVxob06aSgt8Tpw6qM0Cj77faa/evWLS
s1rAVj/IgbT6Y9HUPAKeeSYjQwTI1bxDgEJqhc4RTF1je3WQG8s9QT9j4hcBFTkVtDNhY2ldD/A1
kjr1yvEOusdO3pzdDLFCfsIyeCPHiHdtRGExpR622gIcCWrB5UpsCbqoeFBaIIONwW3WytTyNNKc
JdOTpWsTtm9oEWpujbGQdACxqUGjnx2JhMc4esavL906Ooy9rwLxS8SZJvWnDoxlcKE9s3aaz/aJ
QYFhIWDrAEAlvuse7djAMQ2KX/OvGuPO3TFgvA6HVamPDManTFlHuB4C0JiETu843Bd4G+9SgJDL
m2YsMBYzug8ufKBFLEQS5TyS3deqq5VG5AfoeF/55lY7VHr1aunKUExLjw1OFSiNqhpLcVTdlY2M
3VF5qt/jrc/6gLaucNYMIhPSJiF9Z7P84C/iv7/FcWN+3FsCRWFFZPJXoZa12hVadjPHd5KJOZq6
i0jW3v/dLQOYx9Wkutj8U0n6DLVPJejW8B4KAfvFLTiaTuNFdajXg+4rD3/TLDRd/qgTqVZ/UHqD
f96gQ6KFq8Rywasd3zz83ZYu0inUx0IP/aR2xaAORNFjKb/jjBe0rNDmejIDn/m2ZSDOyT4UKLEN
qjmlHQ/ZZ0PttmKmh6I0CWoFMAUKMbhNI6sTAP5wIEzPzDGtoHyNfUIN2wZQG0a8nvdojCRf3oan
PY1QVpDichvW5q2lELO0teR9d4LNXcZdP1bVuovfPTWjsG1xLcERxx2QtNP2gOrqs3O7fLVwZwRL
eZ+ihXGA2FumpXObFHs5uaag1MSngdpgEX2mXByLNI1XnRwCGl6HT8XEPwVHB+gEe1gfc4J4c49U
rq6G5Fzx6y7Zz50wuPpXIFWnA0e4XgOJPL5yGq+5YszjPaT1Pz0APUvSIULRzGB5CHWBbuBWJRpc
+BbIa0n8NdrtcwyfOENj1ThCah+2HQkBGsQDXO55cUIrzxBzvshqhVf0EjAzowc2bDKVLIIutp9M
sXApXAH7unTF1K3nOQxVr4B+2PfJSDJKEAFG/iaPFebcqN2o82w2t486CxWYT+7HNbcjcRnJOJQz
9z/6PbepU8sSkYbDpcVUNn5MBPrdSXW18JcvFmsvKy5Z8mz7kMVZd/5wjRiNby4JURXI62Zypkzb
T6dXz0BI+91skfKGZjUZUjrnoVC2XSTgUaTgZ6AC/+ctSVHWDKjJAnYaNlveKbUj9ywQFwzxep2d
5kGbuktwbAaNxohcxLTYnKCMXZ00oNXd2/a63SVko3P67XNPZ1XmLHFn92nUZ8sozBhpetq3JH/f
K1Un8K7YPyEprNoLnjhG7OCugrfe6+4Kzo/a75sgZ6wGKJ06XcMlYelDHeBg3i77j8TTplJlRq8J
QHbI1zZvfsnrxdx3KraYRrrdDfkKTAPCPyuJtQTOnarudd9HTIk2GbBUYHEHD7oQmzmQI9dnQuSf
JUK41RExyK+MfRziArngqDlo9s/k6i/ZnaMXh43GT2yF8Ex8OwF3fS1sf9HxpQKKBxoYkzH2DCQV
EHmOdjuPL+Txotl7+IClg/KCZbi51vPfXD58tg1wRbxKZzELNsBISbv5icf3CtiUmCgcs4A/ahmm
4BK1kM9T9Hu+E2jLhXLK7gw8kTPYcWkVjUSR/ona7F2jIza1HUEhgf8Vmc2OlNZQe7fcPnIgLi3Y
dsCt/nqKWI4FlwNqzQ7XGwlgGqZ7fVkGVFB1ebqMAvPgOu4/JNiWKiRXfaAwZ5asPt8u/HTs4lmL
6qIXEU95DqUobXNHwM7dMtManyxDlLRNdO6N4qPf5h3yWtJ3Gu0SfNlcq7zrXtVjxWUPAEYeEf62
NoSMFP8u+7ptkfMLGyIX3Ps3T7boKO26h4MPlns86rYjVKZPxLCvuIjTF8r2X/nq7sWM8XKiVssT
ame8qaWPMXX2NZrEGny6e4wofgn2AqvdMiGm0J5CtjiCbeJ//oKqoY4Wo7u3ZvEXG3/pE8cFwOIY
nT/W82I4wXAP1+gWPXnK0K6aCqPjqakU6+Dgf+xa22k8sTjYKjHM5chCTa3obsqB8kWykDON0D8o
Wdz9b/u9y97Lwzlgamxw3HMp6LSok6rzyhUkAElo6cYlBKyQ9JGN8pludVbWtjkIfGck1B2rE+xu
Hizb2rxh52BXrUzuDbNHcNbPJ4/MDhXgYvDeUXNnJhPw5lhHDolErGq2YdgiKz0Lz/ajnd7hdo22
Kyf9moc6FuCU9n0SEAvXlYdgjF79ZXwR+oDGf/GAo9v+wVaOj9iEPRoZRNaASGwmhHiGPyXLLSyr
8NYApq3LN/EUituO3lolS7BWybSGqpVXxYi2qOv6hu4gPvafuyQ+OfLYmh+t0iViHaA46PUVyjiC
REKAwcx8RMCDo0sVLp2DvyCIp4tj95iif6GfGkigySGlg2xjdhqzTNCK5KmhjcGsAYUxdCVkDM92
ysPu4ihP25h/n3xXTYGLohdKx7n4sm5LV1i9vLcSZJWvhamhKPV6txMWeIs3Th2Xn5+YI1N9HzJr
i9xQo23eVWyEAivMh9l7fd3agGYLSOwXR5krBDxGmm1+GayoHBEv1DWRU31C2atEPv/9igYX0oMD
zcAmgi4NPV663at24jjv71RFjCscCBhb1nLkt4g+ef2Xhloe/tkTIepFcVHabo5EH9qcXGXjt7pU
d8KF4zrXX7JvLo5X+R3cZvcgup5lpyx1KKPJuxLkzcYART7u1T/EYlyG5TeHr7M6JwKrVuFpRTdB
vF17qkiHON6uJryYmQcMb/lPkg+3/g2ynzgC2IczN8GzypoFh2vgE+UFBsxm7tDOX451wlTfaNJe
lIPM9TYYrk20c3uPFpGeUrnRONWa9Mg5nqsrILx9ncU3zXuSCCOpKYsGeRzX6hp1jtdxqH/sjFBx
CuFXNiY2E0VWkOvv0L8HkzOV1X3MqQeyPz6ToKGyJwGAIZpROdMjLE8Pku6GAiqKLZ2LjXBorMwZ
bkIUXaUg5Qoa4J8sqtQ6C80qNvvn7FSKhXXK8V0Xwc1ApHJjral1HCBr4MfJlWyGYa93eYHgLd5g
jaTnL7eXu4sxVdximHwKXMS6kMJEdFIik6RqM6ADNFEsrKnFXgDBRdoK8z9f5wKXasQqQdnSQG4W
7qpZdGQSetDrqQ/D92DTCSDWlf5GANRJlcqJ7EcwThWPGjzKsaHbUWge/WX575osKVxO4BOWZxZQ
xjhFWCjuSsVkij369XMtHpKSVX2SfeNoFq3silNmBjP7r+Kwm7HLt5+Jr+t88o54lrjrgu+wR0/B
VNDA/rzP2EQi0pMbtJYpHdZlk/fa9/4LUylihzjd2sqlSUltanMhIF0JupNw3AkNQjR0qmwlM2Ro
4DPhW4+77IjMkme5SXD4R6o4h9FORYNzncJZ4kabwrqRIySWXkRUNvoFwd6getoMYNWIhgIZUEzO
b8M1JKFvxMDnxSqltTKYsVZPac2IVbkt9nDrpp618uc+OCM3UGdqOovYzeR20LOL2Cqszn2zPSmL
8YpUQGth8KdIuZU7MjPyfRGBM57G0vd6aBrCn86FivPGGySuWAL7sRP5OmXxvO9PSXdUQVgpYU1T
LtOEO0wAaC7gNdBCA42cp/9003rezpkMO9UIDE45rD+iXiaJiIb/xjrwAOsQZrP9Putk4lKqne2h
qZA0tjp8GhtYp21yfjfVmqI3u6oqW1mx2mVj3STnGlPUqlBaC9n1fBpL7wVhyJetkuMVWAMDdoWm
fzYcIxkaJn99U20QAYQgsoMRMNdMUcZxXwNi8kuUwF1I9eFoC2EvCa2xdYdQeHNocGtXlowKKOIw
oKBmbcwkDgUXUv2fDO+38zVpjqyqfEG5+/+bxA1dsKcknZiu7S7tl5osbxYNR5lKamVjkR/g6lpq
7kVYE/jMR2rtMdVWH4Gso3m4NK6JhdLXqtY2fVREATkvARZZIepK8CTeJxE0IpGAnIVjBaul8rFq
JkDutB9xoqiMuRGb4NUqhcGgyw3SMy0uvBa8wClAJfo8qMRv1K+TMtB5U9R7QE2YMyoDz2vY6Dj0
rozQiRDjWdDf12mL+PcOdEQ7EivoYa/lJc5e3ONFlTwGKgDWAK/iZRgu/SZenyrtvyvbuGwxPq23
GWOxDPzqrWcqXRQj3163nqqpeOccm9Bb0sZH2zmZHoqV6kJvwfowTrv/+p0clDZ3u1D0uxfwTYkA
WrkrkbuC3u/97x+LKIOdHAMgUomOV2wDJLCaUCacfxQaBq4GPatLwIAxCrZZiEq+zJ7OvcVztBC3
8w84CR6mtE1XSiYoQF9neVe/ilDkfuwANWkIe5H8yGlJyjSfqGn5joQAaMIFM3tFOiqtPrhZ2VCc
boPexs2boxkl1PDCnDdqL5dk4DoNw7xEEca/mc+hUUrxjwxH5ik25QltX3PW6gSEA3yNkHAMa4ae
iQV8dADd485wokP3KbApr96IaV6+BXgzzQ9JOayVrR+8pEJI/mGhKczoT9PKIWqNyCffAnj/qoNw
ege609z5J5f3O1JtUiZl2632kBpCyDwLYNrjIBJPCM7ojJ/xSAIi6/+tt1gRDgwJpPzwnpw2s37y
t5ktjNHm/H5UQ2Ai7Hq6oLkulP0fMMNasc+FPaVb/A0bCuOutLzPtzSZndcecI2ZFnP0QW/FlxIZ
3mudsEnqwGeg0rP5/zK5WsBF48ulft6ugslhhmSo9UcE+TyPyU3GaLIUJ8xHLD13wjFJ8qnSr2hX
dSZ7zNE0Gg0hbrwjvEFcLiySFoLTBXjhJkCysobXlG8iXIu7Hgigzro26rk7RSu7iIsIReBh+dQv
ZhU/Ch2NXjKISR2yCCxDkYsKJPz0E1r3Y7wVy+8K9H+vf9HP1pTyDrglbcPBW7kNwZpyTAS1JHwC
p3SPR02f6MJZx5EAcz9BxoOgQlnCJl18sWwez65CT9O+IDQXkeLyjUAKAuSIUNYrYSvlDSGY1YtM
HZaYS4566PhwxbfAlohdPuXDg+uL9ePUrCM5f8TDY/lyN059Xsa5i3di1VlICaZjWjog5Awr/jqc
l9be8Ulr17GKue2wj30k+Sm/TRU8psG5XgSFArjDs6WTf8XBg45zRMZONeOIUiZOCjIhA13t9IY+
TbiQRx6yffM3lEeEzGFUgwQAOiEg2H2ZBwjpFU3643NlQxzPeg75N+Wyd/O+A5IRcrbfwbciBIkN
LizZg6i5duF6SloaIk/5PPQyauX6baAf3IMDqYcJHASrE43q+Q3u6M14Bd5eJdaKIzj5aqnJub8w
oHmkBeql4frLoeh0ghYJcTueCGbvy/RE91BCx4yt7B5Up77YriBDAZwpzqCUIplOcdV/Gakz2IVI
wjFBt93kQ66UMEIJgT1u1PeEynO7a2hg21DunDz58jvrAB9bZSklwxoJz8a5mRA2sVhgT6epwdFE
SWEE7edhVSBgK4NAWOGQS8rD7SNSMSZdkOw3iWu3wEdjWyucthKN/JYjO9HioDpnxKo1HEixq8hJ
4iLPcgLu3Vi5YHaZ/UrJb4uoUfCyByX4xfX1DNONTcc+K0xsqxd/tWMN9PdLADY8FaYTH06XGgUC
3m5biTMhaogzjvRVGnSDCJGLP4FYuKK1JPuNZzXfiljkiA1hU1a5HkLHWmDtndXNjX9rsR+68sIo
GK1W3LmMk2mocMGiA1bfV2i47HKIXNvy/PSUblS6xyDOryy28WwQRRRgSxL17/olxQenR/Axehe1
ewSCVHuu8tLztqfWgF4InTdunQIql/14F6b/o/qSZGQWBF4F/ZJWhH8VO0FOhKr0rCgIW0LEEFsh
LLLkut+R2VrsRLWrvKUqfZO9mUE3JU4MShykN0yqh+VqgO6s65EC4GMI4HzJomhZ0WlAh2hwszDl
Ps18vPMOH4Itlotni1ouSFIYymfw9aHVE2700SVMv7k6GAl+FeW/wP+2UfW2yXmO3ywxceGmxzmi
BV/NgwhS2Dn7Cv5E0Zf4+iC09rrpU9eP0BiNs5TDqwMLc3GC/wUflOLZDsem/QGPm5dC+GrKZPal
MoCozYE2+FJd+7Kwj+XGvFpzSbppzUdPzZcxsTi6U53bTOX3xofqiJ8bjyuuxB0rVgsqy2ppkMKb
dbfjGh+glE6yqqxpZp54sLT+ruHrU2jGTliPjlHW+rJawx4XfzTFq/6KoXjgjUGt7mnLK5F5u/Cj
+C9KYUyIx5DBXxqYJ4bRWKtaQDlP0kfVrHOZPHQg05BPIiaIhGpxK4AOyJk4Nv8yn6Gq7q2qG1r5
KYOTDKaouCM3rEV25eWG/IcPKflxAnNe2MGvxl4utBfbOpMGVpbmI7nNFlXctwacEjcitaBy4I/S
RrmgSSVErg2sJqLwKmssssj6oJjwAAuh9IQOjOasF7UouHItyhCISopIOqgs6Te1Vu0aGGox7FlR
y+RDXkyOqB8xOzdB45mi7isU2iZm7U/nIuulSUFxhv9lIXQRZMG21OK+TbvEiWFYrW/1X8PWzwGa
GsH0kKBY6DALLzNywclx9EjcJCAw9bneyXbvrxFTIWF3YGTzmlwXANUDhDNbrKXAUkg9LLS94k58
VOpVNnHKHDqRrvy5kVelMosryI61SuNmvaQ6WeEI3KXx36oKapILoKU4XkFN8TakfliKbgw4gzsm
gHPMKpbD2vHJb0A1H3dOrEo6Hh40/8xemsMVdZUQ45PoQVApyJlFvITJpjCeis4vRG5n6KwNB9TI
H8aqcpk5i+coXK2NjHYunlK4RboCkRLEfdF7aF3R0BdZ0d9ZkZ76DJuo7nZTX0wlT9YjzdYQzOEx
txrDQeBGp3EKnCCmdZmCfI2euJcb+KKO9NqKEaD2j1kGHaXM+nlwetlzQAsvIcALVG+JLuxCvTxL
4rOQb0yVPIpumx+gmFz4c9Kc67ZbhXWpX+fT+eCRxFXrJ+3P8ZUzr+j7SqA3SqDsQAKifPBPfL7i
cV8NgDZ7mQYD67VKkQz+qKTxjj4xGqRIf3ckfky4oF82QStN84km2LyG4nfk8BGGubJnSshKwN/4
Lka1uL60EeWVtd0gmHcCP7kzLI4MmYEJvckWFVOU97L/Jyqhk6q/7D9Fki1jX9CCOzP9cJjXHy6s
9ps3jBnxzPiTPyJu/BojEpXFhmL91gR5SrSG3X1sZ5QIhuibGPacJYW7BX141PstZOITwfCmTt/I
V1Ozy58R7lukTVgY6CL8BG07GDqXOybIj1OZ0qAi6GjM8lY7Tey+LQWciHProHhc5/mEhwxs1cNT
J0Qpa8siHsFhOFd06WGDZ8gMP5ujwNxfm9KtLdK+XMXsxzNfR+Ke13SGNMJq8ys6J+4h3Hyhb5vm
hq5NvdT3Rfq94pYzFwIZg5WHtbxcyJwsqztZRCOphFrpJHh+O5lURUD5k5o0q1CVXdJjei5frFp+
piVACCOw5cmYYAyfp1x8Z+6DcQIHRXnuHjgnuz998GYPQBOgku2UXlB6WxSqwvuMfqbpTkkSUzTH
ybN5GPnRz6L6iDN257lmu3XdrpHloovszw2hC3tnDusdiBUOrBMBKj75ePTt8ICH7G0Vub+TLXC3
YrF618UWeO8ojLBhiebcprBmrd/FBOKFR3FVoB/rlre/kjQTzq+JDOJUYvulU4ExcnQuDjsB7z7q
5UziGxok84s9xFCt9CLkaeC4fKvgyjCQjxsW90FAGwe9pXJr8DZ0jSAcpvBWgL+WYyGUbJ0BaUre
h/AffIEPMsvLcLJBfVpenXhQ2SdjarWkxUsDsvIaY1BOf0QIjDSmwOijP28GoN220zqG187Lseeb
FKJBEx2kP4mcRh+gf3nQifXJ2RKPxo3jGH3hwqHII20tarlYGWFu4SS/0AI2dn10w4urzV4JFbq+
vPI5QDNWckTvalaDtjF+e17OeYrhqngDkF/l3CbPD3FXTYXmsdjOCU4lNsq5hVNpR+qKKa5dBaak
xp2HJxtBHdx6ZVyD7LQ105R6R7k2YC/uIu06EYZkTpHmnTYkoG0KYgA8BFSlo8m4Lr6+Wl0KuTJ4
L9eDuVzvpAZEvdtgqEp+4SwwsYn8mXOm0+uOWH4GnFniTd6AhztsAlseWu8PyvJATcFwbXRPhzMK
j2Z2tcOsspQjchFd9YHDgpEqxw+XCm/nACOELTLO2BUhBd8u3z59aCJdv9SL/j1QyRq5XZKrU59r
9ZCqaNxytlaeso97QHVAQGJPczagtgK3TOdM8+IJ1mMwLCWbm32NM+mpeNn4uiV9znQbAwAm38FF
9ec8bcHzUWrgwoAWQJT/iwbXnSDDlTati3cb7JILDOsNV1C1TmzkvT64QxjQ0SmHP6bQN4dxprt9
XBl6dkE83uF3IVWkR2LtTnr8FoOdrP2fpuOJdHjD/Ld/eRA9jMzL2pmwLv4xna4tSNxmpCYU4zS2
GQd1soGyhyp6/HydDCJC+0eHEF/ofF5SmjjkttAVgr39rZf5NO6YXmxMDvSBnGqGswNC6GZ3K/t9
PzziEQFniU6mdKmu8yYb1euRHk1hUW8UXXzje+LHoxwWUK1vV2MiMf8kUJP97pAdbbxK9LPqas52
Wr/CN7OCMskIEecDbD5Sn9BPg/voUtT1MOKEZum08kJetOEHrjoYV4RWI+UT0xaFiSGcwGlvW85F
DULYG2LfBQFJ8glglvU8ln6eoSFtRKEoowXv3r6w4hC1rY2Zo0jTHBVPhN80RkBpwbLZJr8tbFJ6
Gs7IBOL5W52FB9YkpZKZsqIQKRtnHyJau/bEPTGSdvNgistzH1NVZeYm3W04vw/ahON2bpaXgT/N
U3aw74TZ3fNi86zfAe60mv3WzTTQn8wIpy/vIOINtu5MfUDr6u3utlracatFGlpI6ypsh+SO4B+3
h1hLx8TWeb4GUwyxK+hSS+gL3MY3ubB/I8iYiU6m0TEvh+MiXw51AMy8zOznscR63dbPfvSkWQ73
rn75Bcw9xaXRg18gIPBfFtE05+ZSyiXcJGYv1WtqNibEO5ZkKtOb13vs7SZj78QDqIeQUr2LYgRU
PH5zic0xWi1z2wynn7y6116DbFoPI3PmA+Vf8cjUN0tmh/eAWuA08EvTICU1U912DDGrBprgeGv5
4GIXc69s2UkqpB1MO3MyOFkolGiKmNXXys3Xwbn/Q/dq9kQr9fe+cwUtJ0FecefJL38NKredBk6L
leG6CsOf8kyZ5uW9JQkFaxYDoocawUo4zpgRi1R2j9A0X/neKe98jhB9Pks1IKQnZF3kIl3zzC0b
VLLtdzthF+ExhwOn0Tiu7hX4lJgzw3A5G0oRo77IbGW7pmEOm4wx2C3JsWB6VnCSqrFDfdf1XV9Z
Qtivk32Ev6tnfd3EshplIrLgz4pamSXq4JaCui1WgFcECLdES+ryNt3TMj9n3wCJN4QA3+olxHc5
I9Sdr9PNwiJT08jKlhF5dA9hzfY7+52Awaz+ZX4lYz/cQiM2LN4X3Qu/NKdFLhKyt7tv8OPXDmCt
KyA8LLpwkNlCbeao3TsEZccCFDXqu8bgHhCiGLAeNrTK7TX/gsjoFH8OttDcz+8PG5QTtn3pblRA
HcP0qRhdd2l7Iqyd47oIXrLgkYxxBfKL7phS4y8Zd6D/KgHMwJ6bC+rA93JFGFU1kZ4vplbnzCe0
2pZkHnzHtBPHeTI6N7HnoXjgZezvFWJvvoNAbb2jwoXCbPdQHGgjuZYRjuy93Mxz8FTEb1UNZStu
Nh7Gv08E0Qp0bjsvcAsv1cyxxFTecky69M5JbwSL62khW/qBZ0kcanbp2IHHMKkWrrhUbyk9f0DQ
CT9RfQBj/arBCBvOWAhrleeH9SXpdIZVd3glNO+DeQi3+5+gldAHMB+FsFVjoCHSJYPdAvOQ56Zu
b54blVOVU/7OkncPOrwBTBgZ1jHR2zmSfxDX8TgUUPNBRR5Lc8F7/Cp/1WZAY1BxZrnwPInkKjL+
fdt5yL1ykXHPiEdS2gep5azQoOnnsf1/E9IpVER8yCTszWhAsD4QOEjQ9yM/6ndGu5qgieX63bvj
fPPNM0VpugTxI3y8R/zNuT890GFNk0idqW34erMoZlxPZbEKYkaVvVl0Z1Q1Zi4bucKbug7KQYJq
CixO0nQnaJK14ThpOutHi7VtZdfNN2UFq/kKmEWFh4c/KDV7cVJ58wy722YVHMZGmRiKKIzFcpIr
hfZT9bZBQ5HKdCdz0Gol0SvwFn4eJgJU4wO+l90DUIkXxufBQwXTB17amydAJG/+ShPT8gDHXC6h
+PouHqIGGBP+4XU7D7czMZ/Skpeza+GmMhnSmnHOpLCPbzyR/u4vytfcAJCBM4gHnMEp/cbYMLiE
057tFLOpPB2LK3xwm0pErXLuC6csNZd0bBUADxp0MuGYy7+bskKRVqMnhX4dffT9xWzTZ8z5x2if
dXEGY9BuIxs/hrO38OCMTDdhQ0+ATSogSADkIq1VwrAFjJO4aCf9jbwQODk9qmLYlJGjIaXexmIS
3nwVeZF5hzaH6ebRtwpLuw5Von7Yj8NNRWs+NupCNMBbXrGNsgANXEFvjqZNkLYGK6ZEEHyXKV8b
wrxapS81yNY5xQ4jmWn49WlGMPREOrKrpv47CnmV+9UdNK+dTp0/8LUp1Nsttp/LvQF2xNfnBpRw
K1+I3V2UA8GkrmCOiVCALVfJK1qpsuppAdkJ6/aYK5dye16lSG6GNenI7hChsV0f60m2Ye2kzyX8
kKDutvsLxnakpbISADpsasmQZdZH1VcVIxcR9br/mUVAYQZr+M3QAP4yCAs86B1HkJ/FSlBALP6E
aXyXoqAoMfukmijX7P4ae8cTQD1OAvB4/vtcaTEuKgY8iUahg9P05aP3+nnc0HDptvWqNDlZmLZ2
Gefk7lYgoLIoDhYw1k1yx8urEAbfy4rGU3eruceF1mkbRYiAFjDOGP2tdYt2RWIdJEYRykvtUYAh
9hlLBbpqUTlr0Zbus6ghJTHj7V4zYH/CgbEicmVy/T6DoelKtvCY8ctLaT7uHxOKVdJ9+BcsMUf3
tt3AjWM6yC/B7LvAfxt8yXp0vFiK0Bsam3jJjYkewKIjiRSRuHzROpcOdB4HiUb2fUOccokA16iz
iWX5Lj5AtPurciJM8OL/UrcKZAkg3AAV9coyv6sXGGbpBXbB9gFp4vCPm83A4KD7eWesu/opnpMs
LbiT0VReWq0N6wgxv035f37zBRO+1Q/1M5JqntOfmT67C3sNIYTusK1QZVIgOlEGFGbydUsTFw9M
DU46Q01f60TkqSqUm+ZE8oarEr9KIoIaIUYmxT5svj7sPqj7ddAt4RtNUew2raUcYltzNGJjSQ9A
lmxV6ud5v1/5pmjxc5fC3VHXhic9BzEg/fMUPAE613vfjVV8XtRqc6rQrNhdh1/np85Qyv1r3Dsy
C9vAfL9C216ac8oWbEbz8+fj5zc3BnVUTVaWPx7leXocUN8LhY9jwQ3Rwbu1C+RVvh3ia6ZVfE2U
+xjyqFnmHV3lddVpWBCpzqcPZguONowAL1/IhxJ77xzmJs/5ZZ3yaOmE1tVYXyfvfokySBUl96m1
8onZPqNKsC+GaZGaJ33uIyfqm2Jd1zALqEpcGXqNvHcQT60l7aN7Sl1SmQJhX1b/dz1xgOudHaY9
2UC9/KuyUatQ5Jz/Cf1bGLvIZEZv48f8obxh3coCpC3SCEZXbnjRnMKSdkdPVG8NIPDyv3A475cp
ncS6wRvsLC+6kEO5IeZ+fBbERz+kS1fgMGSiTu51DoXRDtKxaStSfYtDRGbf+p232uOCSrbE4XEr
zJvl1XmVsjGmTnPLb/m7eEP6Z59TDLPzcLwdi0+7azOPcsrlMDxA8AG4/JkSW1o2ozD7sdU9LjES
Py6g2JiWnQbATwWehjtdczDFbjV+Ski1x3LfKWVMetuIhNpB+9GADx29cGHplbS1Z30qqwJs8lwt
DXsCaqTtoZYkjdDAABXebWVeJae6aPHoXk8mdaiLA3Vvyo0WO+RzwGIkUMH2WnBdQLXAmvLXEJp0
r66jgnJgPi2pkuBme1tSfDQhgrQ5p767y8Cr82epOOqCbt0dyq053npxHQmlpBwYj5wDThuEFcYs
rf5PqnCEH42aP2RqTn9KAnIhZDfMcEVhlM7tDWTCB/UXDmaXrbWWsS8ZkzQjTrD7Y8GQ0FbMiYbX
nPz7I+VXAt9LozOk/uXP2i/WwxRBwXw7FvzlPX7l/ZzxtFjfuAllopLp5ftS8uUuRFhwM/H6nhuf
2VyxNx8BnrJNb7R4z0x9M+XZsWHi3P8QotPi/dUR9jSC7vQ2/J3tpDMpirD0E7JYDNWeHe49d5yE
Tfm7FMIFpzdr+1/ClaAa/JfQfFCF40HYi0K6knA4J5Y4jqKjarViOoLcJY/i/J/KoAMdisuvyRLn
j+hlFoHC6L2UuMw1cTHYZEo+8Ws2A9o/GSY60+sZjy+Rc0xXDWIVK04f9sEq7verps1vHlA3M74G
jtogDK+uBYb/bLkkObqGmJ34e8wN4FrwhrM9TlPJ3n5g/1Tp9qjnvxRAIFM8OheZd8lnarhaJvf8
hzx6t7VTVkZ0Yws5T3uITeCAYok0NC3Or960bNWxmqblsSK3ARXjT8CyWq17+QqfkA0cNPhKVX+y
sSh2HnFdbo6yk8mooPgIQaXqRUTNXh5T3W30cTUSXIWbyPBxcvMuHnFqecTfobOvmpKh/85wf1U8
VGXLDCME5HTxU1wYk4qbZG6fqK/DJle6/0OM8t2t3+M7bQwXhtlRuyAzA5/jqAPa953EH7VU8AAZ
CvGO7VzHCQhIAobeHRESwOznA8W0zQwxaf7uUcKILPyf1vpNxakXt8Q7z/eUg//ahcSkBgYx3TGD
Z7g6r41hrvDb2TkzCCau6oCNlp5i/SlB46m51tEICKp6fDipRw4g24eV1Cc2iU7FSDCre9JknqTn
yY2xz+Hpr1yIaUM3y1VBXBVe/s+o2OM4Du7lhplXJObOxYsn7qZ4HUzfBzoKZq2CJBBRAQK7m14i
u8vLuk4kK/2H8VVV93kLYCNrac9K6Md0hmyG0L5EMnv4+a7wkVHsfh0zUBozOZSD5fggZq/TeL6j
LvSTePlQ5pdK6Ndt2ILgOF0IowGF/+30T6SwfPSPUnKRkNoBghqwPVHG21ZaShk26wTLm4QGun5A
/La//IsvyKPG2DDwp/NslPrz8Jx8J/j18rYmLr9WBaC0tC0FI7zGGgWm6Me4hnN004+q3uflo/qe
xKTXnjHPDDucD7u7JOmknmBroIfvZR/1a55gsUuabY5mTo68lpvKBvpsPkI8R2M/Hy67EJQy8qpo
jl/egR3xA1L+kkJhj+qquZuOdGcVYZrQiYgtXGrcknH8fEqmld0giKcqjBwmL3HCWrgaiONoRzGr
HFEfl5OObsHVG2QVy7bAjllFLf63yBufLY6k2KtT5ieucthvNdbqDRi0FOEmOycGjH4EEz/JfVDT
Pp+xxSWe8hQ7d+klrxURDmgLXj5vGqIuBUTC3XPgNRyWXu594qGBbC0hA1O+WL3WR+d9nF08jdve
GJrl2CW9OSeh91v1sGYNaMNZLoDr/8MoYGawi/TXrNH2dEzl/VsVD9Y6K7XCoDiDu/0q4rNQ26oJ
4vpOgnvsJvt4LGpFSd0nFoLbAoeFfpho6Fjarxaw7uygtBF/KmpwtlugQvFcnuaQJm5W8tSKwN7v
04OzAjHQZ01dRirl1bdefLz9OltyXfnBDKSV35YynN5eCOS5hPQ3icUOAPAyGuMCWYNkyVfnHX+d
PdaPlk76i8TAoINeS5RK3NU8i0A6/lLZik5GO17VXBfklEOHB+SzZmt9fiU/UUF9qRdiTL0lMdyJ
/5utK/rxqKhpe8nzTnNTeselc89MLcZm0joci67goxmpafB+goa9wNwNHkq5YAD50iY7wUU1y+MC
N+5n9xd2AF0PBnvKI0+KuY/0Fd0GAgtdk34LIcAi7JIyBE0t35LDMTyoHN2HFswH40fO2BrmBOFs
oyvWqhXrP603x2+SaN9fsv2GWQV8P7Om5Gl4CFTsVGonfJBOUIBGclFJQ/kRWAn8zBVlb+YL5HxC
lu6/uZ06r01wd2LhqtQIUEMdrKy5aC6LB2dLbm5QzsRfvdFF7mBOxxUFBXbjaxYB1EAeK//2nCVW
YXl4Xkc+Bd9+Uu61qB1TcbubV6/mpQRmXyQKmJmwfzwLjwGbjQ46GpCsY8XMiMBVznCon5/lVjPk
zHM87UBtfMWtrUYg6805/j6pJ34fM8+AYHi8gZ/WhF4GM5Nj2U7EgSgQwBcovP4Sx0KMBnd2VAmC
E5QOYwS8S7TFnw/nwfacIo7Wx8Tdg7Yoog0iVRLt6GcxFaAotya0t5Pby5RsdIb8du6iiEddQHNU
qNAZRulq++IWj9FOHk8SG/Hyb+8e8jo0QtRtaJsx7JdPxVXeqemz1OGL954EqJknQWm2XSOfNaGN
abhRIgFPmWHRAtF+2aRL8naanQeZIYdRK0qKOepAUFUJoP0jXWUkx/IZ1jBUrimzQnYWL3wO+piu
9mDDO/o21xFXLl1Yh02kTcRcBlbZ02cc0AgTpJcKAeaynnO+BkwQhVJWZEaaau++F7ne+AZ9SMPm
24HlqgV+s48zynuPSxqGmFGh57F7Ti7F9IKagXTXZ1rBn1fEEdGeNeZ0ue42K8vWCDM7luRKmz9w
uMdHn3qe2x71k39kq3KxM7Fdszlbg5DUOnlLMlnPIslP2ElP9IattgyWqlAeOY8FK0QEOFTN+Yr9
cECC49hsTjc1uGIz4MF9xgLxZKNHwpDkS2ib3Xbwy+wVknBq/YOQCY8uq1b4iYCNHE9umKoUu//t
uef2RNGtAcedG3o5nP9Q2SL6BjupJxpYgxaNr5bx5VdBvi7jKTNMF432dgW1H8auBmCyslrtgVQ0
gKEA2UEhVM5JuSayIyb5BkGzX7tqjUdOLiD/nN4OrnihoZLVHFpxNTDR0N4Yp/97N/uHnPEfg4bR
lNgorjN0CsICRd2C8uc3F6zEXDd9zuKn3Ud/VTqCNSZguwWjBR69Ltwdtq0OI/2LbdBriZ9Oc7iP
4pm14cxlN+Oc2biuKV232C0GiqSn5xqWQTx9Y+oXh/So8fakSpKQJy0jW7rIRPqqYsrSs4MK4DQJ
dcGRxLlu4Z58Vz/t8zRIRa522VScbUipys+TAR0tqzVRxsUQKcTwifU9c77itfM8a8kayCdrxxwP
IziW8laorx9KzJhY2VnNibWmERGgIfOgwb3PwI/tfMw+drvFMQSH8ieUwRJvMjXLlXsLKtuh9b3B
K67PsQGv5mRpEEg6NHHDkFLbjg5wAzYrjGupJa05sf0G4tddUnx0OsxXqf9M3YeS9u+Et7STQWwJ
zuZAWvpzp4xqqG0/F1eiwMAf1xn82cVK7Ci2qmdCJOCrDn/oHXX1byx/BkgkZlZN4uoo2qG5RwXu
i1MS7wmGdO+UOKx3lA6NP7ziFAk43qxPxAEkoEzi130eckO9pfbejcz/JAtc1kJ6pPHUY2TEgMYK
Ox8Gq4UsoZQAhf/WzAz6swoCyWP4CL/XaCLbu9udYGTewfd+yXYyOkLHh31F3SuBaEOKKvyThqC2
fUclzRksOxZPdWE40Q+jeR5QGQ+lZqToJ7ass8dwph1/uxbBRbldf9h2q0NENWD4wFMzOSnTJN7M
fHqhk3/Sn+u0zO8IZWBGZw3hZlLOrv6SuecGkMkpMU585GvhYyugllgrqATF/VJdhNaQ4YczcX42
v9bhYqqTzH8s9ND6Uzu4qqOnOgyk113XMg9SnAPzeXDRAa0UIgVmMq+kyGTD9hB+6PUzEQFUmTqS
PHNFpvLVirZsz54Z/D7ChoBtIaM/p7tOFuW1Y3dT8SD7kqz4hbIOr6Cr8H9FWFy/48aHdW6jsMPP
dqZlyR1dzf74RkQTeRodKTZqzd+MIJ1MIqS9Wc8aX0hxsnVM0WDuxuYx6S7hD7yZFq2Tvkf5LWLh
r2GpT0Ct+R82e+AyG830EfMb/hcMjCEhaz1AVQATCHjlHUGFZ0MMIDhzyOSIvxUGIonaUleBeu1P
R4ldNy8txca/q9du1lUKkrOtXoYeVd3p0rEZ9Mb0bZxJ0mwz5uFq9qO2nDPRuraCbo5QdXWYLmlH
o5VdIc2d+tjB2GQ0lbn0GQdCBsTrH0UVP8dL0lQRPKGHVi4cUR5AbTYi2ZPGpLUR2vk883kKrYwC
mS0PEFgQrIofzmVpSZCmxYxwZBF9XvNtJHR52K0H/x1ah4to3/UX4d1M0/IeSryoAetEjnNs1vPj
GpZNXqlByob6+AR6yMki4IbIhGVsqfBMjhMOyM+z9FSKStVM+yGWhCRTb1QQcMPxj7DF8YhQamnv
qXTOKH34R6bHnuIuSL4i2jjQcjiE986lm3/USyZ3SNH82UXaER77ccXXCnXtShQwBckYiz0KTd4G
bc+E+zjVw2y6W+sph/4HrvKsE5dqQlB+Uo/12brWPRu+EwAmMndKm5kU0wxWPEgAoWQTXVibkVUk
cffEwrDcP0aN65cq8HBJjGzzW2kpN3EhdFf0hF9wAXqzttIV6A/sC9hTYWanrVxzn8Jp3HtqHLds
NPJDuZj/TdGCAKdsCuLr6b5w+qJso5e7HdnXZRvO8IPQL1CBGYL9rDmwxhyQwZhkSeoitolMI127
Ukv7QIhDYbEPpHLZ7EkIJ0YmXlGPv6J4uO+WuvhIPFT09xM3AoAa4JrP68yY3j6f38UtO7TCEuxj
AbsqAeOVQbleqbnsoDr1teaIoXCyK6+VLFHoP3p+d11CApNSGJh84eoHKEKCQ5VpWfHPvieYIw2q
LTKEKqivVAIDhgIzZN4C+Oil2wdSu/OWqL6SpmJoL/cdMmclUG20Ro9F4af+7tyWqU2Ei4mDJM+t
o4OsZNhJWixBguRtKxn2RaXQK5FsJo2mLWQy6yiq/YHI0LAncX4kWTX+0bnS2uhyjBVDBe+MNw4t
Mdfx8bFFC1ifJ7BGAsxMpbirsAIppN1unTjOny/3iSJm9KJJH+GXRdRSC8PEQtDQv/eBNigJ/4Mv
5CO5+G3ojAybjDAyMVR16ArMec5ZBtzbVbhDwLpCs0xIHvrL/vOcevxYKclkTN167Ol6/G4EEVI2
6ac3WpKG8IVwFEXTo6jfe6cmU6vzNN80RkUrPuPTuSuN/dz9+ox1S0v/2bCZzA7zR51QWH1n9rmU
PQ95y14rEWORsFm6UkiIR5FSbZsoEXnrp/yA/cV/+vPUKeu39Wa0GS2Rrh4BqWUfOGW+NAzGF6bj
bb8ZggQE4d2njkDqZg09DuSPd4TnueEmtuWhOO84DYyOQFzRgdP5SiUSo6iU4pudk8/JqvZVYs6C
14NT/1me2HZw9L2rnb7204or5PSKja4iXVuJfVLJCTExMUWdw0Jjj8rWDGd5fNnigfpJYoqacwyx
XGmYGCc5inzZvilFk7Q12t1t2Klt1whsBXY6kWT5I1kA0YUuDAhbL7/xyXHSea2HtlTNtCEbXoQ4
JU0wkXKI2S+/HmHwericRgfzZZUPC/5t+Y9Rmgu3ZuNeJafPbj/nWmYhk1hXO1+fwAcIdzAkDYsW
rbCZNf3OGfwKSJhgnwEA8iKZeBFapfXwNMPpxl3vXvzgrNvXIVBPmAuJeIzwdclElbXsnU/gw50D
bCkDmE4770DOgqJqZxHHiZeWNW9Hvrn19KRa0nShPDlIAlfNp6UUW5JnVAmftduSVCQcQ+QWjVK5
Lm9yu6wBI5G6st93TbT1JA5kQd/N0isYSE5pzraM3EJUdLDA8DGE+t5Wgxd72tqBCyy4geVyWCFe
X9X5tZCoCprjNu09lXVsQhJ3qIaPQty4ApgfEcrdEPxL4ESbWCqeW+s6rWzQh+o5XMyFF1qnyYHE
gCAXrLcRZBk74Gg5MTDxZ+DCwBcVZePmy2CFIOsQR28f0Hk4U+eB75vssvyCqVsgTT8AEZByXLqv
5fHRuYK/cfPDs1fAPTLZa6mTPSjXpKQZWTe+KVq8XcanRolMY+Jbh0ZeKGXaI2GYGV8bTv3/oTxL
NzhRmctvCSld9cowCmaxn9auMgwa8ML+pDAQIdCRd8kfFaDnFzOjaei4GOsxyDNfnpvgvk2fmHwR
PFOMwRq2AIipO/alsriTUMhkA2hyrqYG4Rk6E5JAQTjrowe8GSgLvx2XD3OPWg2n51lD1mLpuscJ
W85Mpjz7ThpoRDZRJzEjq7l5VxT+xotFH284d4/mWrKw1aUM5OrNdShPWwfKfowtw98LS5Q8GfNo
rzTjcyqfmAhVL/ETNmd7zRQrPVblMxHF9NdKqMQI+ghrw49Qs0uy9EhVuhfgNcuX7k1JUAYtE6uB
skOXjAUgsEWeHC42h2PalmnDwozd185mB9gMgTSwWt4cLRquZWlmlGcZPcWbtg+heYDRj1qr3MP/
eAkW7EHhEP7TpBcVSDiAnQX+pbViDjqDnwZBpkw0XnWs1h7HNpkjLArTwAR3RRdQ7A+QFLU0P4nt
Ze1+7mtcopyrR8gUjdZUOtZ5Uciy00JBHJ1VP98cd4Srd5xO52anoIaRfzYDEyioxjNK+TtvIUYe
7dh+7kIK/CIvsKLhW9bEfwL1xPNQBHasePsyEvGKQ0QUBS5IJIUUBi6ctnIzwNl1DmNk3sV+AWiQ
UCAvERJAZaV22RB9ovtbaCYUf77kYacVs9SKQE/TxGA4WYhrbH402EY7uA73XNK/ftx0e6iShxlO
DbKKF75hoTFxQ8cq9E3ub/VIeLM319Xy+NQ9wPt7V3mRpjFQRrjdScbL9sPwRva91xVfeYkxDV4R
+uFAnKmB5wc3Vd3oZpbMrwfLuvjlZSLfklS6tblKZIQVGDJBzOiYztPXsfJB/jE3BjyDIywDUgsJ
kHKcY+7XLfW3FdON3BaVs6tWoNz8dhA/Dk9J4EJK0H2wLQ4dSeGdMz6+WwIe8Xlaw749ZFI/J+8k
sTl1Veu3mZrmQLPSvokIfeatbbUpRgQztklmefyHnrxvP5svk9j/tWmV2qhryVh7Ud62hJes8OYk
di4l/gCWEkAzxBpOjASnTqEzbf6pAkJGDZcScHQzTA40ib/oQMMhWNMssiDaptJ5kih9UrYytJ58
3a7AAB7FFjwaRHA6dfJ9H1TUsYrQ/7vY7bySoZ+3edaNP2GH4F27NjRP0MRfPR4pyYEB730o1Pm9
ySTa6/mjy8nzZWt0bs/sjJpftrpCfGxnca2ET9JZopdWMUvkuZfr0dIxuyQHZMCAYiP2cX3T5oM+
BvsMqTagPe0Z3vaqf16LMnkVmuR7IBYI+Ynx0Ew69eW++ObRfq4RawtJ5GuJN114ASe7Zhwj5+iD
W7Iwzn57fq/I9Yp8H2YcmAM52tRBaYRxqVl9pmYHSIYA2fgBeUDYCJGFALX8wHr31djHtGcziziD
6AGysRuQpo/kAz1GwZtfCy3c+tfLqNMf3GIdwhwBpmSC6n3/ycMHyeLn19X8nr+2z/AFrCmlDc+A
4RtQaPNUEbEkpVRObzeiOrmfNYIxUo07U9WfB9s6OhGHLtqfNynzt4oF7B1ljhd4PDXG0QV+aWfX
n9EDbSTh4phpD+s6T/DQhCHtuK3F5/JPCucwsDmTEAIy9aqK2iUj0gMSJ1zizXC4P711ClrVft+0
3VxQCodfLgnzjEEnGZtjcgrOVVFwiKK0d9QR61D5Iac0oFE1QEGzUSR1d+R/c6RBd3YU5d7Rm7Qv
Fk3AaOp5EL3tNUWaiaQauHnwMbCLFI19bxAfd6aSv7s2eYBEor7Kdy9ExAGD8V5YXiYjLOolW5j6
hEozLL+A6PokojXht8NHzsXwHG9ABqw8rQspokv7capJTGRObkGSSvc92s5089u04rdTSivbxbIu
SkkoQLO1Mpbu4Mk7fvP3Q2WKVhPO0OMHwLpWz/TqyH3HY4Uj3rLzhtdG86+GKN6Spj1xIPbKZmgW
ZN3Hf/0EGQa0epjNhWoaygj6ExanGoQJPr9Z5zXpRJ2GzuALsO6AywsNvyP5tCp4w+BVmUJUBM3W
0vmvmu2w/v7JpjW4Pb1UBIENz0Q1f/WEiUi1hEfyfG/iC1n9PyTmPLHs6DM2iQxZNgexZFSf4cVO
sddMbY3p1Y8M7Hy++sDb1IjDtuxcq02Be7QvYuxfJm3xUHRWRR5oxSzn1Yz0Y1gtAvS0gue+opel
aMBrTnNjKlN9m1Y9Rqe3zaAox7FZC950US21hf25ujQbONCEQHWAsnm9pqKd81r0soN+qAHa/zZn
evXf5CzCWXvcJKAR6DPbWZsLPQ/O2ZUDQwJTB6AuwKccUy8Vny44ou+eCEvm0c067TbTRZjOqWgA
AYoOMnkjuvUwiviFQD8TCLC0xmEKT8usy3arYYdgXMDBKHG270PlPvrblbygd7jIUaBHcZ4ngmlC
DcXuWRR47JgUdH5SPefwu8FN+dwDh3OIfwhcev9t7qXxyfipMSJWCvQWylB5K31ytf1Ois6hodEx
+n4voj15uWaaa3BwCRWZnZmrGiwFEWjHX4sE/1rgXQmdlfg+ebanY+TWcXGNhfroItYOEjeHpmd+
+oEoESREFVOix8pIC/AN6ZOtZN0yqpfGYq2hxLKeKtfOXgYL7vTl5Ed5yPg6ptKIvctfy4igjcMJ
NgOv0MCUaDxKPreZduN+NpfgPwqZR2/4KJqpAqkL7X2n5wKYe9nPhKAt0MTFmPdLTvcpPIpcDa0z
mB5t+69u7K8xaF2UkNCx/DxzkeGnu4BbJ1+8sRK6FOvP3+hU5kycGtTpcJSB9KT1v5PMPhbIiTOt
eQM7xVGeaOtvxcdqO1DafktWA0iJ5idD+ax2Bu8sJQFI4z2x1UwjnnqF5OfvArzYsEAqYie0l32+
ORCaDJ+L6VFolmZypk1fZm7q+gq4AOWE/mFckGNWy3scRWYFGX319ZeLXH+xR9DlifSWIj+7IDmW
NrtAodEYyca2L+glr7kHfVnCSwDGCPVJhJco6NrlZJJ5czp8otbVBHeKLukJkpEiguXEFeQJAaqL
lca+pvKkNryfPKmber36BCcG05fSwqPTdS72oUK+4/qzmgNB+Sqbi+lzpMOlshJwO7GSLxbRqUE/
Rcm1FcWph+2V22AsVg7quwTnhFgepYpXCXiarugtchcX7GuKljFq+841f03EAq5njCucNlPE6Ac7
tU7KB9N6OHCaqxe/0I9GgNt59gaA27kNMz5RjJ2fxrE6Uj3+vJewTxHwtp/J0yAbS1wlWulTjZsI
NxT0ku4DDSCP9cv7BCD6+RYR3FaD50oMcs724sXeO8/qIrGFib2ZTuof/UKmE4idz/6Kd7VQKXKg
cKqsdir8sMpQ+oDTWBmQsK8oLFhevMwJxeaj/Cxyq7Tjv4NZTZvh7lQ4QNhehif2Ki7hQO/Mprh8
WKWgNeIziMBHc/1DeIiW8xFCrZkSDi/0LcN36wazNhkS8jGagyzQbSsY2Bd9FEezpKr1pVX4Qocx
UZFdhTkAGoBnHiGI9bqyZpT0NxdgfCTnwymjr2UX/98/SZ1Cnum6u2J67f9s8x338OymyU0RE/To
8hFmC6tobCcVfy/IBkPovB09RcG8JGPCS4P2avsxZoQl2i8TM1HILlqnz2f3J7y/FsIqL7Uza83b
qkpkkJ6AgbgadBH4tQuiOYAzSEH/KgmWArPFkDyf54Orm2boDbg54lkRfpA845Tm4T7MnpoR88pw
JXPI32sIJqLnrvXd0EvJkApaVIOxuqIEINmC2xv1awFaCHOkO7aVqWCLQqXAMn1H2uRPkqm23+mp
lbwTNANPbmnoMBQZyAw9Hr3wemBM8qWiCNkwvLOXCQf8LEjckd3D+sQPAJljRz8xFKZylVSm/TiQ
eARPOYIqCOjLOtoRXR2U9yvsbmry4mKLuWq+HgvesflWDXLiCttnQlxs3s69NprcoDKUoxYUZibZ
VOQUw9VT65PCXF1hmBb42hS9vw5By+N7u6huR2DnGMplwfLlNhXiI+N70BWSR+yWL0e/LTpJstOm
WNQcyXYDjiIi1k+ryDtm4SQnh+Mp73DJYI1o5QatDowr7sEaXkFwwk13WlPjSakdLuxEFQ0vN/iW
Kww8uGu95m8KhNrKJXj52oHmdvVcI38eclXrPSQYS2Z1lNII6IrK6Ygk/kEx5bHecAwqPG40BEVS
Heap7cu6y5oaPj2kqYPi48BSFviXhBjJ6oU7VgQUBfMpizRP3MdQ+u+U/tZCB3TYGKkFzH9sfYZs
xhIvsJDGK5Q52j4YMRnPOCQtaZ10Buur2FkO1zFz/kqg8sn6/4Myj2p+wsjs2jcpXq4UHpQh/Dgf
axrTKE7aUXY4PvKwIG61xh3nhPi9o9dUjQ/yQLRJzVVCevJn/G+5RjQZXC+YNeZilT4U5wWlg7ug
VB3JGnTJI0wpXhwc2E6gdsbkVzY2p/ZeEcTpBEbwzsaVNFMUDxDWrRfSbRCf3PqGub+1p4hWjfXk
n4xNxCuokw8nE8rcWzOoLXwkzGBLKKwLeCSeE8ptpbjDEH+i7X8IQT/aDY/0dM7PwqVtzB+swbyU
0nrwJZMAWfkKvMLkCu3T76uGWcYJpAdx2iakd4aFytU3xckevZFK1KlAcwpNwt+A4MYaaomGrvU7
WwAcdsqlPU4W1jiCSqvwczkDOeulG6CTk6+/GEgP+NUKzL4YTzbHc9bgI66TAWQZTNqssMVXtB99
ARnY85Pp5y3MzMNXPnPdQgm6JecaPZVxvc6e5LKdQaz1Cd4+5wuo3+5qU3NwsZtErRxJEsskMldy
Yaz1sFN4VYxtYCaiI7juKU0tk1FPg4hJ4onq3nc1VsB5/sr6t01/ISLmybHh0wXMCxzw9dtMiYPi
nkKiYE8bscYtbs3DxLNAv/BKiPs2enemWVk21TvP3SN9+PlD8y0gOy7rktp5IKTMcXnyV5peYVQ7
JUPc/iigT1M7AY+ZeQ0ib4iS272w05NvhIU7KHK0M86oxtTjqSRmVPzI5x7wDX7TW8/XdQ+dZItz
NTP1AqxKQD0APJ5W8bJ888JTUISZaXaZXvkN6DNhHNLsSGp90WWRnS9QeB3rIddATu84F1e2cKsB
M3PdZ6LGmVSPxSTihmZE1h5O8NnbwU6EjCyB4Rh5xNkVHWTJ27DHdDwraVfGm9KGCwllbGPFXmUY
ZNZ3Ltg0zydyQ7mfUPdseK2c2JSGFX6c9kyQTO8nJlQxwMCY1elG6Y0RNGOMIfGePTvnqgtpmmEU
SLFE17nqxmTycI8yoxnXJd0Q2WezoJybbYfcUO2vYW7Na/jqU7SLsrjUCTNSH7ci1BRqD7xE1Ykx
XnZQ5lR/pNJA0IILmAP5ty+fOcWrz9ep81ALDdPZsIEkn1Y3kZ1b1uJ1qZoOngW4oVFDLvQkgB1d
E6AOWJY4fygPumyTzfbzPLNZuZrC/b8JtTkM/LmFXitzczdL7FrahTZSumts3ysjb5iFVX+rPDmi
4eiYOVnSAV3wsA1Dv2R6lRZsyiQc085tuUDnN8xnHOr27+7tZ5j9yg1OUVbqfP4lWhCSMy6JchkO
9P0taknEgiPXLTYVKP10x31t625zG7rIYHwORxridzcaUPxmbldTsmL7pc7dpaNPiaOdItiXx/gP
MyJSYp4lnr/MzEgrjuMEDtvgaaEm9xp0U31oufyNazdB1+NaasY9GZEZjvPrwfF33GnoHaYsjyaM
wA5RRIrpGKXDIVUuO36iwSJ2kuXGGOV3Vcu17lucsGEmjubOUSMo+ZO3yoy6ZiEpsOxwNs/U59YM
Qer0H2D1jpxGzujZxRSvT0xoZa9dxPaxfBZiGFIUJLzbY7gbtIXgHvFjtQyrlCqJSoCGRrcbb0Jj
UulBKlL9bEtcQxbNavxyN9vr871vkMTpYXdScrAGd9FUAnnE7zc5wfGoXUnUaMEHjonzYw7PKw9c
huhR7HV5dCL6AglhYgy4273b15RLH3sYDrMjLqInemyfCcW5AtyZzUgKVV1F/qLYf0GzHD5a9d8S
V6l1Co63c0MHUXayv6i/NxKZ7pdOh5ABN+PUvkHDHSNNQmvOGDr0uakDgdhLWlZwAY/qTlnFR8/z
Ag/fGOpVvV8ptAHjkNsHsUwsjgb5ns0rCZdzANJj5I1D8YhJ4mOEOVyp7lKzkGFWVMgwnDvyKbeG
3Q6wvtzCvKfVAtQb6KFsGdnubCXFhouLn5oWF/rCtlxCGc0L59CUQWeDuwI2hdFkmnBGB83QvQ9h
HxWMTbFO/l6bsv9DKpHp77dsZ93cQWvd8xz8jMSnSAzX1M2zjWw5nxxYLHjFFLtZV1HJSX81ro8S
r27DRPCfyBU0su6BcDO/QtjfidC1Hzyh5R0okg/N2ylRYRwo0zGMfCxzC/zBfpn/leBhjwmkr6wv
VGL10AdcTskzs79k0O48nxL4y2e/J9R5roQZplG8yAJsKX3asTaw1QugAZdMy5WAa7t4VvurLt9f
8hi8ylKm/OwHCzModcfGqERDc4FhmUkJSE5SpEBwo5tfsYSJ0YNznsBv6nf1zRdUdZv7uYc0Zkr1
6wloF2HpmFZGtAOEObE6SLf1iw92AixqWbv/tssmBHexYQc6a2f7/jpjiQIwjcs/sBwv4KcP4y7v
Ee/zgDPII51ws4uj0QoGc7Fau3Ww1/KgBFHqnt34kQ1zQk+X3oW6ZoOQ3Gjy58xG5RFRFz5LgISU
18Rf8FGPCOpeyWSmZzvY25NGJ8Wu5p+5KyhtyuCUY7bgkKjipQIX0pfK6gaptVPobBa9jfcbX8cX
zZS42/hJcK94vpL2YFCVbyDEjvnBhU068LpVyox8LRFRz2m6lKNQoFHiAqXdhOwDwei+kr+4hu4D
tAJ1lQlV9Ro+sdyxSvv2W0iw1ce60Oqn8rwz6TCEcznLckzMsEP4vti1XHet0IKWtcordOZNPYwT
jpGAxTjquDvSrcnoAfIAeQkHSI0xEqsUar8ZKCfAEI/huPy+4dPO1tZAyOjGrPqlTSoxB3H/wXGF
opCI2d/xqKf65/Oe8QizX54TzIUXVxQqI838kPlKW3YLM47kxALcp46QEUqUHwK5ODxGkremMLDN
0wERXjSIY4J67yyXmfZ/tdOTnFJMNSPBnxubzgjFvIK5j1Pnw6Gw34m3WUmU7pexRZ86d6p/JpOv
1M+dGXVjJSTkWRFR1MgVy763Jdr3RVcwdMn9Qios0niOuVlEplHH0YBkgv7+V0vkW1YY7zy1G1rl
FR14yys0Sp/3gk+DOuxv5koPqvGmztzoGTj53XSAkF/jzqTBK0hvecJxYtasWhX62SbOg1EPKG9U
HBnyw149t9qczeHZo5EyETUNPps/3Q42bopLvVlZihLMDY0uihizV1tW/q4i9dacJfLa+7UQ2N/I
r6PAqxG8ZdxNSyPqHzyycPqec2R+WH/0pCVwD4ApEv6eWOxLYG/EHlYBkg+lNDcK+d6ZRSIJEiB6
No4+uhSs33c2DRDMzo5/U73aXrAr3TX5vHK5AhdFIIJa62pi73QGw7VBd9D1KIRvd5FMjAox+EAV
U8iln3QpeodJ9bQfa0nPBAFE53WlG6Cxo3l/NT3zSj9eEcwEsT6MeekVi9qeYNUFrNPB6URwbHsj
nLsXiAKeoGoCuFwjEIQyucngMSmbgQoPBoaNfC49qSZQYnQtITTOKJAHF2hQkeWd0oXpg5MUfnEv
xao9V2H4K0s8E9CSs6Arf187JgQkPP+e6xgHaI/iP6/N+GB1+fkDM+Ub4g9q4jvNVdSwGivXhapt
LiLsYq3jUTB7bvJUBeYCLfLMr6ewIN4Lq110zi8o6K/wm33J1o+zu6lYm4uqULZOQwI02r37hhcS
hoDPoN7gdefq6u2/80hzPybOjy/jHmnWXts3kSbtcO14Hx4PkFEtkTXrKVTIG6jSo/EJ2V/EOwya
Q7F1TFlzpmSGT2n8q2Sod54uif0jTcojgU6JRcFLY+7+rnq0eDyBqCmoN13mTb5GzeB6YV6/HDpv
OHIbGUwq84pf7FiJzEX7NNtoYIgm3MBe44kNdikaTksi+oOdGLE7pqcHjo5XhN5ctSUQIOy8whbK
/OIraVLiqrTVgPX8tpr66f+k9u2gKTX2IvdaVaFE17gyogTQOos/IFCCYRHz0tziXu++o00W4mCA
u/xKQ5e3uyolQCFl0BNOBHqJNJ3RDDy5Ahu7D9tPSI1EgJUV5SmDH9hbTzPJHnRFEzQvVuFYuCuF
TNd3K6UFAA9miQp+LWws6ifvTjn2cvsxekEs/zdKGhcYt47DN+Ml4I3fPYmNs0B6npcYGS01hiZB
q92/t21BiS0HzMwd3BKtLSVQsHf9T33JzB3cbz5F9DytNU54BrYPkwn9uAZxswdWr8MBidMwjCU5
K+jE1no1JJG3LjnXVoIv+AXx9F8Ov5QI1lUtbbOXQZRudtsp4Gj9x1a+vN2dkkGH4OFcbsXSIJv3
Z9iWmGTl9rZchkaeffJKLt6rNQK0IB2YEXLKxp/wTq528CHClqDJ1ZdW7qKEWobn6ad6h/q55Yk7
ryyxZ04/JZ+XqveJvk6rU1GxwEAW5UJhL8iumgNwdQaS54JfsccEL1rWdcQnyT6yjCBLEoUPel7s
Oncr9krvHEFsGe6kow29/UY0ikMrXPIOeN0X+hAJfZxteKkmZcqQ4YnvVHDZSRG71ys4u3F+oo8Q
swnABiqkRgvhri6gTN/guO3Oq9lnq/DftHmVOB4YZJl69oEboZJKGUW5HySRx0nEAqMxLeXazThV
N2T1J3l8+uynT7xOd8SN6W1FPG4I0wBofRWnc+ZNpCS+DNEtqm9X8wJqzl/k0VivygRjm1XMIqC2
bAm2ApBPGQEv9Lp41KmOn615a1HUjqpm4iGCM7RTCONdo9cBKgI3sgMeU06inHUr7+ezz5TR2Al7
ANkzBnsHF/mQtmROUTUk8J820EVptPoIXDqDgMdklvqwSPIYmDB8m9+gCjgQh/10m8IIpN2G3+Ap
3g6xPIlKRwC2ovkNW2C2NFHRKfJOUwgZC10q8FHOsygTJ5Abkl3FnnGzJGRjDbmT5TK3y5vYYS1R
i5kLMEbT2WVyHRAXWqCI41CrmDTxvwTGLsf2HR6+UYuUvR+cWliVpI8iyAI3Enk2lTPIYconPh3b
NLvQpuONWewp1SKL4DRkqdesOZvRO0GNhrCESHT37Bl5PkvKJJWiwBWH4Dk1mRHK6F2n5C7V5bU3
fzcu8TPMLa6SSLz+TjflVNXjxL08Fb+WjYKDEhAwCYXDFNFj/fDRA4CMOAWNPI2UICGAQhfikd7l
hj56gQhMMYN+6/IbgBOG7KFPpqNa40Tayy5u81ZIhFn289IcCISu/Kh10oJqToAOvokWB/qxcUs9
wpupbuAH2DqpO1Xhe0GIVsuqB33xU1XnEc2iLrdYC5A3fJLfbIa0mzRbsDx2lZTN2KjOVDHMsJpZ
Yf0GHCHToXzkwum3OJ6u+rET0Y7DxVIzLgC2SSF1phZsFC8/onTVT9uKUb+fr1eztHmHR6vRzEdn
VVjph6kc5GSEFkp1yp/R9iWLGrNoLxrFONYnuTtULWO1IZgmNY19GEPN6r0s7qxfQzBY7taXnpVO
HRgXSMjwRy1/Zof7IkKWWcZM9PLtnE3usgxnxmB4ELkkPinQ8iA8+uExtbXZb9E8oO16YwlS80vX
tDhIuuzKUsH5ThDw7Bi4L+sKseT7dvwtm+FdPWI9H//rZz62c345ImwqVsgqxWTtz94yWaAWZIrd
sL+gtxsg6HtCaS3nVQ61c7K3rFNp3IBdrTRZfBwgoKlOumsW7fR8tmEkxV4SNonfFQ9vYITw9M8J
2+2MbDplGHASEoAA6i8UmqsAKMU2OaVB4BVvjIpJ0jvBKZzHudrN6OuYwfP4dj8xKpxX40LpfpQU
gmtEdI0mylIVTZQuF2uHtIIFD+Hz0XMZtMLrX1BX3dKg/1oejMErTah40pKWZkAMColSPs9PFrEp
G6T4mgrsVyEdsTJp4ns9hXTvqcY8DyDwOfQ3UvK+qIL+ZBD/HXNzdsi1uEMaR6V3Z2lTSi4ewRVL
4dupr0/bzeZOIPM/5FvTy0VE3bXO7FEBerybMOtyknReW8p9nOXdbTUnkTBAzNBeCfgRb56Gpf05
WPEiWNlXHOIXnHqeTOx9rhF0QpXRRL/Ww4ivWR2/ZhR7Xr9CKw4U+Q7cvlzaOl4rLY/SS1eGk8ZG
zUGBcCS2UfU8aWrb62opy1SxTuZ2oD/mGS758saYExPRaN7Lp3XOTwRWXrA3sqy+e7d8Y5EA1iHv
vx5OdWDJcdh3sO4onvmk9OfjXq6WXObGxYeEj9jpsWuVo02txO3/Sb/e3rFugaOdhylZ7WHsxqGJ
67XmTwHaNYKBz/HuYpoV4ee5Zo+goripGPYSDwvHxvSbu9gHRRovN0J3bJhLHMnRlWsPwUNctTKE
h/AtVQqowoR9ZGjjlb58wpI5PcVsl0bbBfof1m+Ev4tYxxunZczgB4ELrgbM8cpO94e9Dm1hP4cG
vl4XZ5D6LDcQTLE1+Mvp/F1kqYOqQNrihG6M3B1jMFwVZtQ93D3ha0DqUvlb9WAhJTKFKVGsuWfV
NKRIptc0XZ/d2UoVrwH+OXxGV9esGk1Exs1zb/S2okD520FlUDSLlJxwZj288C70VSNm4+28WUxd
7CkA4RUuoR2MbI7wi60CL4KTOKimxEigzXiEw160C38S0KRvSqBqyhI7rrHnaMmf1xTJjNPVGBlk
l0ozSCOOSNBmWQxYg9NE3VpQcV2wp+K94JwQW8B/O4CDUvJ4J/T2X95tUIapr7nzO8Q8mllAyEZV
bET13VoSu8lAslFlazQSZ49CGiC+VpI134qqslo9tu0mZzbwSWpYVN7/gBWyZYlDMRaZTPb8UPQ8
j8JW/5loQ4T3hY2Y7XoTfCN8fxZz/0PJ0k3CiLk4dKfbp5d/5Uzsn2au6niJZAmf0YNr5r1JPkb+
8PR3XcxwlvNjEU7PxwjIccOHuKgtWX+granwjNQS0IbmM/zwKVQ5pmcgnoBGZYjTqbx63IMK7mD0
rmvAU4IcgTLvGtmaPgTBj5oSEgVfmdv/OqJqwICNq4ph5MtMRfhCFPVOLaOJzMrLiYX1ibju3N0E
ZnFcQ7LxEgnUThejqvaxHaCVOzZv7g2hVinzhfEZsH76wJiY/QzupdNVp2/j7Ll40XRMaFpfKoT2
ySid02/6+n42jLkUBVr1XIT/ntsImeZZ2RbSz2kgyhIskumuaqn8R+4JQl+D0MXXftvkdEqd48Yu
yBPIo2MN/rXDE72m8FH/USRyyF9HVoJK6JP0Cr+9r0tAWEoAzd0ZAT2VadkzLkfASOkWx7UfW9gg
23j+jw3USqxCacN4Ih02q1hAyMliyowCTJcQgivTC47G8fAalIpbJvAwEW4anwlhOBLzaoVQckN8
X6WbY/Gjphs54EhY0pB9oT8cA3HtdbIf/C8WYQiWwV/Ob/57Nh6phRmtIFmm98Dzso8LLkEQw7ut
+ix8FZdL2mCs6dfA28nZjpkx/a1rVN9KwEiits2ifaTQnxDBVYB/0Sxn9DL4JD7W+WJOc4M6HWJk
vlfA5ExUWvpWqD8JYond+/yYYdKTuXSUF5I4xqwCRyeRVDzmVhEg9osZQu7hW7Rykqhln8vEh9t6
bC4pLOtQI77oshP4EShBC/Ouc0yyXuwy2huXfHxppx4QeUP2sEkt1c0n3jIyfAtaZPbgXmM3VDHq
BU/DRn3CSAdfB9RjOU2RFXVjhxMEonxam0Bh3YlNitdoUF1+pN+Q2yMt/dM3Q8+tNdEJ0hORrZcI
v0HajZ35JpVHlceT/zb9UvF3UFs6BCUbFvfQgRrTi5Sp5p0Vi1mF5B0PqenmkCUf1I8ukDV6jaNi
I8mtvqz4zWmRrIMRm18oK0GLqXQwU+kOq1Ic19XJWEYzX95jahDXf0gzOIRKzTNrISqhIpd3RO7H
FZ6S/tJcht5XQDL3k80tI5ahL27Hwdh7aTTMc8yF+YhxDkw2WK1W3IDvXNR8n5k5/14NnrBO+QnD
RuXUwzTovkgdEk8sgO1lftLu4au/keX4hmT5Wlijx/EDCZK71vcqfG8puhDJslxrTjT2hAfY50wE
+k/NxT+cLJV4KvlO78qVldLNC8ghRGYka7YNmPJByOYBGHyA8/wTUsTf2kOtss8yhjyy0Ry8qbMk
UrVPpNBZxJ/wHYxdwYfI7DkXkSSC6cuL6bD4YLxwlJjr+SwI4Gi1yjy4tZHXS7hG9uoL5KeqHoH2
Uz1QLLWuQ0v2LhuE5FoFGKU60Gf4pnV50WtT6g+pOFXpve+NiFQ69ynZDhz1wCP3euCqW3pfJMuA
bV0/nJpjJwFtdgyYonbjV0uzae/YQHrdGNhy7RGsmuhNdx395q8MzAB4/vgBlktQYngJ/A22dU0j
EjmojburWyjT24NJYaTu1MHzXh6V9j94KuKE/jFfChr/0rZFiGAci38+6mvJMZ5VUQ2UQQ9fJXR+
UZED7NmOOi5c/e9G7ckkF9R/JGKu5NIrrFcmcJthFD19LYw6d4ChoOUrUjrfFX/0xCLXIy0F7mJh
6CD51WqygE5HA7sADHYfWBFKzxLRALbS7/L7aZXpYokw6FqvEnRoOlM3FUzJTs2pW/QDydhvIIGk
VUs8wghN5tp4h+1mQJHc02dTiwCv+bsrrbiRowsk1xA6maZI1KrxTQw3cNhptFLishrsXvt1rbop
aACDUDxXFQwuCav9mk4WH15JxBwK9DgdNdsNA6v/aVW+URaHkAPm3o4Swz3tdWlNFw6iClCqg74S
f3YwMNHfxXw9WWY/3CMqrcbgwvWxO45q5wmME2hGmhR87FWPt2jnbE6MVgeVzOuZ/rO5PTbUXE5P
uSH6XLvOoPpG276CNgUkQq0rwhzwNqkTlFsa7Z2sfuTrwzN9bBsK+Cklw/lIWfSTC1W/CbhWgUkO
hy//QI5K1rrR4/W8iYR11dK5eqkaS9gk5cuEQdsen+sfdoEh34YYIhDTver+rkYgOGiRRZE6EP8z
ja2CoE1/SuuiQu0MPdpOr8e+EmoXZuh6fq0QIOzVE/0cKKulAq8T3y9HIOOLkD4pP/IG/qcu7Wmg
Nh5mufWanqqyNUQHxTc3LcyXVWtUYV4KCUNQ1qrzTg8JZQ5DT9JQI8bJomHMVtHc/ZnNwb59V+3d
F/rwl/DJDu18fy2RhrSO0NXZzsPWaRGZTRiVA/cZoMx+1tPX6JzCtvExHjOdeUSbQP4HQm3SxIFw
Hq6PB8vqGiOe1VdA8LJ7G8xvWAA/n9Y5da4lHAe3GKmP9lER3+nSfvze3WPYkceD/5khDllqs+pe
OE5ulutrNS/gyyndwcUmujL1131wbip2ap7PFoQI9Y0GGhHc0R4hfAYS2abepvSIrR2PWWkNotIt
ACCaXZUqVe+hyMCUDIrMwgW1nEJwIzaai8S97uwtgpZHxNc1XGMyf8XcvMprZZvoqlnhEjop1hKY
hRlVCEwe4/DjnQLbQ5DlLISo4/ls/uO9w+q7lr1l8xicmVqiUHCUWY93T0XG6CDlgV9MZ1y5+nQb
sb25VP/bvUaC5ICx6kqDI9B33L9w/BG6n8INW39IrZy9HEFaBeHMszD97f78cT5oEL9nO1liJF1p
7EeZxbbhwQcvxJxsvBOibW4eHesiYkWvX78fE3QPFm4f5HPysjHiGZdyRuAjh9A3ktwrVEOHZvIc
1DVXtbhKMlMvjnqYkErw56trq4S3FeJOmga5dCkLol9l5pe8TvwvfXXPe2Kc0m3I7ZiA9dD6ALjz
mJjUs6NSP02jacU0gxTGaeK0yHztCmiDLZSvrywU2LBsG91YP5pygzjOy/qsb9ihb535igMp+HTy
4aFdLA4x+x7Fd9O91J3Qb8uWjvhAGmmmxAoiPCQti/c/7NOPnfQ79uE5f13BxK/ItVIskL6edY1a
nzodYoeszWWrPjb7ZSmUUhqC4X9zeYhsvHHYg1P6He667s70T/5vJxf1wSiNIImorwEV+9F+1/yX
ZFou4QmQDsAX30IyPr0nCdZjHFZuPAjJEO8JZJxIrvx2D1//4aMd0gZZ7tKMuSdvuhQbCsYMZ1dz
/yXIiT6IZwwUao3PvPCLTUhW9QAisX1ytjYhY96rms19H52JnLs6T5dDhybBbeF8WF1iFm29xb3i
VxVvBQd6JbNuLXZAZzpQAMYTZ5fPb0/YxDv9RAxB92QNAq0etu4FPFdwekR921fW2THpr+L6blzG
d83y5kd+LHjEsMcj/ECg3e32D8oZSgMJDCyoCuQHJroRirhcj3GVql/5Q+JFGr9pYUUsS1vIi1m3
b+T1vOOYs37+L30pyEzfqJezaNJhNtUwHgXEALG6VPRqNBI9QPfUgsed2VFjsMI2yY7vGw80QA9l
uzuj/hf7V/PADBT2+5WASvkvQP90T/QP1xFrJBYvv0LBgqM1iSBXYZ+EGtACP4OtSHFfvorPSnig
WHXJWMdPPsT3NrScR713l+R1N72MzsKzb6jemX//UFYW+8MnxrP+p/4t3WNxtWvPOw4tDf/KwdT1
Et7vNmc3SDHnupigKiELytbb0LYn7iQvhndzSE8JVTuc/uCF62SDm1k162qcxSYRDedo7vu3XAs/
lZypXLcg1xxZYILu/8xoR245Xy0cytalFKQCoasxwa52+GpS1FRVcJKFvbCY8RJ2j/5dqlw9iABH
Yq4ikYjRTpf/LnrfqSNBH8LcWFqq+HFy4TG2F/HWiHlH6rvcYZCbYETZsg34dDNhCzA4bjI4ij3R
wuLxFN1NZF09qBv+PsPqk0SOl8VHcEpe9lQynyqqS5RvrigfiC98sXc3XF/Rm6/SjQTrY77Sk8Oz
zcM6MOYdp8LYZ3lLFvyK2FijQaTPhK2uLNvqOWoKLsdP5UaJkt4H3qm5ZqEFFAnb3rUTPB4Zwh/5
F90kiTyc8TLALtJPie99U7pQKc7I4WQDqqtnTlGdO+wVweMusMlQJN6bwI28m4kZv0Rj/Lu1n7PY
x9tQRkKLrjcHjqBaBLVWp/tSvpj+vPGq7HknH6Kb8MXTGYshanzjMOH+//CKd4hcoSeAMLF44YD3
Upm8NAJcTa9AFTsHncyZb2aNb5EBCXhSnsi++4Pe7CeJJwe3Uh7upKhA7DAsCYz3HLdcbzkRCUhB
LWgtYzJ83womV3mO1UKdpIRdKu3QETEhq3HZ13eox09t1SuJpm7hPqnUX93TdFo+jtRSpZOM7gL6
0kqazMaj4+io3kO7QVc1ZJ7WAExwphwy9R1Oesmn+HnpfcmYubOU/nZoLqUwbDHR2V5Rh4r0wQPi
6FW2pbbhiWBmu28sx+em2bxgvMGMgxne6FBj8I1F7w4Cw2Ppr/zKjAt6Y3jFWWUX16AufhIHF8Bl
BVcJ7ePkZxYmT5nTmMDdHlzlXAz+S/C05FTWlrO8ph6Mw0P1tp1yxnVBoR9GALnlvqpPc2oHbCg6
o1JpLRcjmbd2Ulu2l2uS8C4eTp2gF8EuuVNNWZ7+0ZDuXcz6kXjjYaG0ArDhYp4BFZ0B1S7oaoOi
sfyKT8KDZZrgOtDKHUOzR6hM+NS1TMRKD5DhuF/WGoJ0XfaadK/QDLupRwJVlo24RnzbVnGIB2IH
rfxfB45Q5OZTBIbzFLZ0oY5sv9cOchqtIh2P2GdIH2J5byqqxTwsob3UBYvoRUqiBB5cOzQfv/de
i0QVXr6ysg+iabXcKytzPgCoYgX2WC9fu61uVJGeBg2SB56x15dOwHJ3SXH9aZF8eoDwmBbqdCx7
MZEsFlyJR+6XTNeLNOcpwMC/XE+rJDK+fjRGFGodtKMPH+v7Cqlw+ce56ajWPftmzfbpoFcrW+Im
TieydwjIe4AK+rnOGRChrtk0aTcTosCkye6uyu630XOF6FmOaQ0/gpvTFPb6cDUEQ3L12VxHN2BW
eRw/CSwyxiizHfEV5eDlz3jJnPCH/g0A2GL95eiqsdXQSh7Gmu+vde5eX2IgViMPP0O6dLiEqeNq
B2E8qWKlN5NZpRo3VPgxCs8ttip737esxbphfDrih8/j7M5hwfGJzlH3CW6gX060hWcT2bQzufPH
2qmZZ/t2YdMu4VxVyss2ChRX9HG3UUwPI9k1yl+c3FA+E0FdS7ClMGp/L7Nwsae+0p4K1G9YA9R3
Yog9Od43sPl3/PwaI1TKSGyj7Qx4JRVrT3txwOn4qoVGJ7m0YeEOAVTZa++PKX+L8/b8KbNSnmdO
5uzulvhXJ18DIbJ30bnvdQMIzP8OIj0WDb5yC5GqwFcaiPVYBLr46dggIV/VKGGSv0IcjrLNqFeD
6u1+j6dDS4cgnabaxfC3CpMf4Ym2OQgLRUnMCW1viGLcvzyMBvtoZQP87wJG8/eqCvBvg+u68o1q
IcuEYIZOqam6cIxxyp/UXti1j8sHiOybY17GcPj8vlh/8lS4nR4jcc0juwZq7vzVJ1dk2hrzYzPd
HkHcJZjDbaUzdc6ZkIRArslNZ4X+uxN46Zee2wciZLmNJGIh0uBfLpYSlVnBLn9n1QuREzjLhhJE
j24jW6NDRxL4sonsjYsH6QFU4tledhQxtCJLjBBCmeBA853kSbM1umqXnko/otmJNZ0UYhkDcXWi
e3k6eSJhFvZgSkA2JuZmqN7Rc1f7oS9Ii7zRO8TIj/7jw8LjxV5pkuCsujmVj3H53QPLna7HO+yn
5i1gs1iHI3ABE44ZWwNe3xeyP86FNIEPKcAsS+XTXRhkeLWFM5r2qoMLuG8OLoL97eggic4N3Rod
0UVGJpS+DGX/K4sG68nLspCsqPvCqYbtkpw9Pxivrl3EyJ2xb+JJ/KJRjcfUR48tV5BoaUaOCZOK
BE3uXbOxUS3oz1o2/7IX5BS9jo7vjP2bNXPVD6cGhcidMEg9Zn2toYiAV8bFxwMm4AFDp+2yZOzQ
R72SNXfiVY54hWAtd0Kl1pODvk/LM47v6Lp3g+/0p49DuxrXHHo+7zvSN/T29LN9CtuPJVkF1kAd
r+V23JYBdGNFUTnx4lXqRS7Y7iVsJU6/dngABSgLk9pFzZLM7VskimoGIe96y9ofWvnPKNSQmAzY
HOxOZiVrPnCzDZIhFZL7QHAWp7NP6JwJdEwoF9KBJF6rig8shlhptZc9gbAPIVa4xojlo3DRxdKG
QGTjgtwzKo0LMHmSG0gJu+BW7OU5k2G/0S8vR18jOM1pNntsZAD94yIvzJRz14eNdKXnk9AxEmv9
YcKXy/cMZidORrE0YTFMN8ar3L1u6zXGZhcypcEvhe7A9eTiEyWt2O8H86V3iGbyRVGRT6OJr4CG
VxESXWOkrMxd2wBRohQ2CUCYt1hi5blEVDEmHfth3PGIgmnxp1m8r1H0QokXv3Y5x8MFhR4psem3
ZcPjC3jw+ry0geZ4Hg15l2N0XuKaREZnEf79/vIlVwpddhpgNRYk+X4cNr0yqF08YBFZ8a7qF5vB
vh5w6dW1/bbgB30+MEZcPBHwfyWqyY5LTLbNe9NvaQ4JuaCPRwZKqWZKQWtUG4Lcy8Ocpv84wH7C
8yF6LD6hDVH1u+7AFE5QuGyUNmyoAEDpn35oHZIiJKVr0C1AFCsEWKSXk7r10BYVxhGsxTRZjZ5w
rU9WicKHuSq8wHjPcWBF9ze+njuQCyWV21Yc6VFbfjS9NV1gf3eKEeuggDzfIy5Lxr0yOO/Tw9Ub
5mYoUNxKYBp1XL0VrKr8phWgaf/9ZIT+LIhG1QXqGqFSW25NNulp1GSBXoLt/NmfzUEJvdGPDxWD
EhRg4j0V4YpWW7f49yQSGdHTZxVz6KUEC4/lu//baIfH7wnV5X6hWH/2jYPHPISiJ9l4/ylXHSoE
BVb/ssIoFenCFQ3Ua9oGmOGb7gWjB6hCJXHX0uGqSXOeH7riPaLSoyC708Yst7DCEIB+v/363Ikr
nl2m2X/IkNV/w/EhqBZDc+5jlUqPhLxQPUS1OfQZ9WRLbPrZe4I6V6j0Xr8uOJntxoxp/AEP/7Tx
cRrc5epV9WmV7mPmdsxaCEArED0rtXc9G+kGfhXBHtAQKBereWf0+XL28FvT20+CzRlPmwMFcpj1
rqSfUeNbIrUtonRgcVNokfwfr3K4NNtLA2Lb3iIf+DBXhChfKYm+85CIcjVcinBHtJYXBJbritPP
qLPuAj9d6UHXT7zh+Kx2GnWwRBkzMlVHyZUUxtGvPixOpmIn818WuG/1mQ2ltRoi57KZ1I8XwkK9
eesS4GHtmN54jvgBZCOeeisK7m9s2eiAN0QHYFXWncQnR1pwg1BQA3OPou8DG1ZPFElnM0IhOUiz
sVmDJy5GxWMivrITj0svTGtNi/35yv7a9Ct83NKPb+/KcCYTMMD69U3ExpuI1xr9qBklDzcqtpbB
Q/G4pael1yTtp6gOJTMNyvF6JyBi0QphjPxWqgEfJzTLYSPIw/UwVLP0fqYK4hNQgdgZrbsg/xiO
iZ2d8mOxAT4xqo7iUVPdFsBLHVRV9Oac54fyn8OEnNwkOiJcj/WXATrtmlmdUshuRQIsQUWw3TH7
/4n4+www7hmVu/lC+xQBuhGC3RyTy1nUn9vyp2pI/UDCOENuGNrtFhsgpD1uiW0d8kO1afklO5bt
BXJxc2LCfY5R28R6dUk3mpyA7Knt4Ngel6Kv5Gj6kV5goytQNGF5njBemOSn1QJONroOZdr4Ry3M
oP2QtuwMLR9zJvV43Pnr4xRcXj1POtZZAncm++L87RTAJBzYglHm68z0ImqEwntmQOYOZxsu+veT
IM67NmAeaMAOqKlXTG0lwuKb0uGFV8PkoPMO0Ryxmy3i5K3qSEKU3+KknxxHUCUcHlVbWw9SXCrz
0Kyq4H3O/V8g4CQoNenJ7psA9Ad35R+rL9HgnUYNR/S3QdCs6rbcleVZs2MPDuXqpmPDnlpwpSvl
eKrvoYUvwfnJ8GcdeJI/F3gHqwxulOX/1mhnkM7jhT5eE3TklGqV9V66tgJQc8wEOWdTkQoDHoGL
Rj05jjXn++oVI8iiz0Z6BgOtRvHsi+57qMGVgvxGd7Q8Wv3eRS6pOeyzg714JCXk98/GI40sk71l
cvrJ4Je6qCmuBTKmiwTlPifCQAxippsrWSEil6PxRSxBBMzcIUmmwjJavNJCcqgapOV8vH1MFub9
nlKNlbVwGY3XDD/XbQiD8R1OgDSdgZnOoBXjGMwj1H9CJ5qvjaRd8rIQmHzyC9ffgVKdyY9oytpM
SJFf4Q2DRJObPlYSrFqZkOuwzo8BUb+PmSz0vJ0NFjst2h1WcMlXci1XDGYmU/QICc+AaUmlBbka
btK1NnpmGFHyM3HyAPROKvkxYGeZwL8BgzXPxVyk9H+2tqDbdv4YjJQxTWaOt01Z7Ch+9UvF85uV
e1A1IjY0EZXFvZ0VjteSKyoScrY6NNFL5/r5TyhYJnlDfSPhe+3kPQFyrYmjf99y0BaHBcNsIxlh
bLEvTidRDyV0bt59tAH3AlDecUIGSTqts36R3TxcF6SOXwzE9yVDS4wq106dKYUgLBa8Cy4bXhiM
lF0sexjbQ/uwxdSlo+/tdy6lGVZR8VrbkQ1hTx17js28K6Yv+gdL9JAYRbRHw83Zq3PrUq3l0PY7
x9RsRe6dHS4tBLQs0hPekbSUWnGg8AJ64MEG2wk7GW57WMTHGdJa6PGem+PdllqlfK/dvD1BsmJz
Spro1OuCW1Qae1iyT5r1feXIb2NQ6fzRGhVKJ4eMuTTSqnlasAJMmbG646mcT82nu5vYA1B66F82
xhXy5K97MjcQADu06CbjRDDDcqBdty9H0VuW1wMwJC0/Dkbv1DWwX//A25B+aSlHd5PVTosagolQ
WAdFhuS74lF8lmmZVQUojqIVA1eqXrtt34XT5o9PyEtKnBRfSOWvShwbKdJlat7529ITdMbBA1n/
6ryRb3cRKFrJh+Rgu0zbPdb2lkuxgvGLH/C7JRaHR4zOcYcQlXMLomeyqXBJjmB01EDQY4IZiINz
r/5gArN4AawFPLPgiG8ICLZrLCtXMEE4yRVlgn7vZEIxwHNJrVpyLSv8CFgvoFq90+MZmr4u+n45
kUL1estIEQpeKLb8yYW+H4IBhjjZXUXmelTotnsezif0QPQJNmLsIlEkrOyNHlweqc5KWCfI2J2y
QmPjOluebdyLfdmPWsr16TTcqUzETwFep+DZferRtoLBQhNWGIboN7X1S+LlcRUxb1UcwfOHqokG
V8wwuZHc4HPzxgP6i0o82r3xFnLa+UW3w/HmgrWS1BUGvucVoijbq3EkORZBZxrgVOpSOI4raREF
a1uzrMNPfgGoN8Q3zcTxEjdgAdkn779Z6xBm0EH3QTFP8e8ukgDlOL8l7R+zvGZXy27cBdYVUQCv
MeBNe2xOvT7avnaoqHFn9A5EaYkHr7Z1Ttb0qg5T3sbM4gdnbbcZ5TTH+M4VrM2HAgiaqREz38DH
60sQbbHsmcCzwtfQiFNLHs5SAyXylzvVtO1b1cKHC6n+RVVPy84dARUPfpxT3Jkh34QLSKNGNQ+y
aApYJzFUq5fcHtztTGx5zOhD9qjkTkkiaQPB6aXXtDqELInkNk2O0nRxtRWdKHQxdn5Ob+1x3gk0
6/g4JPO3WfcdoX/uxqrOKdJWwxrFYicztB7UOo6kq424nfhukTwQF3epzPTQGHT3D4A1spvXVdR9
zLnKP1aJjkkvR+MbIUzBy7np0VJTqOU6LrjWhLMH/D4RzjM7q/158wOmBhjqpMkR1JnFU0dopdS1
ygNvsfAEHtcnEP49AooAWWF/I6vk7NTgUetdpKtzc7+/fERleFoSgtDh5nl92MTQyP7ZrrYuzFhQ
Px310nQ7vFT/TOjBZq5E5rQ/NAN8hoSn5y7CjmbiR6yHFoAdvKExGpxdJE5htDtl6ouiNUXc1KMc
GNO6cfEGMagj7Be1vY/r1OStVm0JebNRCoBVAWOFOz7e+wQMSW+5VjEXjBayVTNXcGEHsKvTcH6G
3z+QYOpoe+qtbEwpU0pSgYNVB7QfKot8SoSOSgnXLsb+asZlR9q/Rg1sSn1yFkIXdXH90dR/Qhju
IRvxY40x65q7j0Q5b1w+w288kLOocVHgzfE8ctSfz93o7K0bkVhmQ6zfWCysHL7JDiFgNc99uQcJ
1qPWrIqivVXhU5r/dPXDflaunj/XYU1+Rq7bnNYufFwZoj8v/tWU0m4MAeps8PfAYWQhJ53HD2L5
+URO3+JF7066Kp9kJK1rMvCMlIFLtMosICsLEyjBa+swKczLEykvwBNn7K1kHCVr+HhJFWpi7Gx8
5Xn0WyCQOoxH0r+PxXMSQQbWH5qPP3WidGdDRTYqet7jFIgLdqDjhaH8lNC5dPgqe5runKCvDL37
6XgvMqub8oyn5Hrncki/voRpf6QaEAS01dCW7tjCE5Zmd0PsKRbrgAOzv1HSQdWsIdIire2IEqCn
s1jD4vYOL/D1t2qi73MALFlKjFaFVRTmyH/r8zgFD6yVczbu0H8KTtEkknI6UQF4AD7b4aacX0m3
ccHOlcRToL+asDh0Pts8+5ikcP4zu7MEUz3bJeRpQlI7KK5dbEdeaAK9tRb1w3Mr5ivp4h7CqpcM
MDalSy19Fe2KXrkf5ZnhGseBH9QzLT884FbAFqv3HXIBN+YboKmlTjbhs4968AMIsWie323hkWh9
nMYgBelBIriqW+rIDpSxaJa+/7y2YCbe7x2Axn1IgqjpV0V0jxItc7doFBKBfi6HrafBTCPPn2TE
ukFsQKEc+KVsVpOpj35tY8wX7LXhk3oeAg+Vm4jZrFouPzRCZoJEbNzhGTfTDCL8c37SxGAvPEPk
DBEccIwX1EpS3rmVAyyj8s0icsvxZPYqlBPkhZWjQNsItbv5gA2Fxtg13SXMIAjb0CC2HXM2a51x
aldKOGB5gK8lGBSYAVDTsBR+6xySZr6jFqms6eGm6RETF5rEi0xyZGH3mkuwpyUi7u4s9tZFkUK+
30HxXTmM98uEGaOduwAJS6Se/dpiJpDLfPxadQ9lejPERYD21d//cVaTI2Zolg3+0sonPGBfKfRH
eoe1sl/2n/CsheGSjLi9CextFbd1U5GH3HvJjp8Oi+6oTQsEVHTL4/gSf4fjJNP16gDOm9hj6cGz
7bS2kSIEdez9aH2QurkPdRGvnxYLKEgybyHjNbC6GNEQBtL7ozaDR3vXwVrS8gC6rJQoJBDFiJ+J
4MZ8Mx1NPsyWEfybQ/aTiURuJPobc6zJGwshpdAeypUyRfze0YO426HandOIY2m9/0k7DclV+yHS
evHWI83Zff0aXc//JX4EVEcjT7ysrHVGRQszB40bhwtBWcfq1VlIdvDc9jSm6JzZWMHAs0MYE6G/
iRd+DCXh2zN5C/gio8XhhdlKdWJPJ6+S8oJQCmhJcWHk1339rO+VWCF+iaiBdolA2gCZLRCdaSEk
aPzXe3e/TdjfzVZKhugCLlLsi3NBEAVW4OY5ke9bqC92M2hayw9VGzWvBs2ftYNh2J5VgygMY6Uu
wFDK8DhMGEg5uuCfFoGT4cyXGUcuhpw3jQNWRWJtCMZiTwKLbjT1xyYccTiv3mohzejxTrPmncww
zweAa1SISXrffT0Hzlhb8X1kM2EvzmEFBWuT9oCfzxUDvCnSw2soRr09X2xHKgFztI39NxqKTzLY
hcbYaexSQ7CG2PMm880rEUVrms1VOox30HgmU/sWRurY7m5WjohhD8/MHVJtFAobJiiOR1Nm53ez
gZhxruKtcnJL7vx8W3WXLAi0Rz7KdtRZLEcNARZgzNXqMiMHPnK9x30b4VOkWBCWk1MqFOMXFvW+
Yy9yDCWeB0g2I7rTAAEJRpt6tk8CFx5B0HvABK3L0fK6o0Y4J7HaQw0huRo5QmFOthEH9r16rdOR
kEtUJ4a/BKt70pK9uak8bNVse8Fwa+R7mdT0bV/B9XnnM2JXcZvytpV5M+8QnDa7CdrbjCdYNoxA
W0nAa92iSl1EZn8zX+o281v+AuO4q8A8+LopXdi6Qs+ua07LAY8HP6FDSnx9+bwOe4lE6U4PTTBc
8KwBlkka6ObCX6mTW3fgtG8gBInQri3h7eqjIaa0FiF2WfDohKdAF7F5MRytz8TGgtGDq1IkvUMB
oPzre573SYmr8PkwOGJlNpM1KFbRcIxacy+jxTHwaKlWDC8NoILpU+Elt041aceqb75TFHNwNXoj
jpRztUtZWPCoWX1+hkDHlm4dqNMQkfVZnlNAf7tiBCveUhObDyGq/wLCj4YDSrjhqumZZ28oO2mb
o+R8wRa5WAXachJcW5WgkRIXOmO9GdNFnH3SPhkUDkNq/QiPE7y3Rlwbce5qwQz4xry0Ty7AwjhC
gWxcB5AFmHiqLHdfwNQPhs12sboQo0jS3r3RHnX/21HJPFx1yZ0ju51BiAl90HDSf/blpZG2Pt0o
Htbhj9gNku2EkqQOGAgvvio3sLaSoLZbHV6uQzXuqF53bA3UB67W1dbyZdhkfpx2QQAWdCXsEbgz
DW2EnvIESUb1lGXLLfCXThbqO44NvDt+2exI84WmzKhiXqACit/TCCrdSCzokSyRmj504nQT2QjU
FBQISXZLH6ZLE78UboNp60J/XgjAUcOwyhqr1XvnBnYdaW1qBuRxGbX7tQk0eS3TinCxTvNb++v7
QkkJ1a1fkyA0qBAk2QN3xZMUytDtSSBOdEcexZRIN1v58XIKO8BQVvoyrxlv/XHARW0biJ8Miv3U
3K7v7U31ciNSBYZqmKJABkkTj685eHPdtui8Rt7iEF1SHNosdzvAwNH/LhaC1r+eN/PoCuLJ6QBe
Ejsa6Xus39dBnAx8PNPKg4e4zXmsYePF3yO877LXBQynCOnYkcogK5gGLcIV2/yXGv/kb8tK0G+z
5KcJ6nwlZn8v0LvWriV87Xwq4ZX4c17i/31EYqbeDH/AKMJWdv8u0vGtfENln8mAYtKVyuFSa1df
N/1skJZ/YuWYTRALXM8d655jqCV+4XBCkSd63Lu6+hk20Ez5IXArd7wQi2PKtkx+QCccQYSe+i6X
psdCTr6u9XVAbuVjNXbbBQTWA6yv8bywa3uzRFV8GSmQMuDzLgX6U2Fzs5TD7/ltLox17l7O8uUE
LdgcZ5Tk8k4Hz33te8NXnDB+1lnlKGC7ezWO3bh4Ze4wTTKlvyOaL8uU6lWqXbL1DdlkZMJ7wtzt
5xnoyvNkVEeuyLKN8Gku1b+JElCes4anA2L6BGW+1wo02W4j14sbOiiH9svkTXGOORlw1GzX9UXd
3mgoMd+PAV9xB07uEKweahzBJjXDNMcSXXKN+GR6Y7DmvW+4odYzY7NkzqEwA8QZ3MkrUaLV2u86
yTjMrVv/oRDFluK3EwHkt/s4RW47YRG9HlKRJgwVT6EzAMN6Re+al2Xb3K/YDcMwmogQZ/EMXCM1
Yci8FneVayVRmJ5kXVv3mj/1NtCGHWp3wx6PDvxzQwogYW2MvZIlrIx2IHzsGpYCqPtb/fw83ANu
EuxAfUnzmhOD9tjYInRtA3YWchvrzL4GX+flAulhBqQYktY6YUIdi1YhUSxD1X+QrwbiDz4iXOvV
s+OmVGj8HPBOX/Uas2bBUpZoGkQl5JUkq7ZRWGE/kZ3CRIYg4NX1iHZzNkery4o2FxWypcR97Unr
3NW5p1Ijx2kJDC5p36iCmx/Si5ubZ9OOuHF10dwU8VO5LdeTzBsEXthMo4m+Bf6FGqkUghYoBid0
ZG9zxiSJKzgpykgK5Kxepg7VzcVdV1ZrHmcdrxbj0qxZf+4s1OjC9udjl5lS3Mp93quJ4m8z8PQl
DthUgoV40mSBygUJQrvV4WzfMtAeGImu8Eh1OGtGX7JQP7Cvyai+T+06Bvn38yrsP14updJNWsDh
YdLtHgLoZyfnV/1YOPdFg38Yb+LCNV2R708PZP5tbCqpbDeoHfAzwj81OFkdVekbsGuvOW22omld
eP3DS0+Ytf9fS2AiPBROV/3+6Xg+4ZwkI2NWqDZfa8Tt0PKezBbi939Y2GSjvGv8k+yJYhItT5VP
FU+EoA1moKbKF0f/66A6oGLfnnNvtI8yKVCyVYjrDv+IXTqt4DGJmSCzE/7NonJsO/Y/vQSTjnC4
gMEjlLKVMHyXjYBYSq1gASSJ2az9XJYWs4zLXxpLFshPzluAb7cEnurcjgRsabnY5tNEPcbfYT5t
bJwnSrBhKSS5BM8fRnHa40pmkhRZ8yx3MUkRbK+Nj/bcxCqXMHqmnjix6WI8gNIk1A+N0lCkXDSO
p1b/nbuIY3K7gw61QjqGLjxzN1JkLg1s6iByceItzoY/L8G4iedh4+6fFjRdIN2QsLu14KHta0Gq
KFwecVG6yDg90x51D+hRhFUYw34lkjVF37bm2IdfIykw3DJcUBmMEkgUKUkiuK9WzU7nU0ao/X/c
3Z3bRHQhhBQRFrAWDs1daNqsHX2rHuoZFAMKdWZnBqs7Hat7/8YNVQZA6XtAkYszpCwiZYO0x/Tm
RZwhy8r50JPurlzHZzLGEjm11uKzPzwwVvPLcY6NWjBack/gos0GCAnlq1SdB5uas8q7fExTvq2B
LVER/tZSNqXDn0MsNVn8PSdLeZ2Rghq6CqQVRa+34Hb17EqTrK42baJvC7bN8lsqSxv5ZjgXJP7z
ijz06uQKXcB514Sivgf2rc2+r6bqFs7NQ5RwhCJbEO54BwV653M41UC+x6SQvT5wgcKRcvDFXcZM
qCOY2grvvXwUEBpSyUg5UW/Pd8lTjXINnRuqwEGhtcbG/ygsmDhKLbgeqUkEFjG9R3qXa50Rybmr
riFj5iodruzmP0R3M87kesnxWfYrtUtTLYZ7ZuLABzcAPJKGyzqZ9nZjnQ8f1lVEblRZNfjwYw4D
VOjvHRkisQnVcuFupvpEoDvbWM3LArfN+IM1eV/iAsq22CKfqTuIdL/e9wx0NASpFNEBN+xQsk/q
+sKIu9wvY9tFsGyL2JrWEOUcgXAYc5+JdzIBIUzjqgMPBF5V2TopIAkIIwzx2s/WjPvfTeYLz+SS
TYen6SEU8rdOrfjD4XHlX0YuOOeutCrRaVEmksQASEDnI87c2ee/GpgthhkzAOknS4ChGnPrvhSg
qD2c7aJPmK0KUYIj6qwP1YKp51+m3WMYXOMRGIAtBLwZLHErFc7sQuraBT+MLPxjwa0mAV9jr9ri
p2esoVIbHwbXsDBUsv6PLdp8avTIp76mKCW9OfROU3wzC/bhWqSJWPSvK/uucdO3Gl76tmDWiRrS
nO3I3JjynAzYX/mexlAlJIiOyw2kqH4kqN4KA6WrY8fZD5kxaboB8krcWZ7jRKdyMRE0QqSPXhVU
NZkEx5S6LvUyJZQyQMfZGZ5ZWknKl/U6si+thmQKug9+cG1CULHe8Flv+tH8ZI9nhet4oa5eQku2
vILcdDwiL2kXz7zZoStWYumqWCJtn0TLO0laM+OugRj7rO9WX4rdw+BwNg0e5qlu4+3Wz9FXQjJv
eA5ctKiVRIOhzByBdHbETQiwbLVTwekvkTLegGxu9tuMnhHY9JF8rsK3OD26LETBVGG1Qd6m0U3b
x3SSnkJkyGkGDc9EByHaOx77hvrOLEX5dwk3EiXAqG9STRGBexRJOrWE4ORZsbrZzY2VgnrtLUvG
eWa7TNC66dFNVUvGcvPzlP0PWIpJcx03rzHZ0TNOx1VuBaoGOJmffzZxNEjkqfsUjVGoY/eWKUz8
FOi3aRW1z8DsR9vmD5tVph5q2yUYFkXxdDichlZl3K2fKKnDToxhI6o0+jk9LzJJet0CLiBAP2Ce
sOc9BYyhimtwA4mBddViKBDojjBBLGFCFbAGiXYwbxdzZfxKLl+cBGonphf3taQghL1iumW6EQxg
zfItDZ+/27kozh5UXaU5CtkHGFwAod0iZE0SvdGyQpA5NPEXGYP4nkVHmHDPh0H57BAmuK20atDX
QVc/4DxLgAUe4gq7WoLzMqVkwu/4QWMKsigYi6clcn3R8VgFyZozxOPoS37gmwvfrsM+MNS1WlVF
rXpyDVHKzgZOQ8/FexS98Ul0B5kIG0Jj6pgCH4zElRMIjN+/kzFgnSyJlyr+Qv4yILc7dTygcxQ6
8/6Dr6juV2AHWPPNi2dZ99W+xPaOWTnqDej+qd7gHQJyAyx+0k49x3mHJ22ztDrLW4txbDC/vd7p
Bi6Z9HD6RpD0NW+IAjQNsYHm4a8xsxhsLedoCRgBjgkeXOmHHjhdmGZPfc9pqA0y6eQMK7tQzRaz
YBWbGJwYx299ivlc0mmsRPYzUm/xM57FSU0yn5Geaph6ieiAutO9CxcsF1ErAA8M3ZS6Gbr1irUz
pNsKuL622nXNRXGvm07px02j8OaggQNV6v7RaIk6GZ4y9D0vai2XoArhAO4cDzmNeZ+b5y+aprr1
k2DQIJnho4+pObDk+QSQi+1RAkVZYg/LYVvy0XWRSiROj6h4SKNhcHP6BK5j3fHf70cLL89yWOwa
RorqGG2662bLjsKvUkgN5crCJVWFfnEVjFI0Z5lGRsqeCz+m32H1IL8PYy4IZ38IaV+K5tUGoKHt
k2bESB77XzFL9nWbs4hjkgFQ+Mx5EIhXjXByn/375JT1uq0GA6IYex/O0fWVY1xCyTY7gFjnyZKk
8bd9g5hjB7pXb7zNBgQNHBI7bKLLhDvKIzaFcdpQ+6x5AYxqWkgv1VGjkeH3hL90HvNuKQQ45l4o
OZv9NnNABUhUY1MawaxfQXUmGpFbgZ28kOB9JB8N17QpfRvEAxgWvziyQU4QL/RXScT+FTJXQg5h
w2ou5mpVjXtOnFoA5GMW5WtOPF5soloRrtSbAzFTSfHqz+4rtQScjbeV8KfvoTAhJSsnHsQbr3pm
J5yr7+//pJDAvWbj8pab1HH0EtALtj3Wk2XOFsw/CeyP8PqlukUQpIHjo7cdt6zZ2Sr4dCMT/d2U
rNoGhEF0iGOyhCNnfcIHnxAWkdxCdPfUqBo+7xU+4lpHZSJrdSq/Uj0qACZ5LtwklO27SmKEMRc4
jTSTY06HFzwnnLma2rmy4E/LHVfb6yhnK+qcb5Dc7DmcqRJpsowqUWqEnodRr8zI7OzlR45lodBL
34SpgX8/l0XTX4KrMDpgEwj5243kGiUWAc1jDylMywH6BnxmKDy6bPxoVI+Y/Nk/VYUESUU9h/bI
7yxUw2hhdSqjtedtGZPdq9HtBiZ54df4rOGxmsUfNyTq4vhQkP13wFdCh5aLC/4l0hxv/eO0u7Ww
IyCgFpY9Q1S88NMSFkzoCvDZxFOHUrSPsEFvt2vLZ1VUCeSvtcM1bPdGAWLl/oqsgRDz5idKZLs+
UqOIRSnenztsIjL5ZtuvnHHUhpW5qVvFFLjBfeW+g9WyF7yJYN+0oS2ovCHl9zkQmv+F+rTry1Mw
TzyfqHDS6+WhH6kdYQIONDq338hfHSCrEsqyc/jSqCYjLCqgA7bJVloRDpYFoYxstBJf1rewC9vt
aJNyC/XWi4YgHkgsjiyqP6yWaE4rvKT03dUqNH5FElVl4vrdf2zUECv5ffi8c9EOL1mR8Zc+xaSh
YV45O0VPWtttgvFKR0z6F2I3vt9IksejvIG0BzgKNtlScqDi4/AeJameQbh+gHqtxicGi9SgyGdr
c/G8mSjLwJR1XzV3ewnzIRWHYl2CKgIQqcJdhgXcoJNrD8m5ckecByHO24Stch/om0YON0pZkl+d
6fu1nk0SE7xe4eaSqgrGMRqY9psRAOABYxlDbltH7SmJL9TeWz/YCwHP/ZiBHrryU+62RFc+KUcX
menZDAodgM2/xpnPjFUQVE1FIyOM9OhahpDNDTIel/Q/X1TEKhPmXN9sQZEmAWR0VeTP+cvMdhMa
Cf1a9JiYp4wtAjlsPWZpAFNnKY7y7lEQelMy6PhS1eJWAnK/KUZ3VL1OWSiFzU29NxD1VdRkiUA4
Y+Lc9wbJBuByj8tB0MOamY3lTQ2xceFNM4AiNr5kjxL7UkBzQi4F3rAZcP9QZRYXKpN4zsd+wTDo
1+EzIRCWODv7l9/OpRf2q0hfyMdcpZpN8QXlmsSiPsuNlx+glgmz98JwaTfHpIUu/l0Y+hdrdvj4
H6YEiXyZD1f0+x8fypdyNo4isQTiSpVh+O5wHvNmzT9pyKwSSgeKvbyLhQkuyiz3ImuItP5R/tE1
stTwjFkdaQn448xyI9vvNrxEN/KpFxIXJj5piHdxeKRQcnF0h3gOmhBrzLoRA5t/ahacERPjOHYp
0W+99G1rYBX6xLlWS5WkCrjIPRijrMSGeyDplRfuOdyImZrotXaZkuh3lVfaKQQdma2OyqwNZB2N
OyPUzdurfywyI/luWDfNvpoI4cRZslOnJpOSYE7ZrorvKWNb9yBNZiSOcEs3otp5QV9HEBs5AJmZ
FpUJ6RYCqNfXjbptlatxErCVN5W6Mop32cLl7Z+o+WQqXWR86zGJ+NwCGYbjdp9yg1FWpoKl7yz2
Vkrrmm0PSEVGrIoOlTXUUnHEnZixCLkt62ggEEm7/LXBfF3Y2DUvaEaoKQgAinrf5n8iXaYDoWf6
POijcaRxtouwUtFhJItTtZzHPEa9a/u1ku60FMEy3W/eHiHq2OnDDrjrHeeTOb10EIVZjl+hNyHG
gfKS1F02t9uZYBx3ENf4dah2dK8oLl3kZAuefBWwUFE+dqSM3Rewfj2zRgQaCXY6pQ15p8aVlkUL
92CA8Nx7HhCZRgcofbw8izPUT0visT+Q5NU78BpFMunWdnhptrvKSWFwy/gLzpVS08+ebdlQsA0L
UWxNdL2Whghvmxu0YAQuwEX/yILF0kHmz8Kb+QrbYlrRgSR0lL6iqguMucTIQ+Z/hnsfsM7SD0fd
rq/RrlqTKWsZh9TYktyJuyzhAXE2ADnBRQSat/DkrUhjs+iYqht0Qy5k27T8IB36MkaP4hQvBK8s
SNdfu3enZPPDmPqyAiCUjtT0IWZZXnQpETWObVTrLwYIV+fcfD6txaAmryB+j4zDX8J/Wi1HyvSx
y/LB7kox0FQeDGAYLVzKJv6yq6fXUYTK33vgg75wkk1NPvEhjyjJG3HLJlUFfhvdu5MrxVLAhbkW
19laB56otv3hpACsfIh63aK/g3gqvMzDAYd5ufZZAMtLIqqY4d9F1gqpRQwbhNjIvqm39fmYHiyV
W+kYDAMzpqJOjy9Vr8cdp/+OkiLDbeUsbf09cgsGeS2xE/b+rQgdKtb9K6NrF7b/xVbxaYYUXLjR
J6NrbaHIfCpRijllN6jYPp0oeuLlZeIozc8NAjNbpL3D23V2+iO/TaMmedLVDD6o5ERtXaodMHRp
Arr8ztGTk2pXk7pR6BA2kONrxenab9gqX2zIVg0Pq9lhz49cQG/3C+jdH8GAEK4bcAAwwQaD9DcK
l+c+R+rtq0QQqzeW0FE8xzy37HL/i05puKHFPoOthTeb68EM8gI35ap9gEg8U/bQPZEz3fmgFAPo
mnfX2URlzU5730MBKnG07UYBm2pEZONuMGQyV4X8SaR1voCU8FxhsVRTWw7OMej2FpOZl3rM9N/P
VhkiWhqvovNB/5rfkzFxOh8QMWt8MSIViHFan6J7o/ytZY+XgkiuKW4GB3f9kpKQAyy4wgKnK34Z
H/qTxNYkMNxXoszEN4lNzaya74S/HZcMknc+0s/VwNLszW34a7ODWLcyHPqAN6sm2IoSxIvT4AYy
Qpj7ffh77lR5TR0hgRRx77NbbJsr4s2KZsDWoU+6uPTqaZu8s6HGYjzjJrs4oIbnmW6vSPSEZawm
nHzHi/v8WqYGItZ9S2gFuLwhwDaXZYEE6nk4e8EguDwO9Nnex/Mb4IOlTrMVEEdUqoUai/KX8cGw
jg2sU1GqtRVft6FRhzppNsF1eeqDYA7MAK7wUUvAMoIFdRsZMePJlmLQUmj703WjCUj2L+kpNvRH
bRDtm+o+EzOGCOjqfEA4n+oiLSHikB1AQl+ZdvQOY1NCW12IBkh9RrwT51xizEO/M4e5T3wDo2qA
bzKpGajLr3LpY7nrFq7VokycBUlp+tPhx3CD8sepiJ4VAzqL0uL3RrRwRhEXLdHDDk9ZHRzPsoiy
n0uv29Zo9aNeaIDDa6e6wLMOTksmuNA+mZnq9diEacoh163KMVWBXnwDvE308yVwIcf0uusi/0QG
ubEdd223NV14T3NkowKFQnFiSuuqBXIZzslJp0W45j3FpCxYbTuLxV4AlXddUZDolD7IZLxLHaiT
7nrqrT+HHzZ6Xk6HepgZJo1Oc96iw5dPocIF5qQ5phS7caEUcHrUxQKRbVcMwevn7y6eepBHpArk
NMu5u7L6CXI/fayARsKZl5RuBfTPuipc/17yU/tDme7gp3eNNtJAVKvWhDJC0lQXkz2VpMBEIC/Q
ODIlmyfRt7oIL/uG9xNLQK3PeOnSv710WG+IyxtoxCi1FakxeUcpiX6c8Rgsht0+9+OBY7CvLTeR
1pWeWCnKwjKpkl/TUzh2LKLM1isYAlzgZvn0VKq7hQXZbTJY/RerlZxjTPxtHDPMcTaELtMumvBr
zX53Hg5oVZqBTNi8uQp9zrDYILJg4QmZmyIxHiXlIJy0PKMpxj9s+9Hp9YAAbRCanmQU3mZpgzq1
ygEFwwUGs0FjdjCQsNZ3HYx6xkd6Kx0mKAsWmaEmHDiWYzv2FnUv9+xGiZEdoEvRmaC8CqbCtVBM
K/lnGRlCCsJARv98TfykUdTA+UWMlHqfcSsDfd53oEgvSCtQsJ5g/rAniOGV2WBILBXo2EiTEYMV
FuM7beCFLQ9mj31qPjFlv13sEXlq3+I0iTNZB92lKOeTTl4s9BM2s15/Fa7M3fO7Cpt8Aj9M5/4c
fi2oF28Xe3P2E03bAUo96elgZ9raJ3U5Kb3v08GOLLT07EgmFkFYMvlb8RwG1V1nfRmuQZ2zzRzQ
7KaTlezvfACrGrHzlfnVYFXU6DCr0Bnu2yD2RjK5govSdTNGkDtoZdNIhhLt/nhoctTcLL1w3mNV
XzG0HG2VjQzf2B0Gspk/Xbh+beBTKwg9qf0xdhgVNJXb+UBpeoviER2opU/GyirT9cEmXDpHqIMb
Gmd4leMmj/1LbQVwbQM4oO3eDRkgoZM7jNqLCBBBnwgCrX5N+mdnioMWICz836xGGMGQTC7KRxm7
pPduckrzY+lcTkUqWXweobp95EvtMlLlV+h0R8ieXltwGel2E1CUO95sTULiyY1Hf87YsEARoplM
KWcpXrrzOC+sJb+xIKfKqcFnDlVFtKWgYwCbmBwv/MIRvaP8QnvSoqKMnxnVI3zfA3ZuneKpYe+6
Qo7atU7GWrPDVaG3HM+cGAb8lj8+0vFqmhQON9R6C5MEW3BpEwIchgU0xCUwUzQ0yV66+A/pqTka
/2gvhEt81e7YTuXNOtCbQKhEWs5YjzRsEZ00Be1VySrFsyZOH8WhZ2YCdvxu0Gw6PGjDmYe7TZEA
Yz5zqbpiUyTTB0H7KqMJsz73NbQGGsCjOXc09/aqjeW5IzxoqiFxhIB9o5WP/5/EOUs6iuVSs9OB
nPa0NFo+RCOUPre15vKmGTcbxLhsLoGMUfmG60iNLEaBh5k1bv8QN1d50nmhJUwQpcic8jXiEsmx
PPOcbSUTwey+ljXZ49STgy/hoJUclhvhnyzN0Hl+Hn+6tuqMIMqkGXFnXMr65xzrmKXR/gSz49tf
zVi0J80f665FPwWDQxfaZ47KUltJPgiPpiK1KYbQfdGoCr/g8MbGcPzyrQW/t6seSE7tC/Yk3zLk
9UYAEwbBHRaYN1uAK2/Zx1ehIiMuD/t7tuFWQpW44o9TkN4Y1gWQtZ9E8mR37KRnXi5er6/0nBMg
8iGy7yvY654OnQWsRFVjbIv5ODix/72tX66l9JL5fQzsIQqdrVZhdMr78gdRAbpRsNh4GvKBcJ8m
A0o5q/AsqKhQZPOsFHMUPym6nQ+ODMFXzDML9yeybqddWjDKC9PEkyWfSTtSQ0KkA5sllil/S6lv
Bl27beH7yC0FR5ecvOmyws3H6vXKGWCr2/kFk9Q/Md7W95yAFWmPmtQPo0VQ3UTUv6mx1ujM8BKY
nWe3R3WK09kUbGqoveWQxX6lis2xgZNTk5uzMos2ihZauOm9qsl0H9rCPlcYnR5uRuSauomhuN/y
azpueK58Nju0tU7ZGkmVK3KvEboiC6ll8ErPOX5OwtL2kPZjHIolOHShHj2SIORuIU96+l0EL2Ke
WMWUxNtQTlRoKJ2GiCW3Sk3F8TCuiiNkUpUdL3KVgN9DZ6I0ym+o8+ymbmH+7SxBqoY8t72ZlN6i
Y0N1VLRTyhlh2+n9UGURM5KN1aOqLc5NnXyLsUD+18SYKdnAyCaHuFDdQmSIaFO6FxuZ+4SteF6h
DewUIzCR/1KZMhQc6B3pDAZK7UV/Hf8g2WTrRVIgbwrT0EgGA1Bz5Nhh5SU5V56PoJgKSBpNVKQ3
uMx8eCT1TT8JmxKNSEGS6BZur/FeuAlBZn7MmhNbMBbPzM0+/hKuPGdFQiAkd4wZG6RI6Cvmi+OF
HXTx/RMdMz3XMOv/mMxktP7eIl7awoDFYW/PDtRHFTaNAU2gLP7sMzWoC5ao5QlZfYxnOUZjOEkU
KciEJUfySGO25fNf+M5+ownhMUAbPye95Ml6j91w4hllSESxzVtf8wYgDp/Lzn2GRmCU6hU+6NVn
eS2fg4HwT2yCVMn8EzRgsj1wsSKgpmhOF89GdiVUzC3w31eSY0xc81JIr5muhKMhJVO86UK/+Q9c
WU2JTkz/+JHMsOBzTuMGH0fnUZEc9SVtohFHv6oXuaCOkqXmQ7t5sx3+J909cOI187GRgo/7f+By
Td2vaugXchHw8hBYRZuRPpFSerkRbe0hlN/+OCNDF5myJ6T0ejfmuEr9EHHzBIeyDWuSLUopYaE2
wRr5E5ErE/HvgUdwo3pcFfWTe3HsoAj4Liap2yCu5jgAiPvx76nA5rXZBmwRE2c+XRflEP0HnWDy
AqChrVOBX9iYsFwxXydxHYgRWa/aMt8yD3B2VCfzyIpAZEVOag5kaD5+EXZhO05X1PeP5JCNf13p
p37Cds+myJ6+WZLzUPejMrSjq5s+gUQAi1CCKQfa+Mf5bdCWdn7PMGx5r5hbDyuXlOGjLMOpGnjA
2xWHWRtIAje9dez7sPi2EPd8V4zXitpquNbo5QwoblIDm87RTEZezh3O0ynKdEK0RCvM1SVIhH3j
TGi0xg49zaDGlZx19x1+rHe4fkNw1R9x83JgatPrYVAZOvHGcFfLUY//yZPHDHNJU5LqiPtJyVxe
1MFWXaIEBbJi4donRnDCriLh/4qzmcWuImQrBAKkKvgEdModAmBRrCslKU/rOpDGns5pSdKPNlyo
RzG+RmpYl/bZlXNQhh2ohPxJ2zo5wPBDYLy56AwPrUU744tdA0jpby0UY9M2Gx7ZvqjKLwmANNk3
8tfwJel/MnBIbOJD/BHv5obtFUDr0eLmMHfYa6QRTIddCPgaCSEZcvrubeRWvC2y4yxDy0V8zVHC
pD11E7bzLKKR1en7A++UXwOUUZhqFEKD2JicLdZkk0BrhAdKQJ6VGXwqAwzfOvgyEhzU7oy4k0W/
/0R8wpOBfbGGCOSqVFSj2J1oY5Fynb0vo330Jkmtv+lv4oHNOQ+S9N7f0iEQ+7HEsJURJeOS+5HO
fgvua6hMKn1oyjmfRphLfdUuXjexWcwLW0rLapYIPx6kQ3sg8u/6f8xVHwN9gRb9Wh7JhHC6Nn1E
qhZ1pncwMyaem2VGvmHTXfZ670GcEhAz8mUPk7xnGtb4LLSyAmRBMkgF/i8YWG8osB5+8IpD5prM
F5j2aABzexu0aXrTnPgvjhevK1jKjH2GsfIabuHxSrwvtPv3UxeQ6qLRdCxF/oYUatU7PLTteceN
P3IiO1GYAzBgWDDzUHwInK86iXQ00fH3J/bMA7yVIsUR44qFo7SjGN5KyWyWrB138A5YRbc6uzu3
Vc76McfCeC3PR6rmm2aE4cMqDnX23ADg9Gk4Xl5d1G1ZImsZobGlTG9WL0DkKgEZHhFiN7syrwdN
gDT3WZhiF0QrUXenNIKAHDhr96n6J8D1CkJyoujAm3qRzXCGS9RJeO/O2i7HjcbsOoun7PsMP+gz
JBKWiXid2s+fP+eaBefPxFSuK2JAeT1xYlOLlmPiheaW0YGQHWPBST0+ZWZ3A7fFqDceJZ4jhxVr
htyBWgh5Mb/6QcKw16tQkua84DTHjJajn9m7YPnsTyXsLCd0Wuwy85fOLg0lafJ1Sxb8g/WGvt2d
9ZJnrJeHa24xa7CARL+YGOklWKIJwlWN66r1ydFPHDk08xyPU8IqJsdg2EedX2HIQzfZ8cV+CY0W
9SaeK5C/opYus7a1Ti/fuuKpXz/gFfFbk146w42EQl4eVuNciNvF/3me1fXg2OM71u8oKU3NTzVa
PzcKFO7+as0n1ywurQL3yLeL7B9RslKMIiT8BlQQjUEaubQmasqB0wREn8uexC3x1zMzq9YUuI3I
/y8J3pE/3Loy/Tr9jXf0Gm8hyQ3ncWGxNb/jgv7yPxfE5/Jim2jcIVN2HiBvv/HnGZkhrnKbGdnI
reXrmQwqyU4aVhc6gG/UoprI9w9lkuQTvS9gXDd0jrOoxGhVuAYKdDcptxIeCjd1Mew88EXhTWRP
fZdN9QmuiSgIFf61TfQSaOv19c6fgXNzk/L4qm2EahuD4SkQXjJ295aoQEY5JYTVEahb9i711a2A
zTvaKfPw+X4BKQvDhHQfJ0ph7LYhXXTV+v2upuLygYFsp/V+J4av4xn50MXz0XGEkF1H9TqYAf5E
viTUsV84eaPMqAHMA9PuQFY9Qxcm02bG+odWc0wisE9Nlz1dodZP58c/k+BXi3UPw4qChXzTJF/I
UB0N98CJ8J4IStu4nu89gJcw3c0hKC06hmN6x89wAfPnUcQDfeVedQ+pZsSrKIy3w6uADvcqvjEY
ZHf3PQBrAe1Y0LtkLYjgDiC5lIVy292i2OxL4hCAeHAr3I8ff10qucmWZPe8AGCFz0aAc04Sf3kd
hSwQuz8kEbgkZ7dENO9klD4PSZ8gXctm4A3CuXdgADOMRM6PwFq5ZHA2sF/2+uxnpbpWI9e1JiAI
pvUo1RFOm9/4RfhoHVePP1YmNjug2tkn2ISSgq/dllsMLZxngUXWjUU5aw/Iv2rubxq/gVoefXZ2
agdikNmWmEk+WQuUe202sW9abnpHNo/aMPtoWiJ5WXKEyEoUlMXwDaW8kwUCsBOTdEmUAvR1zk6H
JyrXZnRLXrZ8i6YTLj1QTNGU0R7Bqr/CmSocwKuZAISdfGzHwNm6/Ofsv8avBZjv0QgY60CZQCnl
dLjSiK2t7WgXKOj+0NYCW68614mCY2p0jw2iZdBv2X9HFLhZq0oP5YyViHjPG6lFtWqvaWeP1TVP
jpQkwjFeF7aYzVfnOLKZO+ZwHr2Kj7235caf5YKsEaNJ7qDzWT3fPo3EG3uMjFh27ekEBvqjlrH3
O8UMvAM0uCdwVKoank0kn12ArMO/7+qABt6ZX00RBhWV6FKXxa+wmSiwMWyTjfskkF/3NiAbF7Fl
AOr9BW7GcdQMGaArpqFrPd4nA8EtlrF09EMsbgtFYiWumRx9Tu6TXLk4VIRe1FnW09HNSRZ7rLT9
5oEZchzRFyjd/JI5+cdMaqJaqMwZ2aLifnWMitytKDhpabiTeJX2U9pG7T1z3inpCaklenABbn/C
lFf9r4qA9ahFVujnbn9RFMBH/hlD5VbK3h3GmipFiJUjvZKk8B9rhVJYW8eqAGJUpUpROgKFpKm6
kVSHRMXWmBsBwHn4EHeF6wp7Ab7RRhsvmcHu5WAv48N/N7gmVaA9G6lxL2lsUf1K35MuUatduMLB
IgzONn4thVRR0ep4UlAt7dg+L/b4NLet8te0d+tVy02HOxXFJ75wng4gO0/A18xDuNJNStI0nug7
OPwiiCDJaEdJ+zC2RBffYyhQqFlOfd8Qavf1BuDvqEFCQjZwSFCAP+ozCdAzZnASkbtcN5xmR3Zw
QcOEPyOIT6jv/y0GUXheg8E1Y1PpPvCBmstJ36ev+h4VNhxwd1ZmzHbwFrMgN/3gnA1qC/loGTkW
idqNQkoymLvCB1Mra+VqdRRPjrtjyQG0smRv/+4ht0IeKodDbU7zz05mPGM8Rs5Q2wAJinQuhyJa
0Q+h4Jpu/QWQS4LuZw9+hCD4Svlr/6W6fAUVs2VLIWYa/Ab3mc05s107FqpJT157MhX0XDbd7opT
95t9iJT6l9YvzrsIpYREKsTRF2A1DRHN89BITuURHzkxaabSps6NlfglNX/xnR/RRzTpI6VL/DcC
auLIR/nPHG9i7YFOOzaEhvtmbTMKqG85t2uorLR+k5QIDxQlUEt7jn12YnSnmM+DrN11yypr/hNM
5zMw4hmrWpulLJSr8dEaNO37WfN/p0P7xEfPIpNW5HGGViKLK9Ys1sUjIp2HWfFykPyd5XG4LZeC
n9dVDta3u23tFHkCjWqpF3RCXaPZYxiYoHFOUpajU1SmMZ31rYkcyCyf4oZsyeIrDTP/C6lMalsw
lHV2CGzLBlFs1p7Un1GFVufJhUSXoJoZaRYunIZypR/mfR5oHAT1vxdyqaSnz5sHNXYB0QcLln5P
hF0l2SfyW+FJGsdeh7ox2iomYFNCZPfGNsCOMKo2SEtc02xf0y9uDKRWgwAvPGBcEGjnBLlsD3B2
eZq2Bl4Nwt/TZarirWrKb6F/z0fFrTxIF58KvsLcp2VXcPYn5fDhyn8vBhi8St8o0PnDhW5JE4FH
MNbSltSFKWExQ/2ONkSJbQ3M2Nb3zPsMQBDrGb1h6fQQm726V4KJ3ghcDqsiCCOUd3KctbG1n5r9
o0EW8xKtztH8gFUvtPLXF6NnJHbVUqim9ismSE9T40y9PuDILvO9fsE1JF3CTbigNlt3Vv2ep2bG
+gJxvGurXR48BtXbCccfJgk/rrCk9w/BpYtn1gip3atQ7kN2ihoUGTvaiEaAgJOwklWOyaQktqr9
nh6mjbIvqNCzkzoORhsVSWpxVw4pvlSHIL0w6lWhwHyiG8IvNaLudf/jI7I4udSK7B1hA//LBbYC
ZbvEAF7x/yGL9N6jePLesPUtcZpO8ag6W9qpMD5tL+UDZWB+q/CxJ9avNVSoMzHZuqGNwbKxTMko
m6nEgiS+RPfqnkWWFRGNYSLR8luL2fwEZLXVg130Gkx37Vrad4h+Un+BGa1pijypk97QD/WjlACK
ewQ02+NhzYYkMfY1IRg7/Th19iQ7kSU2z0KpU7aROd4c+2yG9H6IHfGHuZ1nJ9q+drKEOVr4lLZK
pdK/pYns2whi/YiA/VBPJPWWGZA3D8drHjB7GbnJt952xR1mrX1/7105GCeSgE1CXGop0uJwW7gW
n6CpCXgzHYyDxhCNvWDc0NQ5mCzWMDfppkf4nup4W4ex5puQ8HOtv/S2RP1oXzVrKCcdrq59uQTJ
u6pIGEfkShARVm2utHJzl1oqeZ1F4CAJOl6KqdVJrOmNF5HVduDdH8cnAeK6A0vilkAEXHH+1+pn
gLJimLQnUFGMAzEVooY4+KfkHbpARLjcJvGnrvW+AlBhCPCy7WDpmogw0o+ySEFg579zFKxdK/58
sefgXkIyr8JbMZ/ATXF5aRZOYNYOJpeKFiA9jyZrm0cfQzVRYjdIHIZpEucierFQI74jhLdQvtK+
HOTMxaJuWVIVMB1P9cPh+svNAd50Uyv1ecmGSnthQa8HANx+XaCiU5P4/U8bOWubpYlKTO/Dafi0
XqmTDjDlxxrxI8qx5J7wM8VfbhHbB7AhBw9MNQIOJO4pzA2Kx2iY/NUOFGUeJZ8LxECvHPfV2R9c
Y9r2Sx0RZD3SMMYmswR6GpdsoOgRUxkRaH2Eu9QnT+/Jz0puYK7kkfn57cFQx9zZ1+Yqqu1M6mgj
hCz2PXn3Xd1DyTj6RMARte8xTWqXFRVWzE5pPGZ/kpDE/fSlCOFqxTd6eQhw7hOpp8FrKGE9z/v6
OPT+RAlXL6gkP9oJfRaWQufFxmZ0nUZkOGczR6QrmfFfMm+66wy3uYmL23XOQ51wGMz7fX8V5gLI
NwTYhYU3sSMA2Fq8psyZ/T8+XW1yMtIX9691L5tbLPd0eeJKogK5Cqg0XAypO7y+cumtRcvkZR5k
naQwM6zknbAzOgxdlVNUYjSDyQgCCvtQ+6picv6liGRv4wXjYOtmw3vDcf5wfT+mYUuAkJQ5fNSl
FFN5bQ73QEZZhtOkxSs1RqV4NXyDIYWJ84Aikf1LrA4d52/A9DxpGZ5soNmxnJJlpasqM7dkY9cs
ziR4f+o5m2mJeaVco0P0D2dF3Nrv+avGc1p6F5PUlVRU2twisdPzw9YQKPMMx8vwOwx+ZCYXelmH
8r35t39ngEO9+/RW9apn7d/EuozWjNnTh/UP1rti6SomB4hH+OIiYStubQZEYzleDjWzBQKYT3yf
HVgP+qVNd83RXvfHZtLBwlaQWEFhvTuOSk4ymWvQYYf0Jgi90VWQByF9Yj846lk3EEeQBC3IXLYV
bUlXthkbgLUpFnzer1N6bKdrqNLM2+NDOgdvZVbqa2KJVduKUaYAErfCRtpvq0PbUGI5RFKhz2Z1
lZIj9MQyC0hnrpGq13oy/K+7u8Anah0vCrUEvS2/RHObiAKKUaNBvGB8JmJdKfNe/83uE+8hZ7GT
KOzg4h0/61uw3+OIuFbSFj0bD32Hg4O3wpD9vl9ARx6cKNdnA3mVKA7zcR84RuzoMfVVLLetwhPi
upCEg+hP9CzMz7HH7Kd+z8wPbjwM3orgkc7FwapKeK5lbsg5rHyjs2fjf+zPdl1sLa6lS0TSOMPv
37fVKhixrl2945t2+sj+KDjiHLQOOVVU4lsEYE+vLQ5LzuqXIrbBzPNJfI2T9VJAYqv2kWPKqfSy
6+ekwcVOeIDjwf0igOJQ4TKYCoETRfANcdrsUg5dL9YcCHQnz8xbFsZpXuQHboh7Y+5cOzQeg4i+
W+41W1fgM6ZFkbcqkibey4KCCKmFGdgJIPDiRhFfHtSFLcg7cM13KZo/sKKbGekecBgsHFaZ1F8z
UW5bX7ADZtAYQxgun3upJcEZtO16S2c3lmiEd+aGeldDmGhi5zniNE5jUeXG08Li3LAlszpS489K
h9Qqbe2t4lG2iOFKdkuLWxzLpSrWTEkYkBP/IQfRmN2QXUMncVEavOZ0IA4XAL81uevdYfIGfdgj
ImKiqacPG83ku4lFMp66cp9mTqVwoqHplG7YONpuNqH1gpCgLVKDYJHUznT0oBQnZEfW9mxRuFrC
pzfAajOmyOQQ6zfWsjIRdGhQjYd5D/VbVoJQ/IoR3uIZuvp0cphjEJOwd5FIlQzK3EkqCJgIHe6d
ywFudK1tMHXWCd+U/SLBfnd5GpyKVRD8PLZPCW/5Mw8exD5UIMeAZby5MYuQr7Y3ywgSlHmdwcny
zV1OABqwKjyVVmU4AILA+cqmakzd3IAkKZxI955YHIpv3bYgOSDn+k1qFPGR2w7qj2dGhCDnOqjS
sDbuYp/QZ3G6kuYvDiDkELd6sxuhVArvKMdhglB1GT5CtLQkcQk1EWRNLcmgU0BXQNesm/A2j3Sd
ybVE4c9hUpvK+0druwuVQiFR/JkbQBnBG8ix7QN6CjOm0hQz24J+mmcwnSmPijhI/0HtPtsm7k4s
RPVqcmN/MNIQPXUR+7Lr/mx8flGTg+u/C784K/nu78aNUVZpBDK/L1nQwxHvYaFvAJm5V9s5fDLk
e6Mh7790mUD9uT8dYY7Df5GNYVS+IxfH6JiYm/YraOnmM7vwqKG3h1r7g/i4UTmD8A0fDaw5OdwB
IQvSV91EEQOK6thHF2ChQfgPzS9+rEt8AkZCVfsNHPth/TsgqqPF+z6InqPlyjlPhjinyj5tM/CV
DQA0qIrZH5oYHbEbufWDK82UQfjmoHSJK7XHUNTSidjAeb/k19p4jxVKni1GMWb6f8eE8YV2f47w
UHVfSsv2E1pvBWqa2YuIWmEGxPmhH7w4Jt49kn99fFdMbKJlhV805LpZNkUD+B6JIbmzEHeI1bjE
bFGxQMmqWH36RBI5fub48wUATj4lIOnBxFWJ+fOyXfStU6QjJlijPZMwpgI89U9foKATmQ7CoNZf
AWORTCP73QlDPeTk6eJebxYc+o7DWzIlFanBGNya3dhPfMrRJnpfUhsuK4+wHsxJyb51rmcyMVna
HZO0oo4GVfd9K5JJItIo7hihE0hW6xGlJP/XPqPKMMxV1NeatCp4WkqoPUXhn7/FsgjnFB9wAVDP
45Zn+K3ySPBUWGjya0eSB0lvwelrLFKErMX57beaNhUYOi/lLnM/hO8OkJ8gihpQjhu6x2Rkd/2X
mKbxknsU4xMACFKxJNRbduGkdf+U+7bo2O08cIUcIRnPoD5pZgj0I8WRsoLMtvduzi6Npts9cTN7
gWtHYHtXMiAxgUcTzy6NZUReoPzIri0cT5xn93pgqm4c4pwIuj85fzgiWiDtjEGo4l0raoIvRkAs
Zki/spSJ3QnWDj948Jxye5YELe2pvnBRawQvqLdUwGScet/JkFiLaV+yqLnLRryHUWFPPePDFPDt
RQ4fCEzfv2vitSqOBIBfZJdaNwIgyZ/IKv8SzoQh85HEIJsAzP53Li3El0+eKFqjnvDEHZCgr0Lc
qvI4Q1d1VygUhrT86YsigZ+EyS1Osinl2UNGD7Tn6dfelHcRBSuSSFK9L+PqmbyPAFlfEYPYZbRE
aAa/niTfetFPy61SG9tsD32Rguk7+aZQg4YgApoBaGITTXgKrSx1jH2G9PZ2KPChIJg4ngZoOCvO
U5mjJzqLwDz6iIbZU9FdZzmUFrmz/Wb1+q97IKm0oWj/uM3MCxFTyX89MoUm9eLN4ZjQs4htlQCr
AH7te9O1pSkQ1m1v+rOyZrRVGsLnXUYwq+gQimnchQfPPlJkKw4en31nje6W/FqbdO7DaMr+bh3P
WnbncLOM4ZxhZlqT2BE/4BYkTj+bYUwuSW4kfQR+Mj39HPMyKybWgl0PdzWrxskgx3psjf32V4RM
dUqN2+Gz1sQPe2x2rLf32/F/m0oHIojao+xg+fYvIwMhHlezLJipyXcnUwu8IPatUMR+NJmSvu1A
FydSOLSZYwGfuWNBfwg5l6oznbJybkoLEbB3i7qExwGJdO/uO4W9UV/T8tKDMkUyWDz8SsjvAak8
/wflZ+zhUoV4kxxC+wN620aQybJv8PinHteZyF2NXRaHK/rXq/YmsOWx41OjF5RsrOBST8fpXimt
ORSsG7TUnmCDWxK7PxhSvICB33dd0Wdti5jYk3SdjyKP/ANbVGbZewt3vPHyQqH87eNS5/S6mSKb
cuMBrow/SN+iekN7qXL42dHnesiECGADuOUkejovEWpMU90n7rD5XR/pMBCEe2VnqtuQCopTGkyy
Cw7cOAT2GCKr84WEtWRfeKJ0Y7U3gKTJyR6vm0RSI7Gd9aA7cIkqZZuy0/lf1kjXGzCIlLFNlJu7
29WA1/gZ59b5bEiSvncbIOYwRR6F+YnMrip6Vs/QzSQnBUs/NtrAKXXNWIh8beIfWbz9Fi62pkPC
cawvC5DBN1iPDAW5jvFlOlqee+KJywXc4/SPw1CAEvL96x5lyev2M+T3k/xuGzPCmg1KFkxyY/wJ
PbErosCJebSmswarAp37WkWpnFqVq7u/v0y8g6usk5JMgptRIsCVTq562hkhNstXd+q/Uhjt3PyE
cD7LFtHR/zAdAxaBKMpFQZUPIQvlKI57DnSwlQ45s6IOGBJdihC7+O7CHdaWaP6Fsdhxgjzvzr3q
9f5709cj4psCRTCaniLkQy5C7OisUqqeWjHVTxUSyAD7pjixOOwWIqitm8xKNtyyWmn+K0K7BZZR
MARlOWGzIz768yAHEIOKzde795fDFOm3KBui6My/CH5q8hlzzNKCmkn6J+8Cum+9lHjEQ+tPzkhm
5dsMeG17ZTrWs6sfrq6884N2NrgBsXXqxr8LMzki7egndhMCOe41NbecoW59dm1CP4sgFMqZ130F
DrfDCBKPcw27tb06noXGNCnQX/0GenoU0yNAJqbcHsN9nnS0WhL2QPO/+UQT+cdSWQAnkI4bRZU6
TAMuf2OiogLJWkT3RictetawzljfOfOk/aUhGgkBgD2ArPS6uV2vJ7OiRRT8m+20qzELy1Kdnj9R
amew0ji/wwvutrN7ldfmEQaLpRGtgVRyeTLfCJrJESqfVxbEpp38s0L7rBySUaOLzQhpFac2BPES
VWvEiC7IHjs1tJN9A53bFArmK3OGeQAKskB7DoT15vHle8OWQ4h9SDfTcdbdfoDcFuIo45ejEdK+
7accAwPxF2eWp4Q6iYzTBenOboCRVgn1vs2bJlOf5XELHtcyCeyJkNJ9Da0q9yT0sXPkkmXT6iOy
vZCBymVQ+Nkdt+R03H3wUSeuSlBWA8yJTpyLjcwuVsp8WqIS8qMrj/sNtR7cM9onX7CC8QtReXcc
eXUJHIofnJ8lHh/yrGp5KfRlMUdd4HU5DDh6CUy3LpAbAb08JzxJFp+cy4imWH2g4ChkDTImTRpk
Nocggdwu0uNZc304kKbhJRnbgengdLY3ubdjIwstBm8jLtaMT67rb7gcHNsrXgXfZelnlhRneXXj
+8+/9AIMW2uIgXlPnUAnVPH/7pAXqQK/MGnv4XAa2q37KQf6V6z5BY0g3AhT1zP/CatT8mIIkpPp
Z+1b6/VwlCR1SyJeFC3BZSL4THVDK7lX+UU0PbZ005QtlGML9hye6bPVG2ItJZp6TrCB5eKoz4jI
uKW196wsZQq8Gj0oY03tfBikqfkLvZy04CGitbTLBSeiVW3Yr3hJYnuLN2iw+5ozE6KQMcOxLm6n
kpM6eLMHVwtD6h24eTrbkjhoCU6YjTHauaicnfzoonjMONewbkj8FUXqHjcw8FEgos+IUzHMFhrN
/F/NceEVjaCAwjA661BeUw/sbzffF6kGw0B3053PedG52ikOkLU0vznnhP75mlhGaVGQBnn76Dp5
VwbhiM73BMGaUDHe3AiDTKpFfBGdDb0ekzyEW7ExPJcQ71v1YU0k808D+kGcXmocrwLfPU4a2TuG
mITOlLXLHsjq0sjJyOvk0cayEHRFPII9JLfmLYz9Mc0OEyQxRABy+uiFmMdpzrPAGd5JlAZaMVZB
w3h8RoZTFScaTM2qpaoS7k6qI4zXIkxMDbSuDA0SeQ9r59onCkLbZU1atI+9MFiY5uc5BsXCms2/
llYko3XsPnnbsBlGuVk/ss4CwDbOYdhohfFe+bQyPKiUdtXmL8zJUw9CBmgZP2WXiQjmsFF2jL2g
jawidUphF3kIUm4S0Jzhytf8okirB5OlNvHzlTbau9g/qhiV/8JBo9GjiOz+FLEDi9BsTCIHzRzf
kRSsA1tQuy//NKlqDGF++tbVPzl677XVrjtJvroLa6D+z620V5QWzTShivOOfaI75xaVtMHEptVf
SRVYf6nHCy/6Eb/BsnDbmAOufCfNdr9C9pbf3q52Kh4eayHhv0yJsrP70ACAsE0fQv+5SyonnRos
5ISrH2nCXNb9R6bz2z/+JGv4vzAYrXUhtXltio0Tuen09uMbUzWswbaVR8WJfZMwAgYyovIfrkWr
wM742z8WojtxyZOTN+xHLjOdAO42sHo4N0rYwH0qMElpY+eq1MD7s4cMN90ZJEwlIXUQDr8XXgBA
DoZfDBvsAOaed8JFLqueTwVEOXSjK28YC2EggpRRcPLCnjL7xUp+h/Fr1ZykeMUs4JUxQKD4YfWC
U6Ts7AGl/041FGb7tqQhv70xFO8WAqE68jkVJ+uXLdhT3plG6IhnWx3O3J5g1Txii3o77MHZUrlO
iKOn9CKb/bAUpl/I302pVh7Z4Z776QN4hnb/ERQ3I1Cwp+KPtbJC2vEDgAIiMOWuDYoj68KVvb9k
wi09S/NgdeWcqRQFCWiXmOuMoDrs6cPDcqzfG0UlJFTVUN9UyRbgaK56QNJ3KM8jRuHMAxcXzkQx
kztegkteTVCucgjMDNcbfTHBJAmYmeUVojeshwDoVZVd8xT4+ss9cmbg4EFz38JEi7CHW1adNH8Z
l7ie6JhZVFXRmNGH5zjBYHQS1pYkedZJqpOJipijo/C3KNdSjuC4bmgu+fj/8p/JOfz7DYlpYyxV
uL/VUcrNsa7q7kZd9kJ5CmTqN8rS33Ze+BWwW6mKIjNRNqnIO/4dB/HfSHjMlVTh/ttId/1O0ybq
AHWrIJDC9A3AxIfvhWLUAwewUPEyjdW+L/jtE/p5xfuoC4aJuV41nio8sUJkfhq9h3V/cmjqyfeC
cpRwpOASTKYpaGxbivSEwEj2seE95ooQsHHHctrK5ZK1oNEhShBIYzXBUh6Jl56tiv9VxLAc8KMC
C+uLkTFt358DgJZ3j5DXPgQ6Zxe1DyGprgwYUDklYpNc7kx+glm/x4x5DgdH6iwHKH+BRPZSjLcc
IyynJ/92aYGgmVVRLnYHAGxWv+hcwliDxV5zWLSRBzO2m/X78MR095sFUCKlsuXKlpj3QzmoAAKz
58A9+Gj9ySpGgAb09LGcn5sl5XjFYX6B8hFYIhilRyDlLhL5N6k5aYNG8OL4zawmdNTIW+LJmPRJ
YoJM0XuC3wqpqT2ks4S0k0xVr+8Fxaq2aOplX3uKPSe5E3lwY3SH5sjk3NFoi3rU8fYdVgm/xoKh
3vVdbwQnIvQBBds9FWI5XoONQ23o+/9ua24N2hXS2lOwu6q9xg6HuuR/fZCbHKmIjICWTqLSdqv6
P4jn/EcfdOe3MmxSNK8Dr7JEvyCzTtqdb8mbqLfKOB0Bxgv0NiQAerIFId9qhepUI0vynzoAiVY7
qUpR2DayW60n14xmYAbJXpd0ngBCkPku7wunNvu3mtcSaF3tE4gl/ap3qnLAO5NbfMYM8B61Lzhr
+C5iuVoByd53th5lna233DnwNIarCc5QXovKgPMt5kWMStCbbMX0i1f313vkzJau8Ym/2oNV+2h1
yvMBBJUq1pxVAtPuIKKcUfDU8aP4IrvuxCq2wsUR6BGUBD0UW8Q3tiOqg0jiqjZh9ZeBmk4Lra7e
rM9NaWZiWTEO12RLwQa1W+fznDx9zZoHONdb3Kk1cx9LlmI+UQZonYkfivX1VZP4jmN2sFqzweUl
PgMqZTalHzXTc/mFNn7pc3p7RYu6g/IQxPXMAZaQCpssZoJZEQyyem4prnnkM2yg4JhHpH3hFzXA
QIvNfI5f61XCsW1mHJINuSwu3Sll6BoC0+/yosxM0VQQMAFLQM5jQ/fRhTEha+Pllxowpd5a32Sz
j+h4JBf+bt9ZFS/zMD6UAa/xyVgtkGlBp4Qq2Rl8U8B+QQ1ErtbWp4+yFhiAoeannmZTXsh6JQzu
HNFdBru4SJU4Sy1c+WS2ucighXvFYue6PdD1jBBOR/i9AjQHBB1eHLBAkXzLWSsDFHOOpSxj/QCj
n1L6pjYg5ynaXgtuyqGnvjupHWOHt5iTrVQM+GrJFP4YhIjURdvpbNZokl6J2rgy3y61gChbYOjY
wVgpH3OIyi3Y5jOI2MNregVIGKG24BPNr0YDJgAvK3U8G/adNORz5n9raL8KNZjISD2dfS+AlX1G
MDMzt08DzoelLH+c3fkqIAIiS+WBCfSGtzs3E4lnDMRQo50BHr6e3N6vZFwvIJauPJWB+pHvU69b
/3yluiT28GG1v0JVHbMUyGEOk7poHk84SClY0ZZV6uopMWGuZfOWDMnZb78Jbh2jELwesHyS/yff
a+b6+pc+mmbzbzmfTizcsbi0+zHyx8LwgtTshKWGJnauS2pCXZcDD+qltVBwqtfaJD+73FtkdrIr
0UicoucbhGKPndyMVLvUH6l5aWSArlt3la5N2bI5j0vt2CMvTW/i4xPILVObxRqvHFVLcav1FnPG
el3+cZFVXhSidxH7dCP2hY5dCF/98/k1igIv7Bb8CBqfEPlC3Wzzrs/ndXKgO2VV6PkL9G9W6A85
JRtpqHVX7/luwPcSPHJ6Nig35XShJUUvdmA8+nay2ZadEYmaDAIEgSW1lo3lzHhKTOsHt3TBUrtS
Qt5AuzQMujWQFw/rhbgnNA2uzHgiFbhoz6yuHlZCPlN4HYXLhe+EvvDhyOQW0z0pMsnOAkWXo3UO
hVHiiZwhvIARtkqbeFxZLv/4CESUOMNxQaBua9/hlaZVal4jbkC3ETbkOBViqPCN6gSsUZXeh8yg
jEKMmykvvMXWAzR2HFVIpK5hevyFMTr5HCo+yrq9tqM9jK1cGEkn+N3WYglAGTwB8Sgl9IgVNJc5
/iR/UKjytvpIvSzLL3P1xgpUTwp+NiSCnmkPnO51Hl8N4SJljcp9X1YmL+kGqoNNLKyRJSHoX4hx
xqI+vUTI9VXMe2F6y/PJAIUDdF8hOFGO5NOcVL6cJdWfeF8bsrJ79DpKMhBYV40Cvk3khwkcT5zw
Da1kTbO3AXWCMYs0Ty2Cl2UVpRGdRgBAVfz6jAMVX5MoeKsreXOiiguYy1f+QGw3QQ3rIEe3o3O4
3ssVR16mc9mgJ22HC016bFLoD2Svg14ELhC7qAm+eAMGiLd+X6gdvd4MIH6o+9yNkOazecUTQgTo
FfYfWornZXaVsIBNlwOQTtHWNzaidQXwqS4GoV8n6SHq/V8qEW8npt7sLm2dw0eJm0BFVGndRjiB
hfeodBKVfeAlp4Vt3JlvPbj3mVoIAPcrCam9wQdbpFd9Zr7RhcVgmMvg1H4asYy1YX6/8i5B5Z7l
sf6PW59Bkuj/9qH5/g85K1CGivWi27m0gsrIPw/d9xiXErLBiTe1ULjU2J39F0mJQADgo131GgX4
gTXvV67zhI7IR06qoznUYUgaHNT9NuMBHFqhQGqPkQy/CEA94a1z33c7yzrZttTNn55fQZcL1Yt6
lspnIycTnKTfLg2RAQv48r8Nf5Y1g9X97ZMjmSj/bVNQw9spOtq2KDu5qE/K5nLBJhA1+UYNl5FV
8n4CAY8tRqgjn9f1qZLCEyzdMm8i6HaRjR0n1g5mJ4XbyrrqhKE3aNYPW1y3xuIHZJnVHSLIkzJF
2eCn5jwTx1QbuEnXNpID0eXrjaBHKBy/IByzShAJIB0wDo+bTMf23j4K8g9CfEul6M+/l3bNS1Hs
B0ouCho0Z4k4jXjSP7VZPE3lukZwAg48SdcmhEF59RsiQI7UIvIjDfQw36XP4ljcmS7TNAhbF0It
GjBLNd2cv2hbSfKZNYoO22kwJztGqQd2NLN3KAUOKxoetF/tUHbiV7LNrmBxD8IOEFNAjvhbgqPU
rJyjVvoKoIw7QQkoKTS1/6en9cHOk1LHoPCfSvfckLpGHKyUt4wAY7QdX/7gp9n1HDgjCZ9BPpXH
pKLJhEiXbxPAaaIzPcYxVYmhJVSlAkCNWkMdoSAfFmjfwUqvBnhqv8eh6eumv4N1YxJAWvmNyk7I
mMVYa0s5HWuT8SAc1s9BhXmzDN4t65Mzy1BTyMpJmWi2Y4r5vJI0f4HfmzaI1jf7dXGDFg89vux2
7TTv58lbZquNaF3k4GDU69Kr4LlIMrX7Z9S9Mg89pFwnGYKZzWGkoveSCw3IakdUKJFJjsqTwik0
b0Qkyaj62iEQ49TNi++fTpnQmvAW2scVEPWknxLFWa/JySwW/c6j16zOTrNuD5/etRsIz8ugWgvm
FOPQs7iQpPKnVt7TPUeHvVb8KqV5k/QstEEXxRqRHvgOBihKb49jAkiLlKRcPO82YM9PibyKMEe3
1NVl24LFcOtS/axuQaWzzr9iI93uBZofZpPRxTKEsUyDfulSxrTGYa99Mdh7Bafli8gOnopN/9BR
v1ZOEVo98z8hO+/dojd042/Jedc/pwZjKg9SCEMaAZYwXD9VtOWlDMtJuwzkA92OVgZY/dRFyi4t
xy2cvTQCrAzM/g28OJ73J1S8KhDWRIJj0PYXHVFeDt6HCgR/ibI2pL16ZLjSfURKcbgWlGnhi0uv
OVNRbb3eaWa1QqG/6m5iuubc2iRO1rxSA230XA1wkouNfPK7HXNdotrBxbh3Z50PjG+cQqc+IfIp
a8gK9lqmvbpys3UIm6eXxdEOFUhCFwXbLRJyOP5U9Xnyx/vdmYvSsWpHowZXAsOWCCx647X5ulXb
uDgm5VibFB6XKFRSHVD0gnimThjHDdMJF2pjnWG+OEUiP9mh2fcdPtem0pBrfcfBdnFzwU95VL2G
/sCPC1lrZJDkBavSIBAOSJLK/Mo9eqmrtWZLDiZrZfdlHzNUfA+CHtCX6pqBLQQlV0UI1I1Az6fr
nHLr41wsQhBb51MV8s7MBBWP5tNT4DOcfP4BNg6Uj/bUpHYSBqqeaba4lP3wc872y5XY4qjpzPdP
wnRoxeQ/ZnTRMf5oIrTkA/s32ztepLbhJXdL6/IeEX3lGYBRqO1FIjcH/UmttmLN+Mq+sa2fC1lx
0hi9nE9WbCx7tlg/+pspfoJhy08TH3yrBr32zz3PDkzs3qiD0sWWBy5qD4VY1fF18A1sPo2UDqrc
vtFj4SYt9uAkiImRYoL2QOxeG7WFTwpacwp9awceeVh82R0+KH6BFRwyG+/DsBb2erMX5GrbN/Qg
uYfsgikh9LMMxwBPIrv+eGUyJn4HfhewuUYy/Nl0CgALpJ2a3Z3OMbDzmuM00UArsaxvEzCCJbwq
iZPzqBLef25G79y7uJjs0H4CrYUmGxqjDcvyoKuR8iFoe29cD7moXhYKwGVs+JhDNS19r5z5e5ZX
9lF/0Cp2iE00Zx66ilGmdYtmdkQHCmw+VHpnJXhNTp4VH6OhPunITUZLNnbEe1ThuFnFsSLbL7q9
AxEM6Da620Bhj2I/NcEbtPF9bHiSeRpUguGB3/tlg5YAoEq97tenLQRcvT76zWj9mRVyyvEMbEUB
app2voo/2Iem42h2TaXCaHFzU5Aeh82eCpmDDLxy7ZoO4Xy0zkzx92KzrA7yHZ3YWBS/e404X6Y3
coJsvO5lVIgDq9gSHyEA45PT/I+Fv8kVUwhYDwF768o7iGqItcQQ1fbgJZwa1J1oBe0ZUb7nKOX1
RVUjVrrwBkIaoMxXjXrGdLC9CtZL8x7MOOhTjp9N2SxcrFH2ygOoRY3taLQeusR+xEL1ObjETGbw
ohljQTEVVkbceTDOeo+/j2wWIiorGNHY8TOkPcsXa4paf+lk/BA+/A7Mffmr6qgs0uM+XH/Ld9AO
98RI0ThtzcDnaxZHd8mqsroQJokV6RXnNvS/cejAtRIjlXk1iUXPGzsZs1TzBNCuDi4HRgqdNdOf
lMNtHuOOwvKY3sLLhlnpfekzA0eoK+68RP/kN42E/DFuLFZXmIA/0depg4mPi25LLvov5okyRc10
BetA8CQsBoepfTJcQVN5Ky66KA1znao6n+cdVGOSyZmJme5rnXG7eOdtsJZOCBUD3UX4UGCy4bLu
2LwsyDCWFTABTkl8Mp6cVBYpf7iyhtfd2BRBkQrBEUAIY4YRcvl7Ohyvub6jWc0BH7RzdGzanOsG
V/BlFQMt7filRORJbus6o2u9Dwa/6PXnhGbQfNLv0BkiO6kwJRzRTmy3NyacOm/5pmcde6n68Ud6
hf/SZuPC0h9gWYh75Xb3krcVOAY/ECeC98zw3JHZiQohAmB8BgYgVv+X7ikttV3sXQSlsyWtWkiK
V0oeyM+TSDwoa44ux7wnnlNqPHbu7Qk+mMOpDG3cmeiFmSoVhU+z/Vru7G6L8Q7wNdx8epQkJ/Al
rtTA/fHg7BpiD6x5pm9FkZEQVzFTI79KUAKb08HYzkUMqoQ+zIxApW/m3Xl7OhYlEAM0VEpuCRGy
hMdqyy8anByt+Q8CvLV6kmiwP1ggM7fC9cJDqDmTZTXKJexFHBZELPyoSvpI9+iwZrZsptr/5UES
XlEItcUajc40OXbGXHUyB4F1GC5/km6a2PnYtTJHe50jWhHdup0Bjo9WIdm/chkKBUNJLC+mXt14
khA0N3ai4qKgKOjtNrBcV1BEENcgS9/fOfvvXNVeFmoDu0iFwwshP84D7UblGF1i0ugqaT/EcEqt
7AewGZQobIShCD2V/U+2RwSWaHwUobaa6z4zq9Faw3I7C0wTixF63UOo5Lh7F7ah7dTBm4rxiUV1
dBJCMR4z/Ui7pmq8oL76A/0znMtOlAMuLOwuSquBlzAmQl8hHv23/0FzRza1MGSxrVodQMDAOu3f
CgF8X1zEGGmLlXzJVuUY+1J+25b+fLhPb1rpwaBPipHSfouC9nEcmjJBDx9DcZtPntxfrEhUbndd
bl2rLhrKtTRfSBnEMX6SF05AT5AhE4OsmZ0lD4ysFaxmdPKJ7m/T2/sx4hwsx6fa/T0N06yu/6c1
O5xFtyrq3XqoXRtoMjrCdqPZuS0djtXT22/nDY6ZibqK6CpSWK52sE+Z6BlqMno6et61QiRhI42Z
arsFoa5jwADfk53G9r2acHnn7ivLNiR/3+Z5TlRoLk1QfJY0Je1t0bCDWYkiL6ie3MeL3u031fic
wpneovRsbh5pp+8JcWoOLX2hVRLE7cD/YttjCsX35wuXS6ksPvPvy9UrEZ+eNmZ61z96YN2XrlnS
M+c5h7gyRer9gBBKKafqamXdTMhx9kCImvDsye2Ygj8FGAhFClfR9KQuU7eqbrTICDPfgND9Dq6i
2BdcDWq/9doaxISo40naTy8f01VYZdlKlwjfXcHrylMjzs8EM5t1f4p0Kf2IxsQAbxvj7DAgsk17
OmO4gKsnGjdBwbhgpQMXUdtZ159M9OCc+KfVjJrhP7Yws/93jgUqxs6vHJT4kfiVYhKW1EElByHQ
2muYC/rHVWxxYJnFaXR2gBatOn/9aez3Qsmjku+ob5PM+KP3Y5CtfNPkewKQkofIrI1A5oc5p+tl
KXKVYKcUw4EUuGJyxIVtZwELHQ/a4gYXXSy9BEpPMF9pDzX2HfENWof+I78fcYUOxH8zdOB+jOa9
BBb3osCxKY/bWKYaewWDJer6Xzt2XAvSKV6K3k1JsTryrkHuL+DphTzpu1o2LjuGz9tnyoBzMlDb
Ce5RJYnRI7WHwQR+80TW5Bd9zyi61A+vw7R5582xlhdjXcQ/PiYocLPNFYKawyHW6E2AU/TgxozQ
pV7473OVEK6M9L+qbfTV6Pb7ts99ORIDz0mr+pdN4w7IJTvpM2mhkIZA2iw/Qm0yW36/2YvL7VYu
iwM75OxZh6D4/XFrW6/QRPBnkjEU2m5LZ6o8++4DOf1tNu1RkDJaC3y7GUoskPSM8DZm2qmBonel
pXShfQkKr4h3oh21go9MAtr/yTIMbRdyeyEW6nH4m20ADFy9BMR/vMPfquwQkKTPnwNmHJJlZ7QC
m2Qj/aOMwQ5p5efDILZ/WqgtUYYXJLE2hmcXBWcl1v1RkFQv5IrsWhYiQ9TwjvbJ/GNZ3cJRVh0U
aBwbyN1fgII/BIMfp1dgUWEOSWTOEI+tcc/4Vx3rVA7r0X9W9bXGvDdu7BBoTuyFMsoAbQXalaxA
VgCqDeo4bwaH1VDP4DA3SvZ/Rhb+HxfB9UdUeTV0bVYsktaAghzMFT4ssGBiP9u4g0KzQGsvkLZn
SDceGgm6uY1SDo/Dhd7SOu2+yJrjL5jckOtQh088eyuyoJ5NxE5S+oUyPIPhQuGaSW6jO8dCDMDm
LICw3RSEkJzaHIFQo1hGcPimGxAg7KLkMOStTNrI4ywIyDRT2xm0cqmHCkLhAMRhDWQdErL+EDEe
gE6LsaIEggJ/Eiz77Hkal3YO/+aVjXw+kBTneD0PR5ZnRzjkmejfbUwoQWsVXiAl04VX76Zow8bv
wjnAED/ufRpa7bS5Ch4ipKDxr9LTvzF2sC837/MiFAngF6DnJ7dcmbC2qulDxAPl8fWOCQXkpUEg
Bpo3vSiiZLZnXrCUab40Xv0X1B6V5wPxzJysUPqFgIoZP8h7k4p6pE2WweoIJnOvZGia4qR1iL4S
ygZNRZ+me6WIotwwt35iAmtbkosCUHUnG6KifUz4L96nQrAFKzrpPpIzfzY1KbnIx3SIdwhD/8a9
gjGMKJ6fd0CCiJlE0eM5F/LxvePMML0uSa9Pf5S3AcFnYBoMWloPh7IgNq0ZbNXkFbF0EAS7ixDw
Url8JUjkk6hanFJLWJZLf0HJ28civPWVX5KCHHKWW4XyaHt+FzsiCHlfVk2V50AofPE1ioeWYWJf
i1ZAnKIjklIwIP7R+XXZ5vuoAP1nalFE9BFDHjioATvYjhOCdH1SiwDjNR+kaPyNUBOqXcpIrZ9y
hHbNy7ccQJwfdOfk5DHmmnAVOarRttGBxvcHF+gUB5zAe17aR39NycDjXUlQHNuhZu47eIempe80
h3iIq2ohyM5vJx+PgdmPsT/e9Zq/6OBx6K4ootuhjHufzxPv29L88CN/3Mwt+wSPJPZk0XmplpID
ojQTPgN7k2yXQyPFp0gNmErd7rSLmKuVS1B7dlSYImT9sw7/WwKYBjfxikdk1ACkhc62/lDFLVA7
BDzM1uBj+wW4yjDe/Y0+s74c+tmRHNYgNf0N1wPeGdAYpUuSUWSDHcYf9sRbBNirDBPXf/lRZ4pE
LQ0puARdVGZOyaQzxEeVLafWTz8XREPNWijGlQQ5VzmQRLI1pgsr//4x0MGtcnsQH1tGBtlF+gN6
VBG3wXRTiGLACM0wZTHCd0XH2Vog0ZiS9RWjKrVhuBeMdmcilwunArf351IBUmEa2wJDkIcAUDwY
+XlidZc4Gc/AxpRBLYPEg0ukktsYz30nU3CKMFEW7uDOMxpBzFwskj61bYgau3yhQj2MACqeRyJX
ItU6ZhYCjymttHEPF8/kUh3/hqVxaYB3qxOHo3MaJANvH5bwuU6vI0KpPhjjNq+YOpoRvQREUqT3
+Uw7Md3eIi1WZu6xbqGgkDIaoHOCXq7S0dKXIEda6e2/uWrShUeMZ7YNEn0gIqzPhVrjo1WZTR5I
P+h+3Vyg1TVOKxZw82mPW2rdG0uuXYY2Ugr9MAnI6BkKJ0bLdn5W8Xqu+n6qavkPipe5Xog6RWFU
Xv2VyO6SI4/wVkCPqEz2MsxiMuVVjFhJskxZxOvXXW62WM8S6vuXQnnt+CDK+SC48+gnKCSgXvu0
PItdjJc3thkETXqtoGAOegVaintgnoNb0jHka2D1/Nu+IGGimbiWxwS8+iHPRpPHuQy0KgyrRJj2
sTHntjWwy7wHd65zVlghr6uI07JrXUKEm5SJ16Ej0kDC6WpabP/qyL0xzYbqAwj3e8kmFrAgtaV3
mYF29IA4h/0A2e1VU5aO/4fzfoOix58EKTRlCys8sKK4TdPuSRZ3m7X/D7Z+l75AGmOBnqFG77TC
KDJhG4/c39id3clBp45gVgLbHNHGtEMqjqx9RAJK74YmQAfelF/4zNKvY+p9Jxr1Q0Gpm5tvbsPp
NlC+UBw0BBmbGSa0NLX+CLi4bkqSuSM7lXlowO8OsbVDOCbQOA7XhivrbCZ5LI/MHdBFLcmKFBJ9
/tlEwgyo6E4cezsPlNSsaUxJQXU7t04zMycs4uYIPUNsu3sWfVNULHOsqZoU17mdfVEm4Irj6bZj
cKZRPwTlhxwJvJOCSG/esi85VuE/XFbsQFMKb6c9xFzuIaUy9w3arbnQjNgH6n1+mHWR/B63/w+8
+diKMr8s5oxLmYDAcxTGKlbqjXOhJRZT/1KcZSwrTSNgO9+bpakCblVZEsVI+ZB2UYJRNvqUAR8D
rehl8I20D0U6PAOe6fTicvZ0l2PlUKvSiVpX+ezaNbLLE4ldrFWtKSX+MzES3VsLLTk5IUD+3BO9
ItvZAkoiCv6FvXc9Yf2L9o/A4WdikI3JR9LYCCkIkxtYJIZRhMfMc3d2WjC62jaA/EovcLfa6ONK
l/W+3GYFEfOQAGQj9FQzWL4ahquD+fcYqTH13YtxKeo0gZZU54pjupvpsDmasV0FUl9BZkXwlM+k
zYywkiiGsPL66doSPObZ27k6F+MVBHDXEp2Qlbm6I0Sad3ohqb841hbJhR76GA8Q7lL6yieDbh/d
EuAugWmG1ywto7030QegYn75IAECD1ERmEq0RguHsef7mSQmlgFZT7EEBgEFOMMYkDqNmS+u0zPR
2EK8vK8oLOrNqzsxihTl+T8KiCEhil4wOdH9dsSLsgJd7gZ/lypEHfehKilr5cgHHpVkcIhdWNAb
OPJm7VD/2muaAPXfI7PrfABOydsMjIy1U/85tWdMQQJkJLdOhSpoGmBqL9ywCTz9La9unyiWKkr7
9gz6NRwnLMoILgAhhJb1SJ/+EZ5G51yn+y/hk02y4VBqNqtroSNKuiqxoqN6bShjpeW182mcYfnX
Lrix66UM0mrRFQUjfAENsNs/vitI5oL3e2BhKIAkF1fzMBEfYB6os6VKehLQ3ba78utohSoN/Ef6
f+6BiqxWAK9mvzdoQcYK33IZZd+y/n6reU6cCiCC9RXxkZhpr4vzEPfT7HZEJVEhATMYs36krlYw
N41ZH75XBOJVbhax76OixWmgDe6OF6Wo60QmrHYcb74CN4I3oLMYBQx1JKT6OIAAV9cBngr4HPu1
CiZIFxK0BRKgR73EyZaCKLyTNYRNmFED7G2OM912HWS9msNTyyQ65Rur7CYu8bNvLMrnLNKg5dhw
mDPebZ3RhDt7PfRZmQA68hFTiCsBLqSnd8hvzLZFPyCHyov2J2Ss1fBDChY6/LyvoGf6Ws1bJSsE
Et20leb09Q+qAvCZOtqFL/+cRnrxDjI2dyCdv3OHt5/Gtk9/mxc2jS45mxLhsT7IyTcG+zO6CgPM
3ICRXON6qpcVrERF0udNYKlwFK5CmTQRfcS0rTVISDufEPGLPXTx70wQeBHEER81cUDoxZGK1+rh
7UG3VtSyDtE42mI4v6jWrAXaWham7SM6GAXhSBDPgPwW06hVv4roMMVQcSLWaNi15PxLd9d6eH3h
259e1x4Ki1PyMPfepZ6Ktkf71Iy2hZ8zLRd3gmudf4e7TAkV2FCa/7O4XVfOHALjsM2jO1HhkDfc
CX4FoesYwHK5AsXdDWrRfQf7d6MTo1IzJURvalrjp/wDOP96UO9rOZFHBQp9+IrX1ultdBa84Dt0
cwNQs9woSGAX1rvtXWl/FqlT03gqoAySnTX9uzWQqqKEJlQ2AV7J++chudUOS04q5BDF77lS9vNL
D0YY0/kptKXe+4MoiS9oZ82UapLxlHMXF8NP5txmgOG6ju7GTBJD3zvurkwsS6xgTH62zPOlYUgP
Dua9TrfBFtJz0d3vsPB+V6QnRz63oMCuu63sAppJhpyZrhpNKQvX+x87fbE2Qj8mItiH1oLqnr+m
eGvr7+CNK7DR1X5eMmqjxe6KnfGxkGZ8PAcO/mgOYWiABYIslcaE//BdN1eqVjKFGMAHGMOJQYe6
xjafhHk0vnpkxEdYEGXQORbZHK4Zf3O8ScVdyuAJbljvCm1m1uPo0JFfLPaOHeeva7StD+6huK0l
wz+SfIWdUYO321xFbixQm/MXhKm8QT8n6nUF/2P9GdN5nqKofPFwjVKJGCvtxyRtYsSl1FGFQTkC
anUKW8M2eomMZ0fiiznJ6GY6q8AfERzk2zdV19c5hLlSFnG9VVuVTHiu+FQuaXaPzUhR2g5MpfVK
fZeEVtfwJd0n6dRtmzzPO3oMs+5I2Gs7Yve1RP8IRa1tf2CsKySl5cvFGf4OGhA8VnkjCTf4PbBL
gBCwh0ioScTxvEeuHPlWmI79rkBHyMkQWr/bJwGw62FvjckBPMkct6cj7PkNSRvVh0avRjr1Boco
lk8tjZPD5BSZwVag7n+WN24CJcUqd1qAMjhE+goMGwsR/5D9qNy5OfpeLQv24H5NCE3m6zoZmB+s
OuCCtlJJr3ZNgMNl9ONDS9BmHO9tfnu8f5hh8dHvCbTTP1A4rWwZT4+qUNV7YNkRfvsQ/vzess/B
312Zo9iE3yEYc+jptIbHjmX1tq/ZVQIzn6V0MXhgN6d98QwJCLL+HbgIUghP8qFeLzY8T62/gU02
sN57JGn9NiOC9MlmgNtzxwYSJLykKnEnUIO69dpty3tK+QXW8NRalTStc2gGCVVazbkGx2TjsDnk
mMDWJfpw+yq+QPvzIb16ty2kgz9dkYGaVuqo8MLhtCoWJIxsHpCNcSmayJJvMJcrCAjknYW9zlfr
5mSvOcvNSt7sznOq+FOju9UOHNjXmTocueqL/SX+XdcBUoD7sO7yYED9KkUa6mwcNJKtnz0F3u9O
0GtJ6wZatLx9LaqndoN/u4PjuG9CDn+bkCKdICEfBTf9I44nRuModpBBJrMLS6Zib0uprC8X3Ppz
vmfZSG1/ZvERDXEyVU9ZH6HEYUFZPSk7s8nGGDTqYd+Gmx3bAMPGs+aHHeoM/8i/cm6kqZbODX3s
PmGnkCYDdCa7XqPoeQYEbcvRODii2ifePaPSXU3FUFjhG6zWliG8qZzSYcWRpdykoqBdOBiSBNcS
fIXm0wOSplaL+R+GHgEtj89ADakV7DQ1dE6NhEcec7FwcCwPTEoI/SC1IiWqWH+canBzNOYNvDvy
Bl0r4DnsyEhxCIilKyZmRH97KptRZU709zAGAlfq/4LvjU3GUGsHJwKo3HOLIX1YdJHfKz420qTF
J5Fy6AXI7Ht9I0Tog7Qrf88WudhWg8kpN7pY2jW3I+LQ5DzphMzKVDzI88BTutGPwUE3VC6nF40h
1AEV08jqEMgXFdtF2OCv9h6Nc7q7hXq0T88TwIwAgoGOYVERYSzEKdHQVqFRpVjNT5LtcjmjliDm
yqKX+0Ijfn+SaTzH6DN2MAiUubSZEZnVIV8LdRYiy1fmSPD9MX9wZWlyvVY93CaZ4x3/2lkbIIIs
5kkij7ZjgzE2pftfo2IquedP5cNzctUkIgGvxy4he/Gx3D9CfreJJzhMsRQ9twoQjqKES4eHMAsP
nzA4EOOV6RKLPt9HAH/8N5Sb4Hebx9g6IlLHvMEyOp97GTbgQ/AYrXA7vu44GOiXkgaCxtdKZU2q
iNhqXmztSQUN9+Xh+qjcFTUSOU1kBRJPx+NK63iyoDWKZhLAP1vSFkLwfdnkN+BaiXKIws3mSkPC
BYNuuILhdqLmsT9L+bd+SnOoQ+aGcDmeZCTffTdHXss0JwlKVaDOLZ5aJ8Q/32a1DSBIUMR8G/aj
HRAV0b6QSpXBTJy4iXb3jVldnYFsAOulUWk+h+JIxLA10h7be25X1heCOoBITMq81DhqUU7r/vQu
DbCMxCshvi7Jo+Ua0Xb++fToa5xKCo5Du+fzlOUYduvla//oqaea49fxvLBvcRPIs8hKhzZ6JDSo
j0GcTLmsz7h5R6ijLI36P72D2SYKPybEFYUEAUVFscwTaYtyhQMTcVofbccxfCli2QkkwJoHKgPl
cgcd1FPp5Epl9iVoRNAdx5Kh5+6ct9ouXl9FWyqyiQ3JeleKJQ/ptOubHDSI54HZwqoMGXTjJbrc
a6P2rC5OPREhDZXDESXJ90xBEjGa4vsqQRM5IVcSUjesQyepNeCQEoiRGDr/1KeVaKI/fsQr2CIg
aAfao/ZYxHFoLjvCvxZJsyRY9m8slVODHzW1eOUyEAHCdBVatlrFWufgllpeHSqNCDusinA5Nmc0
yJT/GizS15GgzZtypfPsTX4C4mAiYXBjG4O1UVasKiE/umcPMJ/Kkol7Qjk5RmamwefnCTdhiwB0
KLy+d8DYRoYztU9B0PKqUpZPsk/3G0Tjksq/hMXIR9SYsl0Hf8B/Dy4pyZViNeijVJ57rEUoPk6k
W3OJklVz6leyZR/aImpRp16H/YAzeatxRAOnfLfjHXboFioY58QmijVQgtc1I3G/dW/x3T6L2zdg
KdcDyjrAgddqavjTAYT8vjxcPu0yJBi7OvWnM1rvQ5G32AReMBTO/VTtw2wG/2CKOFOI2dBR9GWG
aND2E8U8NKSxokqpk27idz9QAo4PPCVhZfwt5akosjdcw5fK7TFSuO3ZrIpUP/l4JUdxQjp3dLXx
vlaBY9yRfCqsWHz9KStaIzx6c68Si+eS0aoaoRKBPmeDxd/mF8xLNBwMr08RlHHwar7hlLaD/Vbq
8ht6RJ8Or0cX4D85lMZ+DP3SZTUZWYg3vZNfhUXAhCBfeI6/Az77g9+9mvLXldweIAol3nVh4Lmf
UgRuD0XibV2BFiQpA+bnXM1xBgMjK0zh51+X8T8/t20QsUDNJ6/ox2MVfQaET9PyEbZXSzUSLYvM
iVCT+d23DRlVWCBVPj9lzILIMcgNb0hAXi3jRgBwxG5eGKCGSkoBWqYoQIN4j/SAQRr/3LjDNM21
uT2sY1v6KKUlxyYrHJawf8dZFIAkzqEaEx7w8qW6ZHDNZNZg/uIEs7No+wZkWfcBMiCtGzxLlSzD
yEqcJvQkteoR2Npj0sC6eh26W6V/Hwye9QqL8OWWLvzWlgXHg6fvV+vs4anaFX/lYwU0jpGudc9H
S3E3ggPwrHfJZUE9u2MZM+D1TUD4LFeuXMQKeAPkag/AM4FTlSwRQSSjDhut8tRijkscgkCgRU4l
vEtMdouQtIBVYA/xmyum0qX+1Kv+pO5Cd7a0EkqK+POXoTVkHf1gb0UTKC+aq3D4qYX65PUZLZnf
UrIkUYpzhBFEEzC0P2lrQJILBRdr4fMzxOSd3Wl4AqmDD+VjzdCPWijAqsBuWBeeVno4lngGgF5c
aaubHebEbQWNN86IeQgl50odc5rIp5hv5ep8GNkt9qTj1580exAUY2/IJmhMj4fXe1pNglvMlUPL
2oyTqdUGOxO7wUS2xsbNDA1kzIa89XpnghJ2il8ub9iNwk2gjvzoAxj1wHruCEnr3YvxyXbY4VL7
EfxGAmpxyxS1KB958hoM2c2oXQ5hhT3YG5HxEkHIaMmzZCPZAmcU1X2DCPmdJBnTbZNPcBBvO/FU
jf5D69/9ETBxTOldnTVWwlq6HKmoat6TZHxlB0kWdq7gkjMGiswNQKgJWAn7haoakLIf3kTd3czY
p4HkQmirEoDleuF94IwTMEMAqanD0uFeUcr028JHnUsPrrs4ac102Ohqj9/wR3xRcI9C9T9m4f76
o4nbL/pRSuqHq90qal2L1CKEZdVsvp7GPiFVg2z48TytZsBPCo7DHqsAOrShIykPckHMtA5QB8lX
X54XNH1yS/Rh4EfYzd+QvwIuI8x8MM+mEawKVIO34gIjl+80ckCV+u15AFuLwLo5mbUR3SmvfB5S
1DCPM0J4OoK27i1BrEu3I0IDPFi1cKCgutYnVyI3/v6CToGYgvxWGu9bUllrHAWCVflwI3LfzxkP
AP0nDRf38D+PUDXmexalQ6rL80hjb6WSPFK1Srzu4/B3KTcjOmyhibj5hrP5CnupVkSuKOoMqYMS
X/IhwxG66DnAbT9W9gUXTxhm77C9ts9VvVo756c5np4ks+/PHJ5zxWDV664k8jggg53JyrKs3B1J
qS4xi5fmZ/5V90srXY/C6YUp9iiQGP9+J61b+cWFiaA7xP4xJCkPjpkBlFKO8EVbUb8in0kkCu9l
uJD98LPSffbLQQDyQq9Z6XHKU5RNpwYGK5zx0CeaBI0/4BFMmO/wh7rVojaYIgYLRYA7kKgMJ6V2
tcPTkLpEqImYG9qmhovaldIjYguaSrux2RSRUtKJO0poyreDJ98K2wXOPvQ2Y2F/576dUvyKI7AX
Nkr8npFc+rX6I5c7t3a4W+t+S2dv+RKyyQhMiFJBglST/J9dFlmG0Z0UCQcTMxJwXbDHTNZvJkgT
CjZPVcqgKu01EzT2bcQQHCDV7w9Srup/+KAgmVYJvXOoTKPnzGPaPPfsRvBwdqDz7r78s9oNvq/W
S8GiL9C6POu1SBDtNmacw7NBRsrTWVr0uIHCmwK5H9/60mYzIm0ez/8bh1X6i22teSPTmCOTIolF
6EZFnnPGBZ7a2vCL2K80/uuWuS3HI0yFKG116YE+6waNKey8XnHWxeAzBTEcRj5xaEu6m7J8b8Ed
JxlI1RYgKL9OVVlW2KMVypP5TTs1h5DFFq5UpErw5VRYx7i9yj3snOxkh0RrzFoO8KsAp9y3cIPj
ZmNvZFlfEBaw7XCw60XWdR9KxEsxhis6kfDw287hSwHQsu+ONJKvUfbR0lfu7x56jW/voGMKvXlk
AABxlC6M9+Mw4ujwmxtA1NuEgwXHJCEVK0kQT6ZXOsAJx7ZaFOx+K8RwiGC9xLgVmdCSYgVELeNJ
8TONwT1e8qZg76fziQuCb9ny6YDOep557GDL7sAHKEXSJPq3sFlvOBrTgCArZo9CbHEDXpJOfGKA
LZtsRPVq1sa5BPY/rKNxx7iDECsb1TXcvLgG2L5soNE789bF+3gDlR71XUWI3yNgdriNlyNbpwUy
ImWx+i6J3fuN42bpCYtDKepFvkHc+KDR4Ax27wyq4GaMDznR9Y9r8ZoIF3w+ovpjY4fsAv9Asjj9
movT5dEsfRHJdTAIKoOkNz3dJfhbn0PlzmjUACFEjBlq/DK6d41OXNlIi6V12L639qnSveH6atL7
4GXTcV5vM5/270sKoVLjF/ZT1mtl/8gSdnw+7+qtgCnRNfQJAPwDGijFmVcSpVUGv8dVQL8MJx92
7H+reXI5x8RYgjJiMd1sYzyNizkGdc8s8hgmJAovMt0/UAluxeCMPftSoBr4mBh/qUSd+9e/uvIF
eGf1YF/HGdVw0EuB/Ke0iZXKrQTblNWmyyfVee2U337QUwEV9wtsPlMTLC0+YJlZMAw85zaePnou
zLWjERJDqLxV7Zs7D964yFZuQcbAI/90fJ8mvIr2zHEf+j3/hWoTiUadfYMG0xppzbCNUK4KpWy2
dX6Ehm6Eioywx69g71C5mMAbEAzns/nNS2nfNxGQR+fIsEtFKWzVSzXHL4REMjf8bhgVN7OSGWu9
lHuDdbX0WCYMSxOsLTHdDASO/xpchiRvoIzn8csuTWbMUpIUcEXix2vYgswAqxiYDi7AprTUm7z5
7AxXpyTd6SAGlhyplGJ3z/Qlv7/GvIqKYb4zXS6FNTbJTRlreyOrBwwXOorzbPgdvj4Ns19UTcL8
6aBGmKx4hSoC5H1kg62BH/b9pnGGoxJYZi0mpMu0UnW94sOYHcOBWj/4zsAwsCO2bxFA6/V/TAFf
t8twm/5aX/A2uNwWylwjKw7mauQLRXJc2e4a4P8vGMcWvxT4weITQnoNbwMNmsswzQP1qdM7lEO7
FvcX3e57MlpyAnVRisBxh/IvPaGmQO0t/dISEaFVHiWs9670DK9miHYyoet2lWgqbk+VUMYJR9mq
nt7QnIGKbcTwSMio0F10uQkP5FTs5gR1vNFaLg2pRGaLvCi6MQhBrlFwzl8YS7lXuJXfHAin3aK2
sO5c0wXaGpHCwVBVnXfa9BRWIjTqMgsaVQ5BNvqeCmGhOtIcVPnbuA20Vm+e2QEI1bkJAoCdFj2T
eaDwvymHkrxzi63xQgi1sDuXwJw5LTWluX+TKPUWlBmLxqFeGhg3OwUc77zoUxkNHe8S7UWkuLXc
+c0SvjU28WUVWNM+tIAHpFXpaL+6J6rr3G3/S5sKQggmh5Omcxu/oz/J528Oayi3LeKlJin1AmyH
U4M3cerDBLsPpUYSmAKMco2M1C9PBcUK3ig8dKs+mSzcVKDguO27ChvNLIInxy0bcm14VirHwayy
5vy24QuI1w6Jaj4Uj+ck85CccSjfgde8PeGe5vF6fOGwbKzhFNOPLMkRRCxSeNiQSut+DBVGYayn
3AtQCq77d5m8vkSEEg4qunRULUEv0ExL+UyDcWODw9ahLaYtne18Q5qevoQWx+o9UM/5KTUJ560N
Z/kl5yKJZ7j2Z2NGuSeKgzMrVKk0TSsLOTqJpdMe86jicE7Rco8tZs4h7o8sBeChoUf0xd9dXWN2
MS3oMs0XUkp9uCKxrA6Lg57VHd5F4cak3qenPGh24Zm0/DYEE5uYHQy4wvKLegH5iaIhjh80KV7y
3Epb465NrcGJQqYKO1UOG6tH5Wm1aWlkTNOudgzBVR9FEeV70/dS4LW26UckNKtguW1O5/cerw4v
Nb2jAEFpTtYD/+BwyxoTswcIz8hO4QxMx81fJHfgtKkS9U73Z0AK/oWoamHk8j+E+PU+Ow24f5Ss
uDbClCOeDJc9yxrwtXj/taDj3cB/iLb8iEYeBLbjG90rysY/lUzm3CuN7x+YgpA353waA/MWUSbb
UNfPdfkKsvH3VujOOjxPJaBAe+4SDV5J/iuZql8TL++hF5yr4C4wMSuPj0hdYoEXUB2VF687RijC
q8/K/ubQz7XYW0uM2Y62L10SGHd9qFJihOhYmd8cd9mDDHuqGyIXfQhRUeujA62H+IHnR0Xowppg
vKh1UlUZSCO3/yTp7qupBB2UqlKvv81TBVczBeQrNv1BGyrEbslg5zGdK515jDkmOo6ydPn5MCcS
JJkqlOVde2Nu2sbOO/9eNmoBIeiLNMDBpM+aUXClbOFHrg+ANtzh6lH+eyXSsvlz4yD7N8Z4C6ys
fjn7elC3RrlYDnIU7Vh7EI7PEdJCSjv2PIZVLKpLUHInQ3ZDTI0Iq/P7QLkVfUWWHPzbfwz8F8za
6BeYKZ6+mueh2AqTgNmbU19YoHeoYxLxuRcrevuSYowuDz8FomptI06Igg00RaFeKZWvHK3pZO8N
xi+zso1saSTcHQs6eE9eIL6DYXY2bGyOOqJhKQPtHuQ+2saqQIymgPgkJBE8SMLoyCI/12ngUWcT
CtwsLOslvhe316eB6zhDlhetSiN2uo8CdKmT1w38Xbmbt5n+wK9jfeW5QA4hD1BTVDnGjq1MiPOO
6HVCDor8Cieo9LZO5h5mxcVqGN1XMwNGgQzkTbMRMP2fdfvs7qlwxxqkOEbiogAAa+Mf1QWsS/QX
hRYI1oiAtFBfhJ8uyDdzQYk1SCSEz40oPeRKQtyHJkJjTQvRxcT2ib2Lm3A8yJ9D7Td/18Ji76fk
6n13BPitdrNZN7x3rCdk/8h+HUvrxWlviyW9rLSONzHdzeCJBfSjfVRYhojeycmaon3dG8/j0txj
4GpLzpgkhvN00xHGgTALUKFgmY4RK1uVbroERGkS37Ox893qNIoZUMFmePpIkU3OQUFVsXMoFsEn
Ad5hZtli/LENfkoxKL50RUQSG5na63zWMOCHaIaVNtimvR/VUTAiyR/cADf+K25Y/ztfhZqcjer+
U5QS39M91VfW4SGv4Hfl/LYSmLycLW7HC7Ihf0K0S8+xXTABOK80QJDk2IFUXmP1/OTFWx7OeqTV
BsdYN1iuIDOaVgKxyUHMwD1vUDAOTchCdC4e540Chcvf2bbNYM2TxM0hbfUji4+3vRCHcf9V8jtb
+NWjKpGfa2DgZNNfHsHpzIH9PWDJ3R7Fqrw+mA7Mpv0vcnnnRSYGe5/EtBaUQIx1C8LHlZX9Ly11
y4Pv/g3YzaxPACmvMscFq/B8//kHe6t9AocuZ6/3EnFeNqNrUGtcjZxzWHXnwT8REZELG9+Ozruz
uJ3LDrCGriK9k76+zv9wQXn3uG8b2tlHnsg7AV9oIo1Hwzm4ilpTr+FiCNdu8YPUzuNVWeXWF8Dq
vcSm9BNkSPvI+7h4AINpVS+I/Tvm+mF+jxcA2SArz3uOt1UGv10FN+oW7Pf/ML2UDLvkbxOst98Q
2DeoLJUE0JQ769aunfVo/pPx1/LRmNDi9rmPs9VimatbE5KeN37EaB2xRwHUuJxdS/gRXHNPFW86
kLVjy4i/QbtDmGp5c8z/GQtgyqnu0nSNTsjl4uXyE77oyQK2RLWr7vxAeZYNoMjEO9vOSmZGOLdE
Xu9VT5J5VMMC1vusFKZF0Y8C1gNpHy7R4MVsL1PEo6rbNFCpsEr1zf4Uv6b0TbJrLCwwtkPjSnsB
XSuSTJrequ8lFtIIyMGw9DJUB4+xrx29HvYwg3yC3in/NsxZNBi9C2IPvouVhFTn191Pxf7K/tx1
BGHrK2onJV3M24RwL3PXm4abC8cOVvSqEfNtTqz93CK++3rdnv008LJRZHPGzJ+uFmL87dWH954y
XjDO6FpZUDsNdZCObfAyJJVpgpyJUJN8YC0YQNWMShiEUsdz6sulJXPOnsgfqFQBmgKFgbdtpDOI
hlx1jsu9J9B8SJFOggSgpVOsiEThFn8dqKMW7RoyjdNeulLEGUh27w5hN78nhYll/XGVup3+V3ei
yeEEQOrVSpxHT6Znra7CI0aCuyqPUUJzfvCTj5kE9MzL8eDqTEpvkYoJkEXoMEqnYPI3g3KVWXP/
bS26LAS7WotOZYAD05Vay2gDpFfT0Du97f2fvbfaF9hMO0ta3jAtioMWizu35fFRBlMMVWquANkB
vrpPR4ghYonWdt9BZpqUeZTgix+GJGTl0G+SLYFarewnqyubGf/6RNMw5EBTa1Nnc7byR4DIFoSe
melYULXrekqyZVnLxtegsoovxxNa7H1mg8Oez7EYWVdb03/K56CJa+L3ieEmwKz1wudnhUEMoilX
CLeRZWxDY5QTWzrhfc7hN4jmnOLq8cti3mZJG8rLY2ImyrokkEmUIEpRmg6eHW2jAqysy0uKRSHw
QyNeaONRLx6F9Tl5t+kWIXUUr/gh2vFmqeOKCbT7dFjEwfbPKh9CmdFU1vSMtb6SisNfJvR9EQ9q
bhZ4yjhnPCuilOqg4E5s8kRbsWm/wYMNOecM6wRTC0JKUXYMfamVQdHYnpYmltFeIUxg3RKaSmOu
3VYKkyNth0CY5wHWGd3u4oRgBGD2wwAwh/M6OwVWplXO2hbiF4z+LPoZ2LQhH94OG24EAaAC0vt8
TcCAPOSGMGYN3iAtfpcyBRbSAKToQiKmvBb6Yp0LUwT2+dXzTTMglmvnagHvznQjmS0utwv7xg8C
5WJmmI5k38dQjEtS5WVFD2mdH/iVRPwWwJtBsGDQb3bUtUgrTn0ISnfcs7rNa5a0/7SpIXHT+QdG
ftIj3prn1B+9weRKADPnhPHdNsDIYXrrbJ+Yt8ECE9s+s0fWQcQCtyUnbmhx3hf/13q6nJGGq8/Z
a9V9jvKbVvBod0sqDlZIKSegGeffUQq9wh+C3FQ1qlH8v6pSlW5Rixilcf1SR50Msdw00I/nxIiL
+fx2FWQR41qfC6dWVG93dcXMtYalhuIVH7PdlPXaeG6JSIU3KxVHF03IPBR7vstoOAFVFOxCa70y
QKEDL9oFxUGnWMZKzg3B3LIWbIX+at1pJ5eyUmi4fc2y6PouINAycfblSgckdqJr8dcIyHL40Qwk
j0DIxWcLFbtdbzJNy4Cr5VwvEAZ0CWbswRSBF4gHRizNEMjzFvU3TZV3Y7ckybkB4Sn306Lxv6XA
C7P0ukNhJwBJ8j99hUBiowKqHPnaWEJDRhYQWo2iUyifrZ+GShIO5FBiXWygERh3WH98evHUSq0L
MnNxYU6upZ1GNOg2+0EAqkegeMIUJKkzI6R0FkBBSkcd5Psw6KYl1zYr9989NgCqzLFPlTXDCPzy
DBq+6h6hamhitSOutIcyvPIO5+jeDNBBRmsbPyTxe5OJSLKhWmF8st90kT4jKy6BxilFc51RYYcI
fHIfqDaswzMjG1aKnP2mO0RBeEtD0pwxZ3y4pkDexO8HKzKEeq+4WV7Au4z3wcvqQvS0O7PSIF8A
pexiqYxtK6cvXOhppCg7Y8Z3T8xSn79zLt2bAfiCqIlxqwQ4CFjCdyE8ZI9pTntomHjxi1ru+gsZ
aRU11jsUqdH4+7g7A8vvegl/cUyTbtcceGqz7opPu3FFXuT0+yJOOPXkqL7bpBVm8CvwhToh0qma
kUelUrzdjzC7FrLdfrMEIXCP/8ZJnV9M6wiv8tnAvQnv/GpIb8e3KvbOz4aRivZ9L2mfJF8xAvgf
lhPNT4V0/LbRYacePZBoA+dcK0T7YE/v7K8EmDbjRRewwVZ+BMX0II0TkYQe8jKfLw8+zBZz2l9K
7h32UvlhCpxKD8BQJbKvoU0FrI921nyeat59KZsp8sjgh/mcJ4ele6E35TtgLdQ3BD4O4IPJSHYz
tMSnN0VDlIpUbYibwUF6F5eguJbyoatqQjviZfTL93ugg2L/lKfDd6hwrZWt5rNqrpSP1p0mIaKC
NCRLRgxSLh6rPqt/g8jJAl24T5jcss0MNO95fbWEKmBGXR0ebD/0s6+DRslVcThX19lRaYbCEwKT
w9SLZGDTFWgaiR1T101OizjCbj3RAlyjtNFbbwG4xtkyyc2+Wr6OFg4a7h8lzbxuW0aDMsbKwkyM
EIfRSt6aQBzbAyo5XOo38Z0GkeJzEZ/8gSJcvr05m+rWn5EDCkm0o6KBIRGkUGRm8DLSR8AYjpSu
LhaeeWHodagKQtKJW/KUuHOLJpN4X11r6FilCR+1uvTM9pGaDvqLg1XGEVxZjNMYYVHl77BaYrC2
58ZkspfQ3LANAQBIXUkFCkW9nRW2xxt1CEkHf8ok6UX4x08e+QaSYw+iqsQ3cR7cGjajsqj92Mt7
SNZMWfLIPyJesEc+7HQv/2abpJpT7HGaiJLByW5bkvfcExLrJfLL96ceYXrUImHgYd2Mi59bpAwE
j482PlUHZvDFSE/wAlPBMLFSRrIM7dpVCHDcWddSa6fgaQ5GLmFE7zGbwjxEvZjmZilUBtqza62I
EV6hpMCqYQH7fr2CPehJlExb9cXupKXg2cr6kTID21CJj2nzTwy511Y5dxklOioYfX2DFUlDIhhN
qhs4a9YA1IwsrEB8MUyp5w6sTgMsby9hJR4daRlS+vsU1yQ9COrYCDNBFn05vy4gm6hieqLfQ9b4
ty6yI0WVk9FdW20aonP+goyLB9SHmgZ2DCMx8azyDvCjiZxipDahLDhDURqJMu8wOhKHsTA1DI0/
QzQkxSwsuNhMR13g6ltqMnYoYJjuqkkh6uZoWgrswCSBjZYJKiSRmybv7UscS3SSggYC9fEE7y5C
RoaYOSjk/O80S6u46QP05gNza/7hSqDS5tQ7SfDrEHoz/vphXVYj7ZuNcau4c06wTjWWvf/mllWC
n94Qbjyq1cGQJZUsRaGCdpe/J+dEy9ePelTbdHsbm8EFZnliHqrGUsJ6fDBFoIN01gZl7uU4o1c4
4SFAzid5waYilKwNH27nObZRJ9Yp31rrYSecqASOfmU/DI6S1EKTi7YbPl3XfZ6P7Hbs4sfve5y6
/pT0WueQ64coDOYPcTgTm577gvA6AMymFR81s28CljZ9mWp+fahyoos4H5phrDGl90y33r3eJanT
61zMAvmD6MxoFBSoNZxE2RAJbpaTIB72/Zvso4IMWEts0yyQxDGDqsHbyCPDqoaQRikX8gjIrV0i
Dz29vt0XOwJgBUKCbTyt1172HJJvta5M0MWlAHRDbAzR+QSQJ+QnokxSse0ngVLMVJ9VaJI/E++f
Z9X3M9jofsgq5c9cRc6fUciN/SbFuPi1RTsIaAgS+T7STH978dzj58uflZTyn8VuGpy4+DHA1lVB
IzDD5pkEixtWwmzQZdm9RGNyt9sf833Ev5r9KHMxq/QH3PZF0zuGQxB4eLudm00gTs8M8hzdBi5A
CSmb1S+BZencmusTJi8lhIiw65x5Gx1/RF3w0Iz4Dl6hAtGBe7M4WB38FzEPeRe175W3IUVRsJAi
kqsG+mNYfLenac9A4QdGlRXmagvSot+FKxc3nk+IToVbkhUbmKeAtPcodtB77LE6NN6t8LT/x2vr
xOTQsI/DlE2SvZQaiJc0gmYokDYqDyS0d/lhchAuvwv9kCKO6BdGceOuLNBczSdAmun8biMf9KCn
3CGE42rg1dg6wnXAky2UHAil+pJbhEiDalsO4D26tkEJ9jmY7EuMmext5OOc+2SAVC0gvUjriFAm
Bb91JW7//o6Y6IIEtEWCgpSDAicUhPbSrjphOm0UOF7vER17dyfjAVVJ6t9ZkpQVG513MKQe52nX
ldj9odo5zeFfrYZwZqybFBBi1B+roH8N7rD3VMXK5eBkIWcvkqGd9Rvd8D/+eIpallQ5SSUG7VJc
ma317fH+/ecOhuXBXT/KZBpPQRgu8sOHAGx6XKTnXN2QjCk9hGUe69ot1yGLllZU50Jd8XkPOsFw
ttaEuWzGebAinVX15YYY8pdt5YrB9Ek7R+MCL3jgVkoVP0M7u+wNTEnsgxYy8+vtE0x2dAPIHA2b
8hb25a7RLUaa5y5U58Ib06YR/N24zSmN88sTHvWj7ZJ5PFdMHrXBZyBIquIV3BPVyATbFbZKGjSI
+ITySq6wIM1zH3ftk7tXQCtAlHkZcOFOmgjsgdz2gqqi335UDu+t/kmaAmsk5eZaDdGoD3MU/mgG
meJc0yGGVYXDZ2XgPvKOKR56P0ZZ8gUaCI5dJouLsRv2O9SCFHCOViIMICPk95hIbAiIImgeF+dJ
31dHG8/EAE3lekjHDTyavDQL3Td8RqD4HI/io3kAD2Sza7/9X0+35PVOy9OvLZd5LhjgLmP3bmuF
xlAFY6a71qIe8TLvHFLUI81fNy55DTqq08d1HMSlY7J5owu9TNJV5woNCCk3NZDr0bMOVnYMWCl6
GqGKdmzD/vuQAntjvDOtjH5b9kjBfT11lyMAkXDXJ9yZZBGeUAaWrbkUlt/9RtjQietzq1miQc/8
HnEVqQO9ZD+biaFlnWwWz56/y1rAmTWzsg/E4TM8TsmZf4GKur8cPnbCIZ22cIox1AsYMVRD+rey
N3N5/oGi5uZhCN7GAJ1kR5q/wGnGh6I8T155hCZkYMcLTbGVlzLQsYh4TyR8srm/oueANOQYaLlD
219V+6V/8IKgh7uqZAf3/WpoBbyANPS0XvYiQyl31Re78x0utkyDyUr8EqyvY+51h+ry9JwwEWbj
LtECMqOm9DAe5//jgUp3CSlXEE9dixFiRZ0AsjFjNH9tH/B5n0C+v1TyXiuU0xBAcUVX8j6LPN5V
P08Pf3xQz5FsRoQlNOSm1DkBvyR9uyJV8WbwCwZQ/17B2Hy2XhiDNfTtTMUpXsWHYb5xxCKNyYA0
YyxVYJ+AkoI0/6tg9sEF+o+VYjzH1vFZRkKsRLnVjIUO7AQsP1n5Hf7guOWhSH0Q/jWFUsLejF1g
fFk9xSCoxd03UGqIktRn1KVnqWF9Jy2rYNY+TZrP3UZCHq4IGDdSoCuqY9cMsPrYXtt6XCvErgli
eC1CLkN2OxYKN0r/Y0fvgmdHt9WY953fczk9cGVahSPuvVYR0xzdDevJkMZURDRXVB05IYWl6TBA
HXCeNfX/7N23utqL2qH3gvmEDS44yBOfXFJMDeN42QWTHG7jy0RgoUXsUKvaOaUSAXvaI5200yoD
WvQFKpUPgwxQdUHoaieUSn4SK/1POT8Yy0wOI2nxjjAteIgwWD4P4IqWDMQNLG1c9XZF14LHgsqV
u8kePsKrDdmWujg8BoMlL/dgQ3TL/hrDO1PyUSU/B5n6bpu8JYjMdNfvNuBdZ206brpOdF4wY3/s
j8s1aS/qy+iZxWJH3GUl7q2QKhLUvkuUhW4sp0he3lmgbLXx411dgFRHYoxGN3Bei65tqDLiI8r8
XJVcT/iefNC1EmlanTxdVFtTsaFBU4Cxz40e+AfpuH1OdD5HAyiNEeF5W/2NcmHDq924DxiABEx9
nPdDFrCY3NP8jrNa163u0PSqWLrxSGo8alFYf5ciEsNwQD0bA6wPVEFmVdpwsb/QFYoR1EmOCb6p
liLfXxptRvlkDRSixLeCa+qEMCgUUr3995ObaSxHBBl6Wtx5EdMe3IHrcKo0KWdJcKdnT1cjIONM
U+BRFPvRtK8WYrSoRTryC62HaR0i2Jy0dEVzzdAw0wRRAFIczFo1dZI3ARKvpz6N6WcMQfYarDHU
+6+Gaj+2NahsZSuBntGEy1ky9PPTIAa2Dh/PIy2LOn7dlyJCeoZc3Dd2N6bM0dJrzQU+taZmeFZC
6YdNKTqaeiwB3mHp63cxSu9rUmYcodUfclx4VkcGduQx7aSEhozzO65YF2ONbIWzb7O3MbVtfhIE
wZSCScFHGKbFjpL8vGWP+6n2LIibfsy9UzU6+x98nxMoksyX8K0fiPSAjf2236HYosoG94Y4xHxn
k90jGmraqKv9DhRGuiZyPvkrYGlJunPJQJW/XlWMc+mVtcvA5HOcB0zTNe7Q4AReVH1a6jLQReH4
H70jZBsekV3xSK2ttOck+FurW9d1+uj5LCLuaI27WPSoRBLpj1NtvdUm+WkvdpM+SyDVanWJ1uwb
N9lkEo75spCNADommKg+9goW/U5H1dwedEPg7zSH0Lr2E7xPo6OjtOAElIbPbAHCQf2QWtV45/yA
z6FNAqwBJSUB1hqyr7iIBqB0DyELU76sAYIhILF5vnKzFvxGIzCa3+Yc0EbgxXyQrE8/46Yi9Ou4
oEi9te2nnvevOrGdegzTwm5HMrlzjyc9LcGm6buPE8X19zz1olq+VFCjjyt97KS1XeEoPVG21cjw
O7v1vF3DJKp0I1PUOG39Mj/ZgOkrHrjm6hYZjSvR6aorYDSh+eNwK9CIR3EueOUyHJsxdYFaC1oo
p3h+apghEesUEiCVs2J9AaUM7TZQELQYKaAtDAF4aDsVp1/sCqLRDebUanNx45A4wur+zthFxC7t
xjD3qOM2QN59VZTNejH00ixv9Yi5kP3YF0HhusIjlxgRqmf83Am58CCK4Dl/QUQdWJFnQjYObFpk
HudfhNWFI9aZvp3XGo+fR6uC5zE/LmbHpoI210uaQA/asSIG8O2Y9GKBK3ccYpkxUiLlP52TkKwN
J7ml/Uxd+w3QNW8pnM+V3h1MR9VJIbfjXBY6zTuzw6CXNdMeC7CbHaQNAPCZxvGHXxaaTyrRJWyZ
UHTKh4VIOiB4NeZb0WA6kuAgg3MmQZvn9nDq4tlKP7t5Zac/hZ8rnFVepqtmJqWaAvItsw/R2SWu
WG9k4LeDN2OItxBVhgv76dxoh89EhaiSj7EBP94d+TSLB1FeXGNCs6b0e2OSxTW2M/kLNauc7dmN
ciYBfX2kHUry2Gibo9BO2a7bLDyxvJgxCYbrRgILShWIsk3iRhFIOOOW31RAGrtmUoPLkmu/8Kms
MjJMZhDxPzaoCkHEmED4nExzuaTk68Uof473QUsTd/F6WNJ/GTI1hsw9mRXRiBwSsSu42YxggUdM
SYrA3ZEwcFugQuPZkCmbmHXdShBmAyaZ2L0Onqqdv9mt9PK4lu/NWW7Akuwq6YZGRxyrwH2k872I
vVoBgm3muM1gNU7RR266iQ7JHNcGh+j6ScSBGolSkj/P3MhuJpXV/knO7XVNlm0vpcxrzxgOZcdU
hjbxjIgy/Ky7Btqkxoh2avpOpALUzBx4YAnwHKeWLOMvhUcdKkoj8nasUX7sotGt+8qSZKp4WlwJ
MmJlEoZjMBdHpZW4Ool6hsiblNStA2vaR2lIWP/+EdzMvpecNnUgwda7oxLP1SA1WUqoKYQTw1Jk
2tjSjazLFOdwLNl6dMz61RH6+uXzT1qw4ruwgAZSOVM7PHXf/fSopGTYTPP8MMVeSH9A/1ISHDHX
9TK9/Vxq6Ncj+4+Mbam2//ZJzjCeA6U1CqhWsqVWV3dh2xbhWT8M4Ucn5F6pNeh4ihF3BNl11W5z
PzX4JrdXHqvvCB5Z5pSMLbkAiHZwaCZwAZHEWQgSly0T2uM02SAmtext01hzh1/jkJDjiKUrigix
SHttbfxD4lvTR9XFt2cE7CXkSv6914YJIH4UYS9S1ejCeZtRmWjkCt/OczFefExm3Mbkfz7dOOA0
SvPqjRKGY5Bul95tnyDF6WdMdWUxFB6sQOc05y4GWLVn/GsAS5qYKmnLYvS7gx84QyRaz6a9CzdS
THUwAAG2PU8UMBvvZMGsAltYVct/Vb45xQL3QVVy0gxf3BdKnJwJqpCBILr+taazeRfQF4FXEHM4
XT1CxuIHNNJeKVHHI+agUL6LIjPirLYdn0vc6b6ejBCU0zzWrBGvyiC2v7IKsTLDleyjY0SLjqGd
OlHUU7OBOiMv1wu0/XzLk7T8NP7GyIf8xOJqK6SGxR07lerTOKnV8173CReyA+/NbttKEXElEFcU
bakyZ/JP+rydfHdbpMDByoAEjTetJUbhc85iXg4W2ZBh6UlchiiyPZwDa4n+OJ/9eGKZSHSi7I/2
xLxUIHq/TutXNqicl5OINh3pzOe+sB5icasSI/+CakRmz4t0Drhr8fSWj3LRnDmw5u/P9AOIvUKf
0WPZwsXbJEJAR3P7RomKN6htXmWbaNIOJK8hw5LMsUHyErhF3VNOPHhVAc/W3tQQegwWNyy5z9A2
hrQl3HzYnUKsRadfGYXAkiD7qpzpp5XB1GvU1VS2YaP87i2QWWBbUkn5FzMNXyPIpJC7OvK3pegy
AoYlAO0Aei+4T9VgWwrBHgu9XGSHJEvOGp+1CjlmHOredLDTTJm4yzMy0ysmGAh/DLEQKhVptnHB
zWetHp5J3HPROrC4QjEJdqYc/T4aC/eI9SNpxHSeyIWuDlEzFztmNki1pk2Z9GFutKdyMMqmQTk4
Uy0hKJwt9AfQzUXD2JuJdWnLgG5qFAmeXw5vCtkWRoRjndzXqq8MWjZxqfqF5B1vVqjLyFF1TCMT
mPG+HKdJFoskF89xXir3Sj+HIE7CpZb1bEYaugQJ+jDKucshi1BX6t7yt8aY1XW6nU3y5lxDxaQM
W/hmIQXnsPY1GaNQCgL8lJMEPhSQMqONn3jt0nfqdr1pYsYbgKJUaheR3axxmVCC/VLCFf5K10bz
iHYRb7T7pYU+Im5uF916OdtIpH0EC6Bjps4v8kQdE0TMuv4b4x4u3BGM6eBnOf/E+6rLZ3bLLqM0
7odqp3ZDfwkPCHyhHQNJq55uQkoTd8zhpS+CB60SEiZ18+uE+8/6ZlPd72hN8SWS5WFuO5EeXuL1
/Kcs9TRxwrp187MeFa1WlcxGdmnF/9O9Mm+9S6/m5Cbu5JuffpsveXc7QAxrFKEocVyJG5h0uqbo
Z2cdhvmCz0VvUH6OsxNss7XRNUobYWue+cqwf46xmDRgyPS5e6V9HBEY4/FcYhlyQWkZy+2bC2jO
7yDuhKvJsLWf5flWpkuinGwVmgb3qV6VviSKdwInahjasaTXQul8BzCqs4yX1zZtu0azLfM4gts2
oO+YjyaSloJ3bzyZ8NH+RGpLeliE9OgCmIgqw0/nRbgNrl9fkSZaoPPsbVL4iJEyfABoszoS8auG
TNqkBlZpI5xENJRYsdGM5eOh/GJROydc/LxKv1fn3TeIjJcZ1F8V4wudcca1TRPsEJysKO3WqZxw
RGvuC/NxLGCLxkNHFyl0FDkd+p32f8JaWDSo9Gq7U7xr9v+nSq1wptdGI7lJZWMaL6c8KRH/57+0
trQ6FJP991QdaOCdCuFT64f7jiQf6M+ho+hnpE1E+cYvmfTmd7bB0tK7STauRvJYiyyn6P3whjah
B00CRLFNI6HJywJ1I3h2sDg1o+imgIgFLPnLQRbvhKtDQMREA4Qgwh0cdBgmPTUFx6BCotIzYnSL
CxC326LgSQa2HIgFD0yb3QcXafsPDFDK+xD3p3kXofYfv6NWe1K1SmVlV65UtGMF2vDDXYGfQ6zl
k3ee7JZA3/4d42Yr0HVWLpwSMMxMKUlwRVfJGUHz1Lrn4kUkIzuc3p80k06Nz0Q/R3yWw7bYMcfB
i+WTu3PghlQ6llIoZAoW+CtsrpPdNRFgYodbzgpaSJK4U4YM2lmUwHH/yeKnoWpj9LbScXLrtdQa
30kyFYOlZSQGFqNuUEPgaEVdo0rWkDz2St+378DI8pfTlPF2isGJjMieSs787zRW1hD7jXN+BVhD
PAGJPVAW5dfuHyU2FwyVRL7xlN5esK4WC5stsF+7yX8D+AVlNWwhwguuv2A83U2zXFgzPMaR0Onq
l6uL+s58PTBdSZEUvwhgCjJk+uu+PrK5yrEJv1EHfpqkx1SUjoYrU1tXM1ggAC17WV1sXptbQD9q
QzqLE9rWygVpGX45/jNioMonVfwHgW0ysP5WQsfo6uaW84CtKh+mJZK3t8/4b9lNJC2y5Zpyb7IA
6PtSb0WdVKJzeIRv3cnhIqt5Dgy5J+fvnz38GZXE+fy10U+3r5vwj8zFf1QS4itIKv9ghwzOAE3Y
Rr0XpiPLK5f6ZeNOU3NTeepuEARzxQadnYcSbiELho8ndfR0Wve1Pwv0akQHYJ9OpArJDhH9gjMc
2Wk86FV9WoI3A5JRktebxfUQGrwxX0fUCa/yKjnQLHD0CsI0+2m7rH3JTEKDKwjjzTGRuNuu7B9N
ozq+u7pydl/q+gxKlYqJ/Ug3OrtLdkkfcbEaLdoiOTTnjCplIdhnL/ioLvB4cvx+1fnqnDJJ2ZQL
AYe8XcQkjbe5CYr2jbyJOu3q8IwrjAf1dV6eHjekaA3HvjHUHVtlxjpVGfSQPwUbnIzAdY1XnC0s
OsXLPDLk4kaUFqkUdPO3xmyV3FCFV6drLSnwUuymHVwVYHhaJznUnJas4zTjHtpUZEMuxU/Jb+Gl
Mbj2wspslCm4RGmSwdNERHnAfbxEES/6nSQ8SqMFk/4l4s34xiB3EV7BULl80DMVNtrTGpZTkpfY
rirUt8HJCowGyVvXTHNVivpQAQyLbGOc9at63Q3gMwnTqkWWJXn1j+YCPwfyp8YPkR4XZK7TWMRG
VX5umLJdnXp8WjUnoF81LoavI2LnW28q+7dFKFVvHoudQlp07wkJ1KZmdgGPu8oGbm/F5EkUAHl6
1dHURuOSp7QtBPZxc5Uf5fnD67/oizQxbzjeiP1czF6Po0/GZP+izm1Cc4QdjyVueBoczrR7MJOf
dGUhYDARJqVfz5sa53ALEIsxYYP6UWRuK7m8btKQe+NwMwqnY/jxLvPQcXwqcWts+IJ0qhdQfuMl
PElFYwROh4/8mdTWdEIAYLKUe4oKDyKdXGww2OY2MiMAH7bzhmEdnnKbmIaQcXT1NgR4GGmJxCEv
MLLNK3qTokJewi3ekX47k0968uCqoQhQetJ2gnBGzBhdbEOYArWNbnyytfWINAErUNUVMUkK0gIz
jqHJo+r0CQAV3dIC1eUjlUOmZuO8Q5elnlHhK+bOlc+SkUmt7+p3K5I+ZXC23OwQP2aV2frfQ2v3
N41KCmW6VP5NwGSMRecpJpCPCQmWGLTAQMcNChbukeB2M2MN1yEAZejKpj5vqXoEdZK/oAc6DdI4
vsXog1PKWniqjZQOXJH3xOqP7qdW4D/mYDfAS4x0RynywQWl4iyUIe+OM364Za/sWRVLYYQwb52w
vIv3zKDsGl5UVGAWriKFVm3ExQdrIjHu5AdfXdP5alvIjD2guSe+wE6mvQu+TCpDop1mmE9S4sN6
cDOh22k+wvL7poI/6NIOzrtNlqrMRyEJgjUPxIbHpVTBbWMp1XhPRcz1knI6nUFLljYy448pWMtg
lkhebb2xNYQqnx2syhTncaiVxF+00DA9CnhNwr+zesNF+4whvxnLvGzktYnaRwWQ9KALm/RG1Wfc
ifjTvuO88MogTa/3m0GjiSOeR523qNUZP0ZsMoLDEi2MEY8cW1BW8qCMtORi3bouLBZxiyHBJJ9f
62fqx777B0FNBS7dh+znFdVoYQyaTcFm9NQ5zyQ7Rb8hsX3TzoOb6sevCu3QcbF1f6myhh16Xj7j
Oj+enXoNavJhUvS9c1soS0m0aWmbcBltmMUy/LrC71SDuVpoHWoIRMLLkNnTj7GdMgRdaf6q187t
5sUoGueTIzrzu6nyZU7s/8dFZlqH0nk1bFRMiJs0QrgqujOj/aTYbx5EuFk2h/WOSebfiSj6MC/m
72aXrnoGgYXJPSnXTFAct99YDUQc4b3hItEtQDSAJ5Xn+E9JB2QHQ7maaYm3hsimSwXKokmqp7nW
E45T1AvXnGV6e1MABcStyKbhdKPYcqg6fwshYdieQSt+lDMayz2rG2uc/ZU1gT4DDW+aWxIlnUmL
yCkoMlXLv1JYdC7t9sW1DvqMZ7RO3bGlpuqzDPFFb/Xe+Pf4LtMZIPUXnh2F4EWYmy06ajWLFBbI
wmnAOQjjJqAZwKEM4An6dow42RF44iC7zmb/8RaduzTL5wqo/9c3Ey2x10+91UUSe44UcEboUjoC
NEulIWx+zCxBd1ThDQB/5SwGbtiVqhCd5fZ9X8v7CFQ80swaE4Cc4PXngGW+VVvP0qsSXKkV510K
ofmycsazwh1Q8iXtzrH0fG29mw6n6WYRW/a0AWaZk5T9xY1twxVcY8qmJwY+QaFowQe4sXVP9DvR
fkEg45zDBTLH4FkB/MM5KXqIdYsMYYxf0KSOU+poe29BTj+JMb7ghvF3R0Nt8mwLAAJrsbJ7lz7v
D80tvl1iTYJ3Nh4u7zCfqhT+thxzEyK268G2F+B0D1R4KksF944AGbWdAFdVApjCC3JinN9j5xRa
ljTIgeR4p0nMc0qsFtqTD786W9/KrE/ffQO/Z1G8UI2C8/0dhfTd+x9+2pH5QmBY3Vctcmfe6e4m
LLXv+Oam4NOmYKYZJ1NhBLy7u6ldfzoU6ytvG99GPbNqbET0yFrDn1tFClFVQdlM1GFeTWUrGCyt
KpWCsyl392qZtilBtOTae7aNfBfLtsAxUVZFMyqr0qt6dmtcobPeFa2cQy/8mOTiqhlWJkhca/Mo
htN+m4fBJGyiz1Hs/iYOT/PqaWZ/0yqnkKIOZE0ms/r6tTDGlOH+LCroGrd9kK5N1Z/PrHnABW3g
aMZd0rHUDqsWSefzGc9ISAidjw26GF7592OPHR5jJpzJz0Z9JCZOV/15gw0jpEn4j9cHRMGRw+KZ
USkJyh1qe997HAoLl+qGxPyjrbA3YbOeYtIe5JVgRgV8+W5M7/FWcoXG1tcekvk8BVdo/lwsxUTY
gu9YHEn7UslzOlt+gjBQr4kUQq1IGetlLA6/5whBkpbM7pXEbcReMz09JMSB6GAv+N3NQXBIvhiD
+xBRq1VIDdrkoHQKPgCBR0VCjoBb+eiXAnP+EBjROCWCZtYOELPytrXEX1Z/j/0ihqeXKu2HLGEn
Y/tf8206ZfRNd+x8ZbsV6pDfFxf0TnmxStkizoW/SL6I5/SPilpfWrJJchzzlF1u0rQFXYNX+vrh
DQXprtBa8jT3EFSxUtpxTCrF3Wn6h9ErTPzzdBvVhnaR0KOe1H1RgcpXgialQUp+u6H/XHVGECP1
cNxm3EMkDjqyuzzJ/xAWhkvAUsz5R4jGlI+UwEUgUWsS1gU+nwY5Ig7qaDK0YqLOXCq+Em/+79Vv
mZjYdi0LWlJwHzSVLT2LWiBQTciGPUTMhx1/NvW+qG0YSxVWzRssrOh47qpALwWiDB9Ug5SDWpAN
MKcZUOCNUTz1FVq6U42ShekhyCQg+YhtGKQ3GjP9lVFSZdlMeNNRrjzg10lf8SEuy4lBluYokK5r
whBDof+U3kqRh5x4jD10yFG8mehoR4Z2YMgeQUXKGKZG02muLmvBSABk7DxzO+IFwE+zfu9sfLV/
ueBvuR4HPKpkoRVZIsCAWxafFJKU829adezcz4eX6nysSeTPEEcvYOU5WyPknlTd4VM9yA5frLIw
+lIFjsa8a5qiIoVqZzjd8h83ycT0Nj/UgiE5EJ+QWk65rHRiLWALB9x3slDpc2THLkI9nd3vyhWz
V6xefoFGmwIH6UxxwLHVkna5Ee1qvwn/SGuEZt6iu6PhKvvN6WKBhvdUp492om8MlsUxJH86nqtg
xFcGQc7MrdxOvtkUUX5hXSiA07ZkkuuEJwQbl1EBimnvPpJ0nw31iYVBRJHNobNLl94AByvAeFge
bjNU6MbaNFkM7V6Wrs3xQitOyDwU7nu2BxHaVr+XftlPQ4SeVI4VDfpWY9Q8u5K8RmdaLbRcja8B
w2WSRc1yQL5PtS/Q05YMAFFQID76XY7Qy5upg3OhclFc6rl9+dcOHyiafc5vrmQm/Y5u746NadtF
R6s9z+XVCzJo3N4vMj4BiNaCbzheBVlQ3WqigFeR/4gZbnDLfniAvGF3ho1WMZOCcCKN9Y1Qc+fP
MxNZWn++eSKh4K18i49es5TXmPkZGg8QVX+4ON353eV5d0M6nipYlhIGtizAV0SnSXuhU30mwoB2
/JdDVhDWl25AYveu+iaij3wYJCshyDjLbIVX64LYjsNASSnuZGx/vxgOVH2SJ0UR4Mxk7H8rtdnA
uy6aAr24jo8XLGQNW6QeImn7Lip+lOOZRkdNTFSwKfelr5ags0bHJcqTOkQDi7Mw/MvBi61ed9uK
MFVLwoYvj6sRs6iCPFI7ub+sH2vRgsdWbpCVJSwPeDTTj7NVhxmtY06muohxbjEgLwz1v0ZjlsHk
gG561wUENp9KkZ+/ZcnoWPCpxFYKrcGnlbdmyn6D1nH9ybvupMOFScZsKmYc5Si5Z8uzAqYL5H0P
RU3mauYlns/DMnKqTw5LKvAjcMgmfFynQCY4qbDbBTYjHMXXElnsM0HFzkVp8YeV9uWSBk550Vrb
PFaTYHBhQ0VuLOtmspJCseLuJaP+7wOpp4D5PxgEVlA8j6mKKjkHe6fgxauA5+0RZhi+ZFJR4KW8
bPVoCPO9z0Cs+d0AA6SZY0kK/SxUazFBZ7q3S8wlRiRu3M73TvmDSsZEY2p5Edc9UFC8kcYKrP7R
Yn4cBzRAV/RhhxJ5RxD21jOPaVlY1RYJ4b+0G3E+zynR5a+4u5APCz3uohZNYYncbMd4lYm42DqN
C7s1RzVFX2HNe+4U4eJPYF+IkYwJ3q36NMJsPiA5Lc06vWTWC84bM3o1OWcjosV8X+XRm25nxPsx
FJZuf/Cd049Gmhw2wZcc3MzTvItmm/iiaXoH3EyOLB5bXeDL9AxVuNeLYsiYhsBOfdD15tgfnzhc
ScpFUMwlBvAxLMo4fmSMJQ4bsAq+QEpptVABX1W80uPvmKNVMYuV87KgUlpAdxV4F/HHGqFCylqx
ULN7FL+AujAG6g6ZR6bN9IVzccH/Pv/QyP/nl/2izNCVmHhd+g5VeMOFfxLkJSJja+PiG2zCrqZn
Ds4AduGfjdOmuO0gFy23fxMgdLv9SQFO3IVk4SAJw3gP2koJL+gkGGHMnrl3xcZxvILRPVj2Df58
d1cE+i2nA3T05Enh3PjXp3Fc0zmLGeuAocYj+kIwILt+6T5PK2UijTHTyNmuia2bMN8JdfCPNb1l
oda5mLEaRa7gnIBp0lGVYQVINxptU7ePrt0YP148JL01dXoCo0aTGW0FFoVmlQJq7mT0C1dd/j2B
zlmuY+3L0xpt03tEQIYIm1/elyG7SdBrylWBq+MQNlSU7NGAx7KBWdtzS2en1RrlITQt6Kuj+3Kt
Zxu97ZGqbzdaECNCccrcz4Yakf3Bq9suXlhLC1rqCtKbBy6d95e9gR2et3eKO3dlOohzMPqS4wRY
ckXKAlk2v5yP6qLezd/JiDTKS4BBhyj8zZSZcgSmDQHAMG9lmwTr/aleR7CnRQp7u/E9k+vLA7lT
lVI1uVn8XYA1RMO2RAbBIoRIN4PeBgBMb78ICXzkpz9sFxxuoXmFb4RcbCfQvCWyCyA8Modraehv
rw8DhYp9gxTMuoODS6gBOhYKI7BE8Ybt68pEmOK3m1py5XUEAViEMipP+0KvtB9cvwDFlUgHHXa2
lPxx/Ix0yuHAO+PL1zZkpfAa3gYUrRg8qhevJdqR+hKVHp+fHS3m1WlTaNadIvkOpOWgt0jY/W9H
z3CSanVyHEXyS7YPPfAMm1rrdjaFbXCq8X0YRuLixjm3R/E9OFwmOHp6yBgko7YI2x0kZCQSXbPG
YbOvGKQE/kcu4ICvPTpeHZlaExsOaJZlsnSiPHoEOEfMjDOZ+7Uy86Z/GL3mE8zlORWhGbmfrK5Q
pktJ/de51M4v7ZamAYzTbTTcCijTXelCOYJxrbg131pCFuZCMFPRM1bvarpFWIjK9sbya3kS1Id6
8CCM/ybSKZW9u7Oq/kRNAS9z9HGLaixmfvkSvMrbSubv9Bz81MwEoftw4jdQ6R0mImsznNkJZfsJ
S16IDyq0cTzCu4wbn2MWrlWHc4mbWBIfKKERHYzYVZVF8L2XmhWXb07saocTkNbBwsC5rMOtj+YW
drrZaYJ2ty3+J6AVtsnU3dnq8nEzZvX2T3Vll3lKZAae/X4tHNZck61Abb9aMoaelRfFE3olNVDz
axzQjRl2VvQz/xXDQgL7S0XYkKDUPtc9sCoQYwb73oQlnkyDPHwztt7TIy7MhtVDfwZHf3EWnNJw
J64QBAhEf6tUYPThVDxWZ+Z9kLpX24vh7gTv6V7i+gpUBq9vJdYOXJWL6LKypReDarYGkZJyc+up
o7lzPI/0VK5XZWtk5g1U5LRVfsIGJtkBOPqeQSlh22Yy1omz6V9l7Qhq1TiYTFe4FOc/Dlc/ZGzz
ez53upSCwcK/NBrZdYU9Q/5s7QEs+uOGkHfqd857Y6nyr2XwJpc8UsJUjipn/uS2m6uEEyiDm5n2
2iuNYEiKH34+Glxz3bBM8X5H+4cTQ4ENWSdZ34XWIYjal8RDdGrSV4aQH4fkvVVwMcPnrGRvxLgy
JLdTZo3ybxiVzbyUBPFpLZ2BGOmAwi4KLatDjxha7ogU/FepEgyVlqKgR+X75yiGdOasuW3arwTE
4RWfoJ8CB0eojxtgh2ueM/UP5NZ+qZuhZTOImpbHnntzLREX+PuJp0hRx1bccDFa673w57GaqawJ
7uwCiT0juvnPxbjxk/77+iBUPrLzz9hl+i35GfQUihzBXkIlQDRP4yigP46HQh/7TS6ayRUBxcaY
pA+xDuNnQ8eIzZily1+9f1r/6JPujeAPJe9YPP49kHTBdvq1tUfxR+vkclf7LGR92YfiV37W4mZu
Bemte2Xqo5fAq0oolXhRQxsPtsWBPN6uNs6d1U9gDpmp/3B41XHKGjasSTPr6tzNVLvIZQ9OEcwC
fW4Yp1rXKN8ifjzBT/n/l9KnmrNAAP8ofoEakYvJdeqnOXPzSjrUjV+z0Zy/hPZXOtYC4k4rqFKL
2A1vkF19wmM1GBMZnLqVB7QeaAmP30TtKLlQbfKlaHfC+GHAIAGmeFxp5p94bKdOsplLAhaMtYJn
iak4Q+UhoGXikbNHykTHPhLPTluLLk/rW0O3RX72ww4CwkkwyPm7Hw0NUtlyXjLpOcdsOOwHVqAL
dFcFEBnf7w2965hBWj5ub7UpIyAAt625eJ5vs/4lWp9Cd7/wo5OtvIaYGk/T9Ad7na53w6gEOi5A
0sFgBNA4SR78T8m0em3Y+L1FwW9WrjQ9qAzHkzZCWEdb+ayIv3YY6jZUxotjjoq4nglyrhigVD0B
YtGLkUh/LPxhn6BuJTpKvLnFRoBRlX7sv+gWGw4FDpNfvcOUAzUeLvL75jIbcR5bxggDvtUqDRIl
4tLtk75MlLt1Sn9qqhaZ8rYlgtSfS61YP9OrseQx1+7sGlDBG0Yd5p/RsV0vOCsuTOwuOFrEtClQ
o0EFREiEftFzadijXNC61RfebgR8alvTtwfgEkeWxhIVAh49TztDg2myKt+srtJILILeY3tRbjl8
UNOus6lF+MCBJAon4fnzJwCvNUT3XsZNI5tlMLncMZPc+HPwyty5K+k6kaEMbQ6+VdbOHYeKmHZ3
+DzvhQXeFzf9F5/uKJwgBx86vBhtI7dXDvG61BAFoNfcfxmUwZPW3DZtd770GFD+9R27wkZd0fWT
xj8uMZrdc7D/uThLbwJ0ZEGjPCmE73ZUQal5rW7wQy8lWgjUnB8FlwhkemSlGqoPi+NLb0F04PgL
3IaWqn+I5iSyzYRNiLSqv54WgGFNl3cYUUFETRjIMVMGI255KFMJqsx12ns8vFeZrnWC1Obj+n7f
8Td/Sc3dvxV3nLOib1jWreIk6iPlkJiKwBNsuKAwTsp/+WjLXrcRc6kV+3x6plKRyDtw1YoYq+E/
b5GLOvj+tNCboTOdw2QfbSrZM9V8NC3+SdhloTpdMM8CXQRtivWMYb0c5fovepYqxMsyEGT/veBy
PvcaFO0VJImUSGw3sjl4eVLsW5g6J1S94M0hgOn+jFj6t3ENO+hMvWxdOBZaz30Jt6h61b3UoWgX
nQLI51eu+7Jblou1kvsZdxAKb175ZBJmZcn5ny5Wpwt2bivuzveNH0KIn2JiJCLep5GVMqgFXDjk
lvYJmgSwh9D4r/c8NsVgBySYVWi6QrtWW+u8AWdoalhMLBRXyvUv0u2ME4DWXMzVjt1R9XDEOHPq
7z4C/eZqo/dRFUWjX1eR7wJTyDGx9ClnMcP8FUMsVILFOe1v3eNDNfCyrYTlOcTJjppssb1CuQHH
o+PsacEz/Kwif+tRPbAujwlyhTM/iq39qmosLKS9GnH0MrApLBNf41ZeClFZr1bzTZWWnVj+juXC
Yd3S+qIOKPqlJMj85kB+xzrhFNbojjQlSHhiP/Na4W+MAsSZFPXoBAh+K4YhWH04JamVkGmwaCqq
2Z7E+W9Lva2CbzEnyEvybtWCag1XvrVUFs1HpatWFC2mw+14vvRRr0K9Qh1lYOG2J9oc0lsH42Bx
+7gPMoWjyao1ff1K/3UDc1r3AcDT2rmHjWLJfquaV1BCVHES7DnCJRuyzi4+BLkGEA2/Qd5eyyOZ
vvF7cXwz/U3PnFGHWzc8kSOz3qjbceED8umaUwmjdFeqQOgytd/PogBzeFnEKZprKj0jJILj4leC
XTbEo9EuVAHpJqiHZOV/Un3/Xak6svZ0k2Eq7qT4OX3gr4nteTUVVb854XgcpSPbLNmI3avvgwII
o004HT2DGo2adSJzE3n+Nm6EDHpfElt02hs5QAUY/ZFclovmU0stdH8qDwoQK+SyUN3svlCGfGZP
em/+H4DiaIz8w/pcPsrgvrmFnGqxSLZtGfM0DuD4MidmOmDspm3DISjSawlXupw4qR1Oyeq62/l8
7IuqRrqdYE2WWo3egYFnWmCMvRNb7g+r2sovkKzkyb2gp4mpr4lI7MqWCz94tEX/SEvqAgsQAIhd
48qaFe/5xo3XO1RVi+DMLqF64muOajyi5nVVu6tKf9fTiF+n2xpZc3D7PYQFtp7ErNLxk1VY7uR9
f56ClW9/sfzI3lKKjW/dM7ErZirlJi04JVFftIrcgwqLUSdYUHoFxWj3W+GROyAAV7kzFq6RzbC4
oAplI42VVU2ho1Dcc1cPRhu9d2D/STGyGL+Sxdxv+OODawqFF/IJg/uLaW7jZA+WEC6e4wbDX98a
ITOiVfPHsAVS+z4hIyA7VgZuaO9XZT8KjvR0oJRDJJszC97kKeyD1/HqSND7CBIk8/mhJVVyTYhv
33hYwAa5YGuUAEWI2pEjwkSaOPm8xb+l08TRhLrPeZs9cNtqEwKFs262H7J3F3He8KvekpXViDWn
HHdc47wkP/vxhm2ZNwIUnCBUuQf3eswOJB+q70dHTSDR+cpnuZY2EV8ZxricNFyqbC0nO1Pyqr0M
V29ArtU5ZPkOOITCbuWnl5vx8cc3amt2mnANXrhCVApYMZC65ye8kUT1AXMZ4+j0gpcV2wiCptE6
HIc1y9gY6qWN3ZQ+zmJ3cSHhQYgrUZ7dgD3h5Y58gpzy6O6uE17T2Idlv0nLNJLNSFKOoHFCs2vi
V/7NFkCfSuUOAkJ0o5ZtRjwhyXno+0TBV2SQNPcxuVlg/ISduoLggTg4iYO1epMSNvs4VtJr4HTB
FQ9bOqmdyk6oyWBMYD6AiLZN+UkyPIs7tUPrLpiHRLEYXkO2RizJX3VXhROGIiVWmmj/rSUbb/h6
ePSCXkjfg268oIPcN6wZbX3z1vF9jNM6MU5+r3cvzpyd+rOELRZe09G4vEkvc124I6dClyVMn6PD
3smqbpUPdtmMOwYvtRGqJ6dRjb/tNicTIUdOMUQ+q8oficsmpbmJxRRZVn50sRfEoCW5fcsrKaPo
4eIHGRQpz2OJ/q4YzAxa5FGdMfyY+bL/IPFtynlj7G4Ui6yuqwcAm0wJ8xfOuaY90xwR2IGGG8ZW
L/FL4+3ocTATCQEw1Mho0sSJ+OhkgYZ9jDAegAJgSxt10e+3lW9fHEO7LtZvwM/VirbrSbbjZrlj
XZ181ta/oAeI4wOF03ie2OoT33OzpcjEbvDfRwP2Q7ntFPyUDbBPi8pHhRoEnaQWrm6aps0Fu9CM
yWPKNwsv8xIfGo6nSX+3P60uEx4mG4XqLSEcAsB01t8tYTQBk/AnsbgT60RRKexrgRlEY/iaI7wc
ylAGjCDZMEvv8cRt6Rk0bkwgu3XBNlQu/p473wM0zGgECea76VmZyvmw0sOIXxrxNkhfciPTzYb9
Lg4Ih04SpESMQuQwxgmhz0xH4ItiaikZv69j0fDjDli/oT/brL8obe+I+eVlvUvW/dbDiUsdyGRP
QuMRXBVssBnsc+XGnhETzHVC80q4/RQwHsBeOxUJAmxpDFIl8jrVLBf+tNfABYXe7B/1IaXHfzDa
/peRA5AwQ0WqsZiXrWc7jpevBbGEA+JoOQ9dlhrAUVZqSLIOXFb8/CZiVRU77HAdpGeW4Yb5ZfQL
nrBN5Ls3QOigNYdruHSW2GeZs/5DauMcsOCJZe0W/tmekq7DGlfmmpHB7bW/a7/gjQqrR8yDr32W
qOKkhPLpGujmMO+qNypD2HXBkI6X6jIMeWZI2AJ5ZjKEWHmnVrzJWIhf0pKsHbaf9/djUuHtYMh1
+hEpvZRSDUVDeJindPwkzcZI6zlJy6LtxbDLdCWn7DxG2NWtK+DqbV2TR6ToRFHDINI5c54ryymT
luioTXYftTocffyI/mgLSxIRp5/JbZCIT+qE8MkEUgue/D9zA0HMa/tmXRkq089CflKrfnM7hbD5
MUdkcHgta4rRc18o+vYTpUNu2Jel0lutNtfMyc1c2wGk4xtDgtx9Vx6KrKfhQ7jmpOshRW9kVVEx
QZQ5eb522KR2n2fGGCJS4+917Tl7/MN7ajgT7j6nY1KigFxNBuIIx0OCOnzcOAhIczEh767vHku9
h0SjfUHmYiyn/7/N4vYa/xB1IaD2bxrsTCWhZM+j9UqAPl9nILipHimKY6KQLFxoY5yo7o9VsLVD
dh95ADh7e2vGVk4P3YO01rlQLGDZB8xCSgZKB8w27cBhgS7QR6MFJqqXNV8DOj32maKxjPcHw74T
adutbumlM07G3wPEMAoejVsUJ4Sks/3O3TYY70oy+RrItkZ48JZydIq3M6Krc0dWSgkHQHl136mX
4UTjTWdgGCUZHY74ltn/UdDaLX97C/Kmk/C4CwI7NK50JiUOF7GSofvVPo5HEnCd78jIkX8sXpRZ
7/txpWA43JKGj195906Ljeo4bB9QBFRynH77x14WEA0eOzpMiZCUlpbr4LTuPqzVVPvpcsGjjXGW
tJFALSGuKmC0xBRpjnSgrwCKXGcflVES9dfBz9xs5uM5ablYQBJ0I8k7rnvi4Dw3V2XO6tt4VF1Q
vzRK31VXAGUOZZACEr3xVTMK4kv+vrB8F8IFjPV9Wn5V6ycid9AFVJ4nII2i1rpYkQbNbahrtmW/
/nKTpyaWMyxSDtoQrX7GBV8ZAS3ZFWkw18GH6p1erzC8j18FFXdI73htkrpmHLKDNWPflF2n9gsK
0lTvj/eonolW1LjL9wmr9hODRY8CJkQgqGsa3fJupDbzUt8A7jHe6NyAyGA81PPIqIVav+2p8pcu
5vPna+De68fQAQkyk5bWV1IAakyBBLTkUyLi2KYe58k/MssjgNveorsYgqST//S4maXd104EQghy
2CXmRkXfmWkDJvaVKs9zuDt8wIlBU9fs/7c67EnDUyQRhxs2jfKoMGuCInqMcwzAvWZ55gGqW4/Y
qskb0eR8Jzjuukd4ZoEd6dYwKacnwE5NTL8VbKYDuku3iIGXq7ZcAULBp9yaK0RV8MUzPwqLB1OQ
aYNPt4CVLAoZGyyjwZ3Uc6Qn7aDApsidnzm4GfIqGalAaJHkaqEctKySWfRMIwiepoYQPA0/DjzL
MrzgnoCcbAgUAY6BSbQk5G7vdl97xv7Q21ljB9SI7ux29HlYhav8qYaIIudyaOYgyMOs+uYmBMFM
EyWkFt8TJmkz74wzmqeBlYVsa5cHWA8oue8G5pa6k1Piwmzr84/KtQtC0qxQou/KM+Iyd/d/r/K6
a2YkEl5y1TRNaDnWK6pEeDOw8Xz4DBk8kbbtjT6YlAT9zc43+vsZK2DiLeQ8KIzIg1tqfehgnvv8
wle3Aze9/+imvfHF47Tk4wuuW2v9wzwYiYC9ml38YJ+LyzyrrO2IWNB2S7jqSC6+OVytaWfPBUVG
a9kCA19a63TG0AwcDMKkPQqxp0o2AvrgiBtY1QqwcxyWSriNL1mQHyZO0NkKZbIjD1oSR2qPAXkF
pYRR0kjNTqZ36XDvz/QzoisFr8+oWvpeXFAOwnEbENYq84HTezHAREeKhOnXDshTwjbLyJJCSyBh
YoW7NstyJN/W8VN1mm2Psi43EpwxFYf1Z7eCTpBwGLTwfosI14gwCUBXjt2seveehi+aFUJ5Wsoh
zeMfhyMkY+mjg6/7km7geCtYMwPyO3JhzOi5vVb/kJC6ESxvanDQuwq9q9Mu/pG9LvEXRlMj9CLO
bKPyhF5igCoco0fExDWzW37PMXUj+p/vVNncE6nNo9ACmynDlgARkIccMMaJQNyr+qdig6vou7bF
8ACtD8OgbogFANlU0imctS9zq+f0f6Mu4WCcHHfRzyQhv+4fgE4jVTNCdVP7YvsG8nr/bAOftcig
4as0mwbr2Fe4FUEtoQDiu9uTIQjQBAhl5Jz6H63tsjmP9paQK3RS1+X4rqMdUOBOYlxxWgazneMh
nQdE7OiHCrvQwdAwuS7pI6Ci+VoMkL26fj3tKADJBUSm0wUc1IraxkGKunKNsVClgdJ7LJsj35LC
cLcjTWGX9+GgOA5jt1FTfbtp1HtDVjFcQW9UjzyrcxwyAFxpNnBhvNmXx/A4TRutWIfKcQ1Z55tR
FUA1Ib1haNA7Yhndkw71fBaM6BC6OJqH3sUHz8QqtNSR+EwZphrsOXgPaSzJGSUJQ6UMZi7864GR
STCm5BlcevH51G8oFSR6mYn4ZK2TEa81QDIneJw52/ryQjR0xY8zE6Zt8apI6e0zG4v2melkFWsG
jMPcE6lLtDA+HEboGCnOFkexjJCHsP/NSFMN+OGfVMydEIVtw8gLIh9ppowSV5jwSHY19t2LJwZT
Eh2mqA5Pr4US2vYGh+8Xav8i2KpuHB6sdhGcd3hgGRXjAAD7GVWrsillCjxAlcOaNXwYgcOdlwzM
zSPbvI+NY+wa95ysfrwxwLxj5NrU9GGS5jrk/XMIE4FeGwXImbbv7mZp1/iFKELeaN+CyS9zqeMZ
nNj0ej+JWfWBAv5fP3rCJP4vixC4AGOEME70o6FiZr+MwdcKb0gaSs3szp0cnsjQ09s+PX9FC1/d
KNITjETOvRrL6olSYheuoR4sNE3z8rs1rZAsbFoi4/b3je2NFaP3xb/OhGRvNwyDqMGhC070+pwh
lT4Jv1CwaKxOyOwvBaIasfim7lYpbGvPxnEROpZTdXWwdr0cLFrcROtc3Rah2jENRye6nfJ/m2zK
FLE6flMKk5rlF7FJ5HXs0eyFVsTk8trKBmDLTQIx7v7HVO01v5xAjpNJDoL7w4QOJJi8nV5VkHDB
uyygRvaTe7NvqcT1hpaJhJ4g2gxwwVOUCYxj5QYcA2Pld4CiFd9kdyseUveOHSRHgd1OLnfJ6jnJ
hALekmXpjlhlUHTArQkTNuREnauyGSUuZagMnqqvrJT/AZ3cJeI/LjGeFBg1dbaz5KuShGrWDXjw
0STdoZcCeac3u6As3+2fkbnzbPPN5tFwOyouSHNGttpAP5VUzGstup4pu+pneeyqrVSVXwYK3Hec
mSdhXNDuLcqVTiUGccnpB8v1FHg6hJ3LRZ8WEeoMoFV9/Ubw0TNFWJ0KQK+HapJB7ztnu4SZ8wAE
2OKA2bY2Av59IVmV9qbYzsqFbAMe8DMpk7jylw70SLHLLE3/5qAZqdzVEVkQpZY10cs2ZFqwSuEA
S89g/KOI5y5038wG8+kgiEHMiFTJ+a7MIyI0IcV02snGk79ClnPVTNcNeK+iaSzEwp3h5AdUqYOO
w1WVqZLdXBTSsnUnGmmpQXNJ98+LLZ3f365qy5J7+2+xSnAZFK5QGQyidBPwzSDHnFX2Fixpmh4p
i8Pyo2gL/9N6UHiQ4lkgVH/0ovIuCYGWMvaR4VrDm5BMe0ahe88RW/LdjuVOzyVVjDxfFXAcv1YQ
y/N3TTBEuzJzE/lzaoB/ZbvugtAp40VSAcAgU0mbW7OHhVr+aw2hiMMZlyzHldGeLrROdBj9/Mck
lN6CnnQxagRnU6MFClsD+cM+hWCcm2wYSCUhoxuAOd7j2uu5DaZXSP7d57qpbhoaQo34OfiRi3mL
llFdxIw4YiYrZ1rEC1fW/YEWp7XFbbdScGkAwfb96tAg36DdW23bWK9sxiGHTDe7lOe4YJhlnHrb
ykaspZfPrHz+8kdERuE+iTNj/h32Z0OcCNs5tptNpqArUfKHMoNsCX+fq/YJikzKKadYXAl3GJCM
BpkkoAJZQNUN+5hopzfLjaV0twOFnvNNnykFkvCwMHlBmCrTnZcgakGf3LCIRP4GeVSRK8fAMotM
27vtCYgVPnM5sNo3/fG4nkFDlD/+QVMBCRCt1ag4yMtqLTwwlbHD2YZB/TbXyEamBoD/N4UU9LtV
MFq/m825Auj0LdVv65k81FNgfEdPPoqsT1rE8NP/16kGSoX3/E83Eers6FVqNqWq8mW6IGNFE9nv
Z7QdvI38A7wV+QcLzN8P7CkrYkP32Vrw4s2Tj2MY+zwBtNCnK1HmYlUnZt2vHn/+EQ/FqKsQOtsW
y67vuKM7ytuzAWkUQsguRqsvkXFSf+uKuEXycNmdbsQHn6XOHpBhdDXioTgDZukmc+Vcp8GlV/kF
QTrMPql0TB1K28wXsc84EiLm0Hf4qt1ubYh0GE3e24yHbUhD1G+OIjmQmrBRqMhBM8dijJ2ssBLT
BvsFlGHEjTaB2wXn/obzKsPwcOJgATqe2vPiAJwffFW54iDMpPStHO5RcjFAxyvEpJur/ZUASrv5
EuxJtcpd+55pv7XpYQdRt6cvvBBHS4mQu3jemPZ348cj37jjYdDLDZnTt7vyAwAoofezJC56rrDy
9y9m6jOWF4nw3vaxogEsfs+hK8BCcX/y2TutpSSUCNhZNoFTopsfusUt2TnnKXs10brlVySAEsT+
YQ9jZjD5pl2p+AUhAxvHQcHc9K1T4vfq/BmswgsN4sm+Yopp2E+OULfPJ2zMJySiPV24cN0hsftg
NinKjLbXQUeGFhxS0r+3JcInFMV0wub0TzIaO/o4X/LOGEFbPhEfymSQZUg5ygVp/6LuLzQJVGrl
xn0ctwuBTPLydJQx6ROhzWr/ncXIFQnsshmelNf6+UByo21qE+reYaRFPtG0snULgt3qyODbqF6B
weknzFc2CnKqxFtGc++jlyfQ2BeOIMYTB5bsovIcYNnw9xF+W2zaZISttQuUOmxDWju3FxXQqnO1
fyY3z25XHjSJQJpA0o2ay3dd8maKg9uzbgQdfxfx2rvVqKKG27EMukAVT0qR2Yozgpdwa2ztthb3
Dt5dnRsthcIJrzQeDYlLmo5BS/y1H2ZalMO7URsvksOJLwDkv6QtmfHl4rokzXjFSnQGuWKIlW1H
qlicICbcqJQq+/omLpOeo0RdS1SVlNNH82YtE2NAC3B2Ds26sXRJAjpUmmmy05nbOtgApqOfy5r1
KqnavMlXwIDa+JVS31ydKWzu4btUH8O3akMXDSmupA5lTIyizqr5uVNvTIFPupYaGK4mqfYwP2bc
EhpqsQHDfS/g9cu1wLY7lBk9LrXrV2CriH3t+t8RuqP6z/m7jVrvUxI+nXPlDHmrJ29ChGHYOeXt
4z7kltB2Qzf9pm5vTIuZQHOOMgEd/ZDcyICj/LLNDz4sOfRvHPbcqiEPvPGxAOe1cG6gVH+cd8dX
Ubf3DkjM3i9VH6DKvpOhR2hbN3vF5mMxO+5GyIEvOILuk0hfSZsj2reyrCHUtS4jiNkZ4WZ5G7o8
SLHJ7tdPHLY02CR46NdWZnmwjPCrYW+tKLf3ZDjXhK7rwUsuI/p7HjVz4iXVi/HYeK9u6A1dzkfs
a1sEPr9TUhSS0rYhcDop5R41f9bXE5QAbyCGXyq9U7xv2IdCV+m79Z2aj7rOu7tpLsPPmmZrWdDr
dY+acV0knUpINh0IbMtyV1h8ITHzhvFFNGw5tfY3rINXe11zzC8LPvrG3I28Zd7s1e23K10ttGVl
hn+lp883bN+ICMBANRTbC8E+fWLBTOFmwQTiBro8UhcLjfMETsn3nHLeYPxXIBGRiC2PsijwVXF3
irfvpGXYDpnCRCSCzE6qqDubcc5anEICF7MOkzNHYg13/Plgjs8hRWXqI7qZDwM8mGmVBWgvd46s
4w517BsF2rCHlmT5dg4OJFg5s+3NhubhQ9spfRvZ4P2g5OuefEMT2SJ+QO9DwIRmBvTpDIyMXyGl
DthDK5mp4NJal8htSw9jftXW0E5ei/Nu9vbnqsVMYAz8BDj4noq51MP5qGfqN+g1LGLydEGjTFdQ
4O4xdnNMVZjJ3zwjcxk/ddHKh389175iowH9xv2MPbSxPIDlO1tB8V17oVw90WBFL2c2XUtGofu+
rPyJhaY6EZOWPuK0CNbUyulS8q003orheEp7lUIBLAsRinUH/7FSrDbvXRaypxEIZGf4HPeaiwCR
iB2BQ2Ridx11SP9Rz0IFvi4KPxf1FdVdyqjsAojUOxofVR+CtYzVHIIOBUutB/UQ5dBY8LjgGlGP
fKuvbrPHg7H2M7g1a+J01r+fDh19GnSjA/llyjnibfgla632Z6cnMhT+u3IjYz8WfClvJiAo2K0Z
JYQni9c+p2PDndcCBJA7flEU0PGt1JKLLT3fgHWMqYNyJTsDelRSEVm5G8q0gvpORhpBpkU7ooMs
XoKd5hrg5IjqQNIWB3X3aIcb6Bpk4StTwFIw5ua8GWvbhOUq1Jn5LYmSAwWgCdcidU7ZIfUjLKn+
daMHZWQ14PeOL91NpsXdtChl1Qiu1kxbYNhNa//hblroZTsmtcsi51QoqGdU/6Wm4SP5Vu5SwakU
PFDDFuI/qqy8pWeSgbCBwIX4VpvTRBPvlZtNjPA6pnc3jz8dhBERdvVe+W0TnrOVferCVSUrc7Cc
dJV69SKwSymNUDRL95JSnrBhE0G0rCtb/fKxzSgxgBcMlcrPSRguyJAHFKyVWr+jy8GvQXPPbOWC
g5VXYTjgpCZDJb/4/g4Mx+VzwEwAJUU7v7b1WFBvVwloZMoKIve3qvMy/pWI5qM61R2vZZdV2R5b
C3uAw6pJx/EEgGyUy6bWdXd+m/nvB9MMUl+cPdyv39irUSufRVStYZzf71S9UU9AcP6sGUtA2XlC
MzSneVevVL780nwCcYb0zWsOVa7W7Dh6uHbJ70URlfuE1A7APpI4ZG0b1XhsJ28bU/xaI+WgHs3e
z0kzPK+an+Eatu2xaJgDEUf/ztMxsBaKggfa7rvXW8qfkjLelrCi50zt0kcFYw1OVuXcwSFxYe+9
gtXvasyyx6AZWoWgyiyTJrS1Xuzk/AW6OFEnI6pGtL402AfpEV528+ER2VmJAtN1Ri7gByGBPrOg
Lyc38SBwmeZnDnDwLHtb8wG/waKqoZxDDlT7OigWEHWLI90Mmpb2QqlK43ZMsqKoP5zG6ALBDxxK
GkD1Jf8mirIuSXBKWhHIUYObpvjGDq2TNOxFC4HvSyFQL0kTc6G26/QERmneuX+ccoR0zUTmSvl9
XfLaqB+pKU0hxSBbZPnJcxaPralmw10w6zTgMCnYD1gZz5lN3V2AcGILNQO4N0rblGtompjcQwnS
KlMTzEFGqs8CgEGQeQ3qWdZhKkCJ6YWI6JWkaqd0K+uvxe4e3S51GAlALivI7Etli3Sfq5aMd1xc
3P1EyR+XpEzqSrOApv093fy24vg/gy2lWtYE+tenwtTd3SZ81HCVkGxJCyMaOFfC/sr/L3lDP4NH
wzqdzIjTfeF86ooMmnhBn5O8/6LcdM017V/43iuTecGSaSTM2GVw5NNPN5w1tFA2b1jxKhueDuCT
A0cH8WTSXjuKT9tokTYC2AjjPuVekX6Yb2f58oUK3quNq0VG/oOcnfx6/AWXHEQWZBMGtmFFDOt0
LCRJUDhxCukknZ4rUhKr7LMKZWoR/ZACFySspVINeysdA/yKmzrF592LvhGqplA3bm8ucma8qrfB
BR7AuZ/ohX3sntUa3A2BJgdastO+iPZCmhWHQ+eutvyqrcAbVPB5PNRHpVXOhqDhohNllZPqZ8PV
g+2CJomkK977C5gWFQSDtw8ICMAG93f4D732AvwlrPx2lVegKT7T7+yLAIWyD6fKZRaNzCegDYA0
kydlqrZbr/W94rA8x2QaOOWv349QuLaacnNFKHyNFERK1Fjn68IozMjRtczyTO64JGqMXDKZZkLe
2xfcz7D6kXiaby6nWDc0JgZFG4JJ8+IvuQXPnMdPCfTLSIsCaQJLEPQNsGNqgFhz0FXX4cAne6c3
4BqYgkD2SvSJ38EluuiNw48oINeQQP5KdOuKBysm56bXqfUFE5urLbrnby2pYafEk3gH9PnRrhmh
NK3QUu6T2C9mA7okYjoOTNSiPeuC95JYdwAbwkWT4/trZm9XJnPqavpEqR7Z5LiYkdbYTAycp6NO
JZgiNiVt5+6ZFG5S2rtSBmClqxsFbT9tiRQNyc4nr3Sxz6+BWY0mD6ru5j3MW/G9Cf7ADEqQ+GpY
Vcx9TStUuwPu9yDBwn5E6ZWKvY80amOeMwyLcCbMrcfKEEkgzVQ2rj5UDWQLki5gmMRLR/Z/h4Py
0SdDxKcelS0xRYDy54d8BXQPAu7XZ4c5rjNobya7Jmh8zE6iPrnaREvR7P7Q5klKtXsXC6snte0b
s4Guif1b2fr7vUOe+2YT+bGmnH4HD2qn0f58ez4az1yfz0TkXDjCSefV8FOROjHN3Jkr8OxVd6Ie
Nmwg3yijFLYEgX95to0/e/ZvZaSnv82flNgeR49KmcsxTlRuvIg2m3/4h6WV35+P0WteM3WuEZZK
g58FC+9BUhKpP9NeNqwQiq0ES7toY0TsPvhCPVIJngHHMDySBCOeTkcbYvUMmanjk3zfYAR6E69Y
dhmy+BrzQFhzrGov6fSbkKFFxE/FwmaxgCKRKMLEh0dFGrpMaaTJNoqWKMxoCYspcHL7/JCI5SUh
9AUuSopk9i/Pxc2Ucn5/UXcokAcnVwU4JEBWaQ8Tm4RLZ3xLSrrryxUG8jrzA9yiYLon/0570aQQ
4t0mcrlsLvu/OisAZW8TDIJaHMnNTVxBUW8T3drz+f6trS4LQ9KbY61/AqviCCHPNxGEGyqOiF91
fYJ8XeKsW4F/w+f4hUiELJgtyuXuJijc1xHKR7puytjZP78ZNYPkFWR4agH6qJilSXQ01/yUtoRa
KYgCevAM5ebZbZ32caacwxws7DZEziyxFKjaT6YzwwtYDSzbtJZlumQYCg9br+pnXpdf6pRkC6oj
VuDGUFjyC57tCB87I+ZA13CmoYsMKvBvZPtjiL1s6lYnNdZUU6Qsbojq2xCn6i+gnLW6QVH/1D0V
LhYiMN1TqEaxZKRdF7o3fkg9vzfX4JdCx5VD2S1VjBvK/dj6Z4s7oORw9eP1iLgFb+WomAm9J0fy
jsFZ7LdSRTYKWRPfG5yQi9KtuuZiSlv64t+RprcBxGjJgCPOqgVYWfFjNxaI/T6iUmnSs2rqFN8g
hRuY7VtakKnp7g8EKh60XK1jPwiIrKKhOjMSajZWXBP/LuI+mLr13jt2KdLj58+BDm/NXyKyEsOF
NtAKrcMj4+ZgKdUHq3My5fXbikrEatiohicU8QHJf3d7z6SUEtKIYwiveH58PV24DrSsueTAb8xg
M/V1Cs8zIFTZtQFdvBjtqdbF9gMCURT/u5eAhCpJDaUYopcLXTH7V1LojMx0fJUgLglSAa8/lgap
TddoTse1d9ISC2AFzJVNYfY/Xg0VH1xtzUlM0e+ELNIAzSGtnXmiR4d66gvreZCXAD4TusKxt1qv
kptLbYatEtYRvhJnYl5W9tpfgMV0ejWRFF3Q8KZ0VO63U/e6b9Fk2S5Vwn68T8kgPsrBYQDdrU4H
CmlYPuIJnGwRUEIDVDYZftBWBr4BSDMF8gztad6LNn4yrfXyk9rHVx7ALmBMA3XGkdpb/bcXNRoc
srDUBZw7fTWJYiIYS7iwg33SNCXBfsPDgm+WPsjCGZQg43l8tpVWpQETGsaH3DjYrW2mVPPJcFhl
gndOGyGDBN32yP2j9g/yH9Clsk9cJz17J8FM5s/wg6PuwEVM/awLz1XA6RijvyTBZy76Q90zSGSy
3bPHZlwjsD0TP5zcWRCqAX7HAdcnd/N+XbhA/YWkIwb6vwDu98e1T9CYqQB1EFJAwbacMuffhtPh
GqNLO2COxO+aoY0UeMHkp6NeHPOic7T5qN0bRLrfyAvuAmsUXunIbTnw6JBF3kzfBR/cEoUtkHRE
NrL+oMkFjCniI4lXFbzQX4FYwLkxkLT4SbDUn1Ykx3sHRgE21P1l1rxgLhjW8iReejB2+ko17lfx
fbHWjvEVLnEuE7gSOHmLC3cU4suTSdlP5RiFjgED9+Qq/tdSpZVV6L2WJtfbxGKZQWnloIQ17e9I
VlNCqVRoHkAzuGoXNPjov5yrq6dAXVNTXEcMIeG6XAi/mzwxew4g8NAAV5zsFxtHFoWGYToM3rdt
xsQdfxmy9wMmAK690w91gQm0T8q3n19R2HitZMRW3St6AA11itDdvEQDSQzPM08wqdv3SCNVkNhG
+gM8o2tsMTU7HJZmrMVf2qbcukSjLJEcLcEW5+m9mp8+R4XRP3/N6Qnk0HYd7KY5x8WQgPKCMwLJ
GqH9dLZIfPqf42XxImji3Bq4iiXzwHjXGerdTRqZ2fGB72Krt/i+DRTr1tH2B4LUxy/dToRxOAI/
dcQ2Mt78TOloAEE7BCbYtn4EQINohyMZFZ99ByGTRlfkS4G34isHGnEwj6GGB89IpFVBD0tOq6kh
SBoincAaMetbjusTNwPRkIbp0951m72DkMojkq/Q0FbejjFyiZ5vh7rjzk/Yz2qes9IfiKNmmMdm
xwYd0Zkn/mYRNfkcrQRlSfQtZSZ1cXhIT/Af5DtmqS7Q+2pyv1jdg3DYrFHMW/SaRiQtHVSxvKXy
Hmd5c9aARAON1QElI858Tg0Hqh60CyXmNP/pKaJ9qNyjDAzWHcIo4y8OA7CD+JGUoEOtJ+tZC/2R
1U1v1j7qAoYC9kSYeX1N7xRa69wYECkpo3qtlGwogemBJmJiUDeEyPruSvYLMTqTrqs8Ksi7NYgR
OoOErTKoWGEuaD1YX26JvAH5RZeImaxE77zDtW9AMLu8WPBiz1vmRoWvOjtpHh7wii6NK8dEUo0l
/qR2HoUtdFS9lpEXaJ7XeLoHOvmbV5mu7yjZPyKSt6eqJYUHwqcMPWYzULFfWkzKCISGFf4+9pch
fQH+oPVH28gJziGXR7NjJPDGzIkiwRDF5FOqofYIyMsrp3X899vaf/+I/lS3Nx6zAJVUMdhDQMOV
qDlhEjlbeOAj+1LSKuPkwfBmWBSBv2N3EymnEq1VzMp5Zcgq8272/WWwQzPjtstk3l+VLFgvKa3T
oBefMuhcgtH+LT51jKyQIbzzOyHG3ZWsuULcWYOs376xC6GassXommFZ7KnzPOvqRHv2ACYRxt4V
rgmL8uAIKoVcHwZ3vXyvpToRKbP9ro+oJPCIsQ79y/Ip+oHRtpOsTXts8NTfHVo0mZ1udtbU5M8u
FB1+cI36a5hIxEcA9ArPmLvxWdVK1Edudp1Mcq0FWYMvomYKqUWY1411i2lgblwNWjyRSDubKDXT
B/5XRC4ctFuT4RYkjVApNYndTFDGZOE5wx87KJ/MVkq5+cPC9U8HfE6pWv1BeZeCBF9NJLlRSkWg
1PYKqGIsywj8QKVJCZOkRgyuYiqm4nzSCJnl+BWqJ1GqTeDR1c9qxStRGgOQuNlvIL2Nk0zlvXL6
0XPfNaxg3RlMACsv78KrINNoq9O6kGvAKqcjo0SMHKuhUTMSIWqMnI1SOdZRi1FV1yC1Vdi9Z5Kn
yFHFnLE7n3akJw7Ekwea4HyO4bYq7J+GqZ42chWCgbyvcK/kZ3DuBolgqZJAcfkt8jsjgjWtBXIK
Yx6MwGcGUhSO5prIDNx20Q3/og3VOsSpjvPMQe3wLv9bX5Ib3LzbhBZRuvgv9W/9ZLganVBjVIgS
er2ojyCFqESA8VwT+3Cni5PEHjtmGOjKIOB1DxJoM3m6oq971SDt/Hjn/Ha50h+/S0GwRD2MEent
SpLuIlAXN2ij1C14WmKS3wFLKKzKaueCYQ2ltRfxoV4dgPFIYpXNzH5cqjtsi6xFcvUp9MLewN0v
RpqhJno2C89j6ATUbeJaGms5/dPFNxpFWjnHepxPcV7bCDUnwMMfxvpI8pRJS9167/RkHlhcDPxB
ypxNHiGlzHk7zTwT0AjihKpYiJUbQ2512f4wdVn87XVqelw3P5cDae0SMsQz0zRbeu56e+M4KZET
UmYQLETrJeionont/bN9gwS3LUUmo3KdM8kquaszRf1BaDtBoRRVLnZ4ozCRvd8irrIhjqqjj0ju
rdIZ0PRxdZ9na2Uf3sa6cNFREpEP0klhA6aN9Jwg8Y9r7H8USRH2uNOnAnec54ztrv+BpzAGj0ID
XpaSK6DYQaeAsCOFsXvyLeKvsIQqbPBwCMUGi6wwBMvhgWIc8QZVJSWvz9Z8IukdWaI3WIqIgln2
C5GQrql5EuqYhqgFSL/BoBiNPugcMD6sC8YAHqZybzVHzAtFc32quTenDa3mgXMRdoitGnDpLzRU
6kT9s8G7jsi100Jw0+ZenOtC9TjimaEcJF64Jaf3flAKIk+GOQiX3bO2OOoqBACnN1/M9yrR4rtM
Aoua9kgtyDkO4h2LMTkyraK7NgyUjlw/oWwSW36veXGn5IuXWtc5R8cgsd52kHItY2MZandZYBLU
dn8awFuZwUa1fOgQP5bvaW+YKGWtzEJFirnrzt8ORB7ue8Y0sfFJKOshlLJg/J8sL0IMQiJekNH8
Rv4SGEynzJieVAR83YliLO2PZFWms56TVjq+2VLEH7g12i4Sr0WJxmodo+NiSFX34OV9OoLFJLVx
0XjMaB8Fr0HGsYw7uKQj2wV21Nd1YtqSkvIcqYK+RLEwkliTiHHxaxrh22/ElvTuUpkRiz/QGX4S
XX+HiVO5DqXO+F6DaPT62EG6IiWkaPfcdLF3hNGF9PSQ0FMzssNJMqC6Exz3o8Uaqa+KubDICabF
gTlU9TNJi7gd2DLr+Lx0idEGINJ8EfqEy20O+Pj2VlVeUqdl/dax7uIV00lkP/onPLlKokoVT8vq
eRNyYoADtQIrrJZWJIP6JLI0YOc/vBDUqu4hsdiMP4+QLMpbmq5xWLXtflVzdzy1QrY65fpZ/tEb
8Waxcjjz5UdeJVWGd2gV54HYWk2dVr+bjnKQDzNVQ4NkpH+4FOaOi9PG40ltZlsQDy4lkz/IUEKV
qhxoQqQg5wrKu0taURdpXw1qJKzJ3jKMLtijZvpB72OdIOi+T/q/Odqrrq+48SEr89ijj1kLpNPs
+s9Sw1TmYtBks60N9sj2a4B2JrtUGR91Qo04a4U+ZTOHcN4wO+D0Gzzsc8UdwoTYArUN9f11a+TL
zrp4bYsy+DNak1Bp2rLOCiqxroYweAsHvg489ErBuxPC2oWGlZJ0SInqMYDLnCbxUkConNeurHZ2
ACC+36U1SAw8XbjUfkSi8RN9YJ0b5Evg7+44kUvdysntbUxz4RTDBB/dKhGS3f5/sOh2I9eeFWqO
ZYpMs7TH8e9wUkE9YB3Fgj4wz5XV/r2TjZP6CJSMJZduJxAwD6GL9pYhw6rffuI5KXpl9Czt0vB9
Axl392J7nwtjiQQ8+ref9jz/rSsoiQD0rMqA2kAhh6qRq8qJUtEbxr30c3fMQA6lnkwLe+yf8lbA
b/c52VGbQ6AMvADIZqI7nOW1pVijueypGJa0c4m9sQFGBMJl97qw7X3mcg5RmcKq7NYsciVvE4S2
wXaweIw79ZswA1zCHoJn3VBeDi5w4NkkGdTS3fdekByd9ybgyxYYil1XIRCgEScsa2DG0Wmezc+g
o4hfGckMvuu7H4kikj5qUdsIEZkj5jBEcy24dfm6AHCvns6vbqDPZu6VUUONcAoVdLSVeAeyRsgC
ejJGdalxdZB2diMQ+uuDl41oQbI1jEEA8SAIBBIOPBUUhEw746WGrYh+G3l7d4htx2c6PjrzNHr7
CKnIzeod/klV6Cij73yfN9KUTeky2VZMty7ujG68G7Yi5msBQMdnGQ64fm0IQQV/3P9fLxoZ2YY7
7LGVHihWlxn6LMAC90q/y+eRSJ0b9/y2WOQUU1wuPF72706xcEkwdgWcupbdm6xr3nIX/S0nAQf6
3TFrTMY/9dzYLA3RZhARAECR0CqNzsF6H/PgtvWHZZqbsz76vx5K53K3Ufosxbb64eW41p37z0Y0
deiS6KOM58BaIUaJm1BxhPZzbSZWLBYNMFZyHDHPN5OB2zkJCJqZcQstmAe/ykiKUiD+FLfbFUS+
5ODcBtNfj99kVzojqbaq6htNSrIpuwJXW3zcdk6H5dZaIVbXmwdPuwhzy795wibH7gs0J2Kgnwso
UFJ5VI2B6HjPWLofJQc3D8dMWJkqI7BeZm46OWBCfWWMEuoqehPVEtvkA5zz5826OWn63Yeb/4Be
jltD6Jd0KCkaA5Sby+45jVOZxx236oqoueSmxQYZiWrQ/Bw7+dmxG7kwMY9A1jpU0Wt5uMQSFu7c
YF+/3BsBjcdQSd3DuUuZpSC5itELnyYjxSQCr7RheDM8mwV1ZifJ39l1UrD26Ets+4q1jMwofh+H
B3dv60cabN9mZRuYVU8HSTHpVvJ97nyQbE1EQFV1FQujOJnW97wEs5vvQav4Ph0+nUrOEBZJkMnx
1iT5548Z4WMLd5DUIslbA9kZW4t4FTL4JRH89oeItJj7s1dMYpMK4SqHl0E8QCc0GWs95UbYzLKY
AHS8vdA27PLNOeAiigPJUXCP0yRBIa9gi5g+fFo/qvhC1QvxbHxt7v89n6Jc2Uvg488JUZlfj5sI
I5Ny+VP8LvQJ54b27ytN6Uyml/47fZIDzONEApnzZb1NCOs5xkncCh3j8OqbvxC76QRysDwzrjUu
Cd4vcO/SVVT+HR5kQsnLO1ErPZ2pULwYVqqrYlfYMbfJr8QKA6wAH2L8+RDIgEtthGGxhThcHemG
1VGKr87XgiDxTkraKyrPB+qS+y+9Q98dEokRMl9l30/DBw5p11DSAWmP/82KDokTB2vukq+WUC+B
WzlH5Y+ayGogyzGqphTKhrlLNGzN4dZn1Qsu9LWG6ACD3Sa1mQ24hIuS+3K7TcZWCdG9FsDGIqHQ
YdUaDSxyH3MXhNVKim4A1SKoYjNiagD8tDA5Evd1qukCvbt1hMQ0WRXOsULeQMO7rtqb5qTNwcd4
0lWAJWp5XdJplTcANWhPe4t2n5l5ZS9228EwLaVKvzMLUzsyCPIQaIFN/kIirYtqMoLvRnwmJ1qP
5xk5m2+y7ADy8h89+8jpg2E/RGp2qv/+plPtPxxegs1z3QegmG2EJvSzHhLPJfs6O6sMxogmufRC
Mx5RE5WrIwvNyI9SC+rKIL10REaaEvBXSo4aQQgs1JOd9j6rdAVBLJinDbqNA+TnWh3n3Kuw4CKZ
YVWTJ6SxKY0TPA2R0p1BcUizvSCMW/v7Oe0Zci52ZZ/eMZ9AaVL72tYCcW+WJCH4/fVWDLfPts4Z
v2zTB1CpP+9rW3GPDggCUCFXMABqhtCD9kEt02CmRN/LZRthzHtpEDaTBSH7WDkAuFan45WvExbL
cZvgLDlGMail5WOmgqIj61G3rybkw6WJEzzHWThIjh6VzL/wuMcVpwM9DgqbDkYdGAs8/WEsb1Qn
mcLRA29k0dtSQ1mOISTSSGiOGRdbWhGPJMZRgz7P1sTiVjPjovmKHbeIBcSpNjNkXgYC7CtXnT3O
JtuTZblq93ujvGwlDFU1egFWxLU8OgljMSG+HP1fmemp2p0CmIaV2EA3bQewJTeG9HarHK7EGPJm
ZgEzUcuHIqKrfcPiTvFaF0i0jFA7HdPscaPBIMBGuEjuGSt2OD7OVHhrE+K1t085akv85RUZzhNZ
iI//8lfBTf7uiFFqrusVVNN3az8bDGGv56TLO/s3t5KxR/dWhw95pmWuPQLRcly1LGBKdcnxrHMT
ha8KFZrykogjuxr11xI919X5O7+bamWNGpF2ieoEwUKjYTjyu0zenYA7i1lqPktuJGJJpu3jp1/g
Hm+gROccWRVulgiBfdDGUFyYHHI8ZN3dnIkbMd58wh2h6DR3N0iQ21AiR97LDdZFcUHqGm7QnXmZ
7vsqDdfPd0nDVS/ktCkWcgxUWX1uVYbPg34zMp2WUb2dCXYbUKicCyyByoBtCA+eiO5D/q3/AcnG
4T5O/0F7nwyAA/x7jMLJTKtKl42OK3//78hOPNoaaN/RT6NnVZm9DQEay30JmmlgOTMq9+taBsz3
miuiaru5JCovUJMDJ+bHQI9lSn/41wLNXCHLK/AmOyIsCXmjt+wMQbHW9Y6z+5z8dfuESLtTcAc5
kcxpLV/NMdsyPx9XOGRh4OXmLn+Q5MzzVHJMDc+csH3037nQeYxvXIMYj9o+OzTPitu4Gk4FwKkA
4p5YT9e6ARBabWfC9wgr2E9/+KeHht2HukXrhU3YurQCZqOQy5tqUp8jJhehabikmOYQwAl0Mp7W
2gePr7TWCSzZSlY19X8Mqt0uPFDMbb1yuOr36fbxxtciTcwTlvkoaUxXWuIE+FcbXCcqafRJeuYT
T2WLWXI5odGtytml4n87BXIfBrJ32gkeqNMkOhlNXBrMIgMxzN65AAfXQwBznd21K8+zUTtum0dR
UtGMxkKyYLQ+2EI5NC+vbM2c4dM3pFYRPnFRmDzglyXpOOHDDTZaimPYUZ+WtIbC72CoYoN7pzHo
TmuDLwU28S1P0rFQyZO1+L8pLLKIXL4I2L8s+3S6Qol4q5av+I2vuKBbdQKfaBRganGFjr1qO+E0
oUMLAMVBme3JPnY5Ue4F9sCogjFFfJ51300Q8hq5TYxqzy/6ESrwgqW40XN0Gyua9MWpaZSvce/b
z7aoF8Cjyz1Ai7/sbNkbpHyE9y2QYKS6zB8t4EE2gbXWC9/GmZzU0LjaWU+ymtNc/ZFj1h3Rp4HN
/NjFY3m82wSqfjxH+8efrzgwlhMN8AqmQrK0Tb37b9P06XOnMbvVEMp/ycevYRn9bWmiha52E4aE
oy+2awzHwbpjXDyxMjWMFdWQ6v2o4HtdVJ05IeNRV7FEwxOrcwuLXwF6wQHTS5HP2J5sx8hqfosp
catORJ/4Hun33ryYE5qwFcy6tBs7Q5TNgiAMTO6KRPXNewXqT3QIHmFNc4eWvTmLp01xxvCFIZOn
e7bCba3w2B26gQ7TCmOnYwUK5oFcHV5nCnq1W8rT+KIq+fvQ4mgWxwytjRcP/Glg/i/WNZdRwUNO
l9U5CHk9rz5LqvloyDnnsfIXnuRIqocJD3tszUihxXy4oq+8E/l/dg0cd5ggHHrlLhKj9GxlrYAm
ooZ2KCp+OdvdiR+b6vjQQWv07Qh3mQkhKKR457/Vl0/pnzToQsvZS59Pnq1ui/v7AkCrADuUiHwc
Zmve7GtXig8RQpXY2o3EfS1lftEY2jDVtFkiX0X5XXldNmtx8jqy2IGoXZRfvcgdsXIdouOuRw6K
EvFhJx82xziacfJyli019PGsbd4JS9sMYN3KmzhZ3fLK5YdR3V1RGKVcE1vQJKaB7zZOvqL3XLYO
T54KZFLRnt+cLE2fg8sGHSmE+QLqL+lv5GvlXDhqxjqkZkO85cbMs2XOY8UyKyN0zG26LMhqdo6w
/SLhDUBdmNX5fAtRMI1w94D8W3eWUEAcv+wcnNlLgOW4M7nB+Hqhl3Wtos9Fwok/Wg/RHYhT7kr6
rxCshqx4ApBejxpnpGVSXpjecZiM3wV+dj453PhIUb4OykeHU2YiFLgYgPHD03xzOgZx1zjRHeKS
U/+EStuWeUAtAIFVmwupeRxeRX2e9AkCgTGPgHnUhx7QT1pw0+0y35BjMV4dnfPlvGgnumgX481a
+e4pCTo+jaLjlLn/x5hehmu8IyCPDm8BRYxtfj0vAMVPRFYBbiukUlSaT0erIyoskgbKrPuuxYuX
pk4Yezj08c5OdGhx9RrSezPM3tOprAUj+enBz1muNJDcEtQE1gznbcG34odObI3Cpi131T9GupxW
Bqb3nmx2sO+1a3tP6x46C6JV9iAex62Vp8lzsS0ZyyhejSRQaLOdNK7mbiOuaONOA4yUGAtuQ5Qr
5Uc2lmmLOWC4BWYVUTzuA0ELjYyC2v/u2HsPmTDOp//dsb72r4niGbl2Sii7x8MId9wvsCtjkz+7
WMb5mOPZDdXvTTC3PnzlkBONniWoVQW6I0yUJXUybayztAZsjEijTrHzLAayPNJy3RFSes2s2Bdm
ymveYZYZ5U7AWfxthILRvvS79sg3uXGYE+PC+d1L+aJj4wP5c2to+yTkfri36RpvkZB2ZJZQRrtg
ho+OD82Uy+dinl1Iy4mKofiOjdc3EdXlbQw6jRjVSvBk9oMdxvGYD8ooc8oYpFFUs6JfyU5+bQyp
B5y8nu+BmaCsTpzqlIbbxUsVO9dvloL9JE2WAjri1alhHWpN2odDEXI6PyrITLQsROPdvAWubvQv
9IKabvGWBofPOvADDK8FW+aZTHvK0bIGPhWZy7bkeGYw6gDnuyd33q4HeOx8Duro0MpDMc+up6zF
4sLGI2b1fCv5EagDZCOVdrUvfQAM30rVKsjvk5TBeseRsluY+Cys0y1L3uzxqhfS7rBMYdMeNOpg
8+Wbqg1su9Iw9sL5oXiZ9QamkrcEio3lHATTZQlJS1Bmq5WLQN+cu2md4xK2/EW3rqlcK+oCOki/
SfDk/8jCfZsLtQdURtbJeErQYqf5mFMBtwZnGqcNcgxwVtyBW9SIiRMgWOG1oF+0qk6T2g81ywdT
KSrvIB6bzbsVeFno4L6leqoSfyeIxnZo2DMvwuCipdBKplVLQrqs6YlurxcCJyQTomCFO5BhGjz+
YLL43INHUG/NXrJj/wThEuTLCQoomXc7zs+uBlQiXHjX9U6POKpARDN3ETDQmowA7MFp8zpM4lDp
cImh9NAmmDmY/1j2PjMWb4siqFlGDWI2TzhDQmZBvC+kFEBX4/yGmI5u7Sg0UPMaIWt/nXOMreEz
tUygXZGU06JXvqtgvtfgRMDgtVsCjXdxEyOb4CExUFBvZqYZxb4TEn6RUu5+A121GwXmE0VcRJiB
2kfYJCM91rhrLu5W2ycUwSlEYK7glVwuA1myxtn+kpg8QN+JZ8QD90eVqJgKX9Vjg6oJpbMmx1kU
djMORrcmKv/1/ptG3RiVTLNbke53VLE2xD+UmvQagPKm4wwjfOpY2oR3yh+tgKXrcceQ1MH8I2bP
9+Br3gms+TpPm7tzZPM0umt91vGQA1I9qmppH3AvlbaTx1MeciHp1JB65+A+gfn5VKL3tB5YR21P
cwG/V725mBWtrwcCDP2bcXvbm4mqLqzeJ/U3eumm1Oi+ODQpDYV8E+LVg9lQ8jd8BVmWbN5eAGVD
Wk6P5LRG4YUKOXw53Fy9BlG0YDaFL7b6rWtKmusiFEN1IhL98Q1L+w02OD3/Z4AGJQe5CuXKpkSS
bcvzzpQxfXetkFWVYInBrsgq4uTP3S7lV89gFU71zHRdbsG5nEVV4Aj1VBni/SADCa8OZX1A6t6W
/pXGXdlUQg/aCWBPwvsJLtJRMtl2ymIi+BZLp2tYjDHh4eETONbDIsGssqHqg45mBXjhoM4COyfC
Ztwr0ohK9CJvjcgvLT2svVPHINRIWaZ7G/kEs8b01EH5egHl9dtuHntQVFgEZljvAckV6W2wkoHn
nknZvem6E+zvcxVPF5HgprLwekCnYlgRKMDuBVtNCLvR251IZhhnbp8bPlDopvALBVweM3c84Mf1
fcSc9bEOYHUnMZwIG+xCxYf/jG0U54BAlIm0O16SlR3Yjgmh8RGALwA+apYs5eafEsnjkelAtr5D
Ifr0P+S44JvL1uUlEg8h0RwN6u5Me4+0oKY2/kLYzNYeK/IzFc+jMooHoyjiEh2OSbi03QPLGHxZ
Z0JtDVQjqF/dwQvCcQPnveIrG/2VYNYMPZXDotsGepfiK7i3hHkwGIHpt8Bmo2tavfI3y4Tit1lP
0aPGriPW7s4ZKSxURnLb/jiferim5PRYPkY/ACiGDC5536xjdeBhlAweAlF9mAJDU7XnCcXY1wvq
DFG9pDXyH30PIGlzptWRMliBDMriKfsRbj+T3WF5DK2Bp5dzoclkEqHk9d6BDvVgjwmOZ4xw89F0
BmvSHFRT3WYKhbqOTpwsqBHbG2LglvQFZFRsS9nCd33kzJAsJscFLvWBrEkguq8Vu9uIXH3hgpjl
b5/UgvWzC3cBGXjETMXMSoAjv4eKODST1I9SR6vxXYuh6bNlEtBRItVKCc07FJ+oJbYUmkTnLymG
iVwRklR5S0i3BJG1FGT+O+2S7XELQjNxeyy4cqbqYvP+wwBF+7mj5XZ6dTk4XcXDQP+cY6qpnyB0
TGqpTSxUHVPsGUw10bgDYm7RSBFr7Gkn50gooid0ojy0Xu7V0vUZLnyXXcBRmU6pNChws8eSqzJK
muhhKyyd37rsN5aWbVxHeIdyoTSiVplDe7sHR8f+40y0VYYx0RKAODmATGSdOfJa2+nK8muopb5V
e9clFoN8/YEg7J+2kpG4HpE0xWWcHS+5aSjBuztike6HKFBr9BIdgnqvkjAn1l1JM5Ww2onn3tf2
VcroKTQRsccIUvoAR41pwGRlu1QPc4kNxNj5LjslNbY6pup3GR8Vgb7VqXVlOhlLk/DVnUq7s+UC
1njisM8i2gfX90Z9Zcc9Hy3MIXxfFKjM0U51CsHr2l7L9WJms3cWRRv7zaE/JbOj8PRiLDq6Qpob
fgjxOPDtwDhs52BIA4TEFQjTJ78DqmlC7AhGgWEgqfHswef3lFP6LIf29ZF4jWWiOkEnoFKAcwGi
cwKVgk7bObWIGrEukE+lyR5z0LftHyPXj7gcC06+a7mqQ9yDWZIw26IAHNGDCCO3dPzp2U0/bwrS
IfHmtgj0suj1upHTMgSUXaMU6ob8qQOADeDTmAYx4ojYSCxjHeOFDWPBfMxnPKXHr7W3c5aVDvGE
gze5Be/ld6mlkhU44eQdkCT/fGJ78OVihA0y2wqKjFEzW3FI+pLr7pZWSPUlxl4GPvxvtP+EyKnt
jrdWdWEKSi5xu41uUhgN2GLpL3HYYneg7KF4yOqIREOFgH9lKcd31s9/u9Ed99F6uDkhSkcWOsxM
q+NIbbCg5QmxgpbfK78dsA2wDSosEZ6W7pQIBYFtYs1LmJkMZ8eF5yVIwNYvmSMN3+HQtgw8tmm0
SXhNOuk1wVSJ4klRZWD1GH1hdTyhpLDQ6pi4xjMITwvN18okv6VNdlMInRhPp/wp57tw4386qGqy
trMIGDqww+oBz/0DbzCf7wCmBBU6H8wP4f4lwwJ7vfq2p/OIZ1bsI2UoAZnbpUtCe8OI+4gZMDNy
xDWPNRuIzgk6iEt5yOySRQk4jh+4GaznL9EGBNeaJXLZhe021ct/rYGIh3wNAJW2lT1LAXVfUui9
DyxY7opFq5hrJ4PI3rgS4tkqHadFt3BPlF3nqeVGxgp+vE3zxu5oRzwYvqO9xMBKZlyAwpl5mEc/
Rd65FUdO8anqccvZbsawxOFlQD93t2Hkb5gwreWHoLkuSenZR79epZeRCeInN57UhN/pnv1XN989
FeTcyKYg8Q0kX8PW4LMMuhh7ePw6ea04HaqXfJ8C1O2RkPhHAMpTxU/yqG+MoEX+EiyfUz9OkmWB
Io0rBav6mh+rt67X2ivLBqzPcJ91XkwjNUb3o/pGVp+BxrDVR4t51DbcJ4ZKWOpyaaxT4NdOQU4q
9hrnkqmC8Vn8BfjzUYkIIfGnQRaZJGkawe0LnhIoHDcXg6liT+Lv/UkdpvMfpKF8PljY/uHJfxrs
W1+okUHWuw8fiN5BvxxkoYGcIc6WUsllsGi/NPsMFOuO1wYURXxuwyCdj+gEY6mTHIfK3s3iWqa3
MQT+lzXNHblff2YBGktJ89cefBsVNrsxyTxSWGtTG7WohuHD62upHfcsCGdVFsMWx3TTCZ5Spy5F
jrS2Zt7emuOizk13bxra/1dzXj8KsABhm1xdexrqDwqEi1DXnDkxxxCaHzmYQSenb5O4qFbZbHqe
W89WtJ0qfj5ZXrFeE0V9hjGPJCgS+ikbpMZkcAiHEp7rznQgGnU3hSOEFVF8ihvxEaIjYNfN59VZ
kx2JXokRZk5EZVRXHAH5K4iRRwz0ERfIsH9ti4TnGHVehnB07dkU55Wl5gIhTQGUfWczVFzCtJFy
0dUpZgO1U/GLQxUPEQQDKxKlYfOV4HCDD94m3pUTMvK5aANsGjmdlCEHTXIgAfr3ojj2DF6NIKSm
Bcd9bhSJzNgSUlgJ5Lno267Lyc4U2KCfkLXxCozivtIRWihZAayPPS8I2UcTCn0GgzYui3LEjIuG
zMK7inXM6GTwxca0mjec07RrKyi2rpey57ndD/pNp6YWVEUj2/6QfhcN3lebweDexyjQGn7eXpB0
fJwrf9u5ZNYTri5KUhn6yn9Wl1zl6Z/zaA07PlUM+oXcJnBQd7oxkHN4f/qnCPWg6wCBEsNdiYYb
Ywn9Rbv0cRpVrCeDfXCebUbIH6jWZ0izunw/eoWvDQu7sbut6bktKT95lAkazApZx5LN8EFZntOf
jG+LpKhZnZwlWswXV6MbQqKOh//Y0Q3uEH61n/EA3r+INJDHwDBt3ScMYX2VB2GvZyVmXBD0xIim
FvLG0qPwAbkQKWjw+qi/kXf2b3KLBWv7ZcfopFXJq0JUN6mEx1RB11k/r0QiTbc+Mau6d4xClFZI
9lEyh+pirTRXjdtjfbDG6JhL6tMSGCSMaNZJyuL/Wtto/Q8+a8i+az78Go/NVa/wzUKMI2NJ2Mno
DAABBMhztepcH3STkjKAy5/bIJQexJPRg8W6k+wKzevTu6+vQOwtWSPE2Qht1l8WElOO4d6/w+3U
z/fN5BbOq01l53cQAfo27WrVkOJq5XrEju7joqbf7F21bvVgr7ijmTORt35Ouh174FEtu8ziIbDY
C28m2y6qcACYJiyZ6t4E7fp8ywKGx7daNR2MXvZIIgsXegZnvmGvn5EdsWY3we+izvfokKzJ7K+3
U+jDQohU/zI/ApJ0oX3RbaTSyYUvFWSa2R+X8hjjNLq4s25NUoRzyxjgQo+L8QBaQ56dKkpLXpmr
TS0FjIxe+2hJIQQG8ZmIQ6H6KQPe8XIiWiC8yYSPIZnkksBgSMIMHKq9AwwgG+JwRD9pa/0NDPRV
3kP0G7ehebrXpo09YRd+5P0DVKAogTCfeH4rX9Z/gQHrEH7bI0okzbWhE2Bx2vUs5b/Q5MNC121L
oYTKMbbeKCaKDKiG0ZE7HnBGFMKyjUIZxlCggcrWTx2uZUVR0ELQ9IUli39AJA7j/F/oHKaKx/6E
HO7zZjTViOZcjB0KGPmTWtw3glho1KE1wIElw8ThhgGoLogBHfoda/33WXMuzozBkJJGINtTEqfp
Ecb0nWCCNWMHnLaRneomtxRtMinw0e0myL9xf5fBRzuLGYFpV9WHo4LduTs7/byfGxJkz7m8plkS
eLIesUM8tsJx+5kyuI4S9LcZ7UW2Huy2t4Vpm7lzRN9IhYsCc9XKqNtvnzbfuBnS5Gdv8p21jzZz
UuNJcfBETnng5QDSnYTmCA7CzX4OIbOhCYyNX5445SD1Pn7JmDe9JcjSdlMXU6jbsLE+BjVegjXJ
pkScvDs1bYcfuVWJbBQQwfktJossM4lUKtg3zRZxQNkfZwaKJKHqBNHiJqGUVkIYgjQWJb9OXLom
bAlAGmPelRvVjWUrgfyXeauxCKjQ8gxIfpMJQjik2h/biAAeu2UPV76I+GsITpu5v3QuJd5M4UtR
ShpQmT9o6G4/nKpq85vaFmYM2FFbrsC8PLyDgpN10mPot+mTcFQdepcsHS1LxMY0ouSbJK0CTIxN
jSI3pzf8j8OGNTT/TClmr8ZsyKyAgv3dxYcNvZd6NsKJsTCCj7f2I2SDEpQQXGjz9XME86JxcO6r
FUu3QKOhdMYDpjpuVHX0dGlKbTVSUf86DlkcrTBtuHhVFGMVWbfTpnXY59EwLpEyn8mXEkCzaQYr
8SElwDnUpk4EJ7IUUwYAY6qyQhRPVIlE5GA0nh/GxdD6kqgL0WfMhjgLsxGfw8teqJljflWgELIk
++iuK+6YgylHuYLAcvpB6csZ/tLeGL4fSTw0QhhCGf9Y5sYr3VihPpLt2xhlbjspKqcFKiqXbkHb
+PGBqVT9BUE3q0FrlzMgs1aV7bY+WYeO93G1ALjC6tfgFF84Cd+ldc9Kd4g4dEzFij9IivUDbYxM
jdAvK56nSbc0rLDCNLXh9DiwvwDlKtuKxPkCuru2HW4U04fCNT40XOxc+CRKPn5Fxl3zZLM+mbCt
ta7xXZH3I+kWtttF4OQJ7v/rDHIt29d5uLf44P6kjOM1uusVSR3eh2sknMDb8dhkjZjxgSwNEKr2
v/tCVTEC9VUCq6Hw0LoKvSa6Ws9FvA11QzLV8ePjzxa0+yOzIR4G9BwYU76KGdwqJ9nKHFEp5vR2
3WJy3STD7GoojN8SJvX9As7exEuUtzTPJj7Dge7Rjivl/bVsgTaFPhGxmG9odvFF7OQ1dpFxZy/Z
rzKlBuE9+w4QlFX2yBrw9zT03/wOVYtHFLwOZ10OvkE4RfR+MEaEsh2WS3aGb153b2WKHF4o3uv0
FDqbftn0VCI/1XHEr9IRbX1yhr11hsF+lQY5kf5AZDBb4W87ljOgA7Ofq1Ri9tL70VF2BiMrRdEt
2CTfgdVQX+93LMRs7Noj34rqbbmdAgiaiuHt8fmK8yCOFonunBUi+M0Y/eysFsWp9uTHBQ2ItLhI
39NKJEnC5bjMZZmDtFpzIgOpwKofpY66RMk82AouuQIVUy8os+O7P14YA9GIYoVW73OxM23N6kH+
zkKJvBOe8FI/ZQGVH1+IM3qwNyStbQfVeaq3Tfv/GavdDsicB+p3wQgIIpeifOdVla+L4QDPn2L+
9xz1Pqx3z0EAg26mtFbKkqe653+wL+eg54IsVVbCQcpO5bqbsUEOx32MEygm1EFg2/u2PnJl5o69
0w3D1qJXAHWUViK5ky3y4L1FEC75/W2Cg6JrNqq8XEnrLaUJVOl1X3GC0/kViastFNL5SP5whvhS
ubhhugb8xE58xzyPps1jSsknsyLHvdOgaqL2BRElj4bqePZ4cXjI5fGUHJPJARYdZiRLd/H0ihLi
2wjbREJGu9YusTu5oeqUYyDiNjBACSDesmYPfPl6I0cKn7lNQxmIWhhm9sGOIAU13gi6PISwU3Kv
6kcg/CIrOGPRxm7FYWKydxzQDY3GHy6/W/Hfj2gZcSqllrx3UvnomprzkH+p/R3G4sF6jMcIQDhu
QGBpTqp/4Pk9vaPT9mLbmVP8e43KsjTy7f1O4LTVxn8bikFHV/NBN3numtV7VZTMvzaoTu6zfY58
UAOKe3JsjO/q49AAtv3Zf4tHv1q0PZciXZrOH/Win3nd+LXMb/mxgiISlAieQEWCfKYwLAhmSnoD
j/9Z6q+ThVMa/y8ZXlMQRKhHqS7P1JoL9Nv1T02RQkNZ1PnKp6k571bVYZdkn30zuNWkL4cETbQi
EQJ3yy0j6Ysr5Dc87CwL0G6x4v8ZBXmQq7nkuo9Znilm7V7nhTZQhoKdMPH9zy+hu9PJr7ntllW6
zteHI3WxcLkEFg1fcOROUlgby4YohdYElpUFN2pk1zxOJwe2c3YsK1NDpU0wLtwH7tIYDtDyN17D
o3siBzOEnGWQP1AYOqLhffdabG3mLhIXIOdHxOyVrGwSx83aoQkvggdTkM3wndDnNT8OuqAZsML9
Eofymdk+BEndvr0hTm4VsubDeEKXVWCPryG45exC5g6F29knL7vJsL/TVH9paXGKpx8ai9MiDPkF
ssiZPpycCp6Vmg64bLiMvtZOaf6lk7QxzGhXtH/IAQRbiMz7x1q+S7mgYSS9DFVtftET08ZxB4xd
t/PeairqRm+2VcAS4AsXOgH3uE07p2UWxdRRVmYwDMLnVVPvwnIRL93uddCD/vpp5ZSeGSanl1gt
1YrZkAbSKIjkqGt3/RVQ4G4cOK/uefV+fwcNacf2G3Wxe2JlFKJbOVBTKrmCWb55i9uC3iWyKmMU
yVR5yITqSOt7lWSmhLjWb9EQEDr5D3BF5CGkQO5z/N1D1mV7dYs6SwPrs9QadSGMzoz3cn9nNQPa
30k/T5sPfbpZUwerjO8YJY6hnLhaUbP/CdGhdJ3iPPWLDihVm8TrMpDgT+EloGO36BHi/gHXdThZ
wimRWBMykuYfF6lZiBl/y3c5toglSSIXmfXG/nWLqv9G1LpbUIxjUjLSnEhReN9vufSYSMLlBlUN
m9mmxGFvyNvqi0YnynihwkQlJlQ3dGnCvbaK+dEFy+9m8p3u2C6CjIlStod/gEUmgkNLMcYRISYE
w7IT+FA+teOHhh3jHEAE1PZpLXu4+jC5Lbc7I7twPGrLyRb4xUkIfUjRwN3Aso8sVT3yTG+1M4Sz
jhUCj+qSRqB0eUtTBkBTj2c60LnLTSSwsIjuVM8ByqxIp6FOlpbRM9QJakIrMazzvScPBb9BJ8co
/1WYURBhjJ5tx9hfWHDLaG+RoQKHexHA/o2alvyKhqiT6De14eVRPFNPXxtkidyUcMR8ugJmkTtU
zGRvInpyFrWbRJrLN9S/odLqe6Owx3UG1RvKQ1QTJg0vDF2mX0IvUaolmtRzdW5PObYYL18zWNHP
ghtAOTJKajZaYrKofJ/qAW1J5ArY5LUwxZ5CU1Rlh2j7+iODe+EZtI60mMQAkYWMQ2IYnkxJBMMG
UNbngnkJtNR1g48pQMc7Id6YSdZxVVrKLHKf0B9kjYAKNNw+hlb2ZTkbJgyI/6BrF8tQQJmYB8os
Ojzgnrs7mQZ0z9mh1kOHiOVSxbtVG/Tuw3n6mN5xr1luY9B5vk4pq0OgLFCXWrTe3qRqcdnhZpnV
UwXJsV3v8txn1XC3dWx9EtuTBUqqOxJcukndV2MHEA1x+RrVOYkxcmJcqq8xG371p6EdFRsg48ku
CLlz0YJGyxJX5mDZsSiqreUjwuxYKgu/FgMeILZ5hH8D/Kfcj2iLVAuxTHcjwrB9Yt5EBxJrm+Vc
hkpWwp40+N2xC5A7UW2e2ntiGtYHPvwrxqh7uwOQHLvXm//SbHyRUK416VcHnmNgsKm9HkVsmTaK
Zvxv2D7dqgCRs5UD0XMwYbZerw8JwsroZLNZ8lRnz9Ip2iKJPfSy6tA1DzDPrjvKzv4RMINNLVFw
jq5NXcO083zRBXg/4pC0uIYHFMjGd9R0n35jCaZoVBFi9032jT19mncX9tSR5f/aCNceRT7z+vOR
nTMoF5b9yMx7nick34sI7FwjJSfuQRgveliMiiS9OezPUjSr2lE/+BltjDx2HoB+ZcJOGlI9Ly0G
QQaQ8pEszWeyiOPt/a23FFvBopI4nyAW90A6wAE7N+zwsOA6EHal9NoXYOjnkbdN1ywN6ptEig0i
M+/zAhaYC+GRHQI+EKct2mN3p9qWHRxT/jJHUxHzsESM3INPnArwINxlRclcGKsNpNdARVoppqTS
aznN7g934xUH3ALMwtz8RTyPj682u6+GZuXYbNEqxVjANr/WXEcvRZLIEHjDQ5SqBrFr8Sx9PmYV
4iZQ3GkDQm6R1mETFu23nDd5RWYnn4o8r7Sys8rxM4yqJkzFk1YD04iTKs2N2d/PiRDMvwLaa9DG
0hoPuiPcmiW5Vrv+7ioFNtMYgG2pHsG31hxxYY9wLWrsOh1bDBeL67yl3H3cYrH/OOFp4LO+JV+/
OPJyDAYbk+AyiDyWjYeHTnhCxlqKIIkgvJosnabFRKK7o45aBJQw0EwkvGp5erVuX7RIBenkMvaQ
8vyDyyO9hIufjDmdZ96x8Iy2JBuEvD9kh10FbkHYw6PM5clJzwBZRLO7BBXgwdAwHpx+Vm+AFO9g
+0fEeBHpcovOSyx/0iDuJYVDXBPCCVJQYSt8OkLAWIOpPchTHqOsJU9rY4Z4Z9Qj8iE1nyuNCad2
ggtJcg6m9ptU3Sej+7WNWqJKMbvklnYGurAiddWj0iMiGiwDes6LPLdnW0nCQgb42A//qgE+IV1D
Y/jaZUzco8CRdxGM0EaGXej0OoKmZIOVRJyEtXUDBhODcer4mkrF4Op+K4YAxHVab85pymlX0qqu
G/MXTzpnjxsbJQendZQyKCVpy+dMHRNXSBAMLqezuaZXgyqidYjqyr8qdvtEIlm81G0L0Fpgkzlm
c0VV9jE/5pFmaid+B+bVAYXhJbsgJ5YyB6FAy5Y8fVt/6GMMOu/89TyH6CS0xOGfh3Bi+a4oFce5
kpZAc1p2f2d+EQdr7H/Y2q4CUrx9ywHD+mzbl3XGuv3rc08TSHoAId3guhvyyVy1Krp833gobx4a
cLnLwEmIaYyc1aJ5GpLanyFRy4McySUV4dnYrS/hgYiJBaDF9DeeWKNSpEb1PSrdgBLGE+1iQ68W
BCA0b/vAHqTx7oaWceLSXaOd8tDr9kC2pIhukNBDoAafJ9Q5aUqXOotFMYHY5jGefeCGQ3Yx8BgT
otkIOtpIVqQFXg7Ub89HVhhwuO9q5t0M7Q2UApeQB/TsUq3dcoPRsWLIUOTdTALUs2YPrWlxMZzl
m1MJHly2TiDrPDAnXJMdRZRfg00ggXcilBuLEuivGlkYBlrUIve5nNEIf4lmdYQ7dyIzZfucRZO3
6MRBiQ3LmKlgPtXFWtPWxyugD9U4WnHlTw109qDGzuSnnvPQbgrciZudRJXocK8zzUOtuHKatBxy
5+e1k/prriursEk+nl9Yuj/CLwKIThKzaSf33fBXh9F8D20jLWKFO36OgIhiiUJJzPKIi+FVpj19
RC5F/KTEuCj0clzjo+vwU8rAdXjkBb50owFMH0DaaQm+ST0+6xYDLyrVIw8oJpS/M6d8Bew1q22J
u1I0dWDjjGO2isBwlHmzGp4IRgSAzdhyvemJrQwtaImdP2j+ifGX1A5/tMT06wOqZeZ+Pcvns2Sp
N90cRgETc99ovzgYc5ZOt4dD7sXrn+UxAh8FYRg82Ta8+d9kSYAKalclDZpoMK75uwGbm29Eyy6Z
N6P3UYVMb+vFSmJVQLndZImj44y/PE+MC/uEXbz4Th1oOsdNW/D5WcNtjsTSfiLWu/hGtLcmpBK/
eJ4d6avqESki4LrHFzL2mAm0nAmHkR0/2OAQX6f0YXtQHCg+oJPsrmcJlCXVK8bMf5M8i0QGL9ee
Ql6v1GWQ7SzuRHv4RzDjNHSYYTRRymSapQ3y49y0+GGtK5DGD0ksSWm0Nofv5U88F3z0IwgMu7IY
Opuuiw2LRnPVTpdwPnla/V30cEJh0Q4m4jb9tkHSyWuvOHQjHMoLJJugnN6luggtMwerfXesZZkr
uVOguZEk4Mv5NjSxph70VhXiT7cJYe5poNbHH7BSzQUtxRHwL+dw2+b4dfcBty4Alr9g9W20Anpn
P57Xh8xc5+kPhpt7gtNQldY/ewlkTUGdx5CYreDzGY27XP+0eTm/20haHo8pPvyQZeuuC/CwDgFn
ftq6n5vDj0o2IdVLfDgf8844ofKQYENC3b7yCePbo+tafnT6DWCcL021hRECBYmLfM4hI1AawlXS
/jNMcd2iTwAXzZ00eMLAH4hgBRlENc9eAkKv6WqICNM1VMNy8hhDJFSzEXy5M+/0tdPqE91Rz3A1
JKAAJgqV2SIFpvUNb5jd9JMNXCcDy2MS9rMtzGd6m+eULb8Q/uOK+cuI4BzTI/u0aD4YcaSBfXJy
eNe7o1o4zOVkmMWsyTbKzFFVabLw1qMjp0oukyFTmn0Sk0vv6cFr0hXY9khiLKfKu6XmCtsfZ7iz
r+IzLlCHzIIsLnDeNxHP2Jv3eHElV6YtZsd8a0ZVVsw3pZ8YEShthlRmTIBbesKId/YJItwLHkdx
sCFqs5CRx42MTPgZGRF4kiuwOUIEZF7/4PnJ+5Wfvd6oRbS/kX//Cbr4fbcKfaHk5Z1rhSgM+ucp
Hzm3hprOUvX3zXXlMy4xM5Kgr0hSSUl7KXAbyoSZyUTjNGPGWHuPLuqbWmOKJb9QUcR0NO4niMq7
tFi5iIaIssoSqXcKof/rGmGI6lCUfBS5xDitEtlZ0MAudKzrZYXZI/ooPgoFXyV6jQwJdm3Bkn+s
jcP7NVY50HQI7K152OuCxUOvdPkVi0Xd1r19fy085Io4Ji4IdkHOKtQELHiZzpojsWFeR8SLyof3
6pUo0YELJI+kGiaFldr/HlpAsnKxxFRfJfohq5v0SJwaEMFj0SrW/ar3K0eLt7oToiiaH4C06obL
YK8neLhyu1Eoi3yiTmloPJ/DdcfEskh6gppfYKssPUxz4+/3cI7fXIQqRKTgFL/T7kTbspl1ScMK
6WBmN4GC4Q18I4fE4QacgoI79O6POJeJlUWOTN7yjG5JX8DTib8CmPG9JI7z9X43zG9JUEzw6MtQ
zdi/vapUZaIP15tgeB2cR91aBzhZ0Cvvh8vVjVUOQiSAonvvu7mNCN/nZHaruZmDxpeuJ0kO3iPe
mG3fDs6z2pj7CY9voZftOBRClp5UBP1MjrM7NXXOv6VOvrC49/oJEl7N8O1d7I7RT37xc0yHKgga
c4d+Pd2WYPoII9K8Yrn/z2Ui4pZLz5+lcpgu3Xv4xKMtipL+b1ooNAS5oRR7BzSxj1KBp9U8+Wf8
8EMMFL3bQ9Ccj2irh8vIlnjshtgptPffO3pwlzrXCSS3n2OzaY3yxK9zIHn7NHYUfPH//9iDGEcQ
o5k+Pz3H9zFoSNeUyolDsMmQhBN9YzSPM5r9hb+20zVbo2bA48JNKUWHUj7B/jR4iKeBXbf2b5km
H1enfKSIFavCfQreyXTNQ328MFS0FfVaXGwn/1x8ktkv1AY8rPMLVfRmgZ2RJ2TO0eOYFnK84yDa
gwAVGL467lkyfu9N2uqMTZAf5W4lDG+VGFgJ6c03oYAi7RPhWMH1OdjHMPGQ831jkEJuL6mHE+KP
LtV+G3xrC44w6LUMzlpQZgpRykMhymMqcRQvA3yYwhtZ7GZDqcpITH86qGZJTyYR5skBr115QPBY
Nz5+nOW3uTLRhYGseDc4SIXKqp/7AVhY4K1IsNWkKdBIu/TM6nF31FqOjDN3lPpDQGxJhhGtt9LB
4qu8TzkKvINqDlz/vxUfWdE0pRu542FoKGA0p94uKvrN+5bowzZt4Xkq3TTUQzNp0WrhXCXlFJHm
2pOBNwCiMvZHd+/99SALrS9U3FGx27Si4gDQmBdWqhVY9FV9R8nxNUeHUES67ak46RG4jga/jP0H
uAtWcVTL+pXd4yklHFWs+i9/l3Rbu5BYYgyEFuKI/DEjaGAN72x38Fe7NI6bUvJkptIwhXQokWBc
uddQmP2uPnKuQ+fkXfP0/mgrawRuBB+4OTKhopE97mNUGZlVb5ixB5N4S8t0NfMO5pjFnvQXEIQn
XyU+6RL3FWSUgBZwFMtxWYwIQdznthoANjdUQWh3MhLOBXKR5mokcRxZK0P7y51QELRTYRTls0lu
6qlzKx7m7wlzMOpgy/pO8hWhQDlDuSdviTj0RdPads3B2e+SzOuyvqy7CPbVZU57PgF5qXf6nHQj
1YSGGjjJ7lZ9taEOloRFDHE9KOBg++QULnK/1zz4dQo0S0+9X89LwtBjvrB2JyyOSIKbNrxcYZ0/
7JW0V3P91+5Mnn/RdkU1h1fDnbpxpiIZFjo/O7UNxPmRJl9u+R2y6yXWH7ulrD2lpVaL44F/w7rS
trFGcVREXfx9nkYSz9xTZ+ooh3/QGbtFxxw4Y3zESt9zNNmz2YCggrXhMu2BCOcPlYW45mL7IVFL
ocgCKk+kFc52OrFCVmgFhEe86TqsgYOR5PDI1bOXKsRakXnMyeEsRbM30MrjUwZlcppOeNxSwz3S
HKqGWPJyxEik8Z9OxwRfSwdtrQWj7xwvyvK1cP5bC3OvMxVMNZyDWXEfEtettWZpWerSWjrRCcA9
5g3LE3t6MkBB/iQ7+xYGf99HVBNBaJp+MwZLxEYphrGq88LtHboj3hAFIJvS7XfmkYAMfW+G69Lx
soUzQPaOtWSn+JMhgG8QdMsysu98bbr9qO7lnGEkIlvtl7CZ8yqPKjZ0JPiOVvAryyBMZs44RpbT
F3glLki6aoIoZ8kfALNNH+LhkhY+lYPXdm+5SH22c5O7O/YyTv2vgX0hjkuXnAwMhukSSlc2G3RD
dqQck0UOU1V/1898l4K6b93uBKsSeGYwa4pSKFmzddrjKg7vCH4nU+9IBK0hX3FtBKrZbteI5fZi
zhdkRz9cb3NIAhITOargRf8kv1u3jRHjYtMpjZeV6eEh03aKw+7lFE0TamBsOivQvBcH5aN7fYaq
vixiv1+P3tJg3j/4CIJan9t0ezGmY+56B6DCJeZdL5utMMs1GMO31Vdp8xKNYs+8Y6F7J+hxPCxp
s5P3h5RpnhpQKwMgOuWlBfh79n2sDaXIEJrbAvobZSoaLdVC+ex2wbAc7okAhk2HUUCcRaHl0p21
cFIqO6lmUSJl7Zy0IoZ/kojakX9PXW8/B6PonJONvzexnC4QtwPlfmzqUrlK4m82JxzcaIRU5Wm3
/nR+0+MDTtrJhj+KWjksYD/3NQdVK2AOzY6DjeWWrzMtlY61jOLtquduMWVSnAzd8ujLRYHOAoST
yZ8cGLSWsq2VbomK/1qB3yaHV3qUp5zM6Z8mm9GmRjLyFXCgmct0oN9c1jVpRV8fGulLflM43m+I
078OjCeoJ3RZDFGOLbqcZ9ngQvrGdYVxpSEAn6S9WcPsFX3kt5a4WTNy2ISylC7ipFiM5QKY0FGE
ambjL2Pp6c8T2/sYB9fu2YqF6R66VKXChl2VPxGNdJjMRdDYs/6EQ032OS/P+iSk55/QXhR+BvY9
ngAeHGm2OBtTb68N/imSzBzx5dYNQqt2KRznRNGYHls5ffEn1PX0uujPgJZjMt+4qh+8NuM/b6iR
IB/da5OU6OFD/jsQtBOea9EYtrskl2L1Pimr3EtSKUGc73rNQOX1M/PAXpgBpQNf1aIVRLXq/5/k
X0sYGhcQuS5cAkkjtHQFu1p4zLlyKyHRg/t9bAzU5Ot6dUbUbMniJdd7EiWwChcM/QZqI0SbsBld
kKkDl4viVXXKX88h/0CjFpBrZK8LKRhYafg+Ls+m/amkMunL4OQmJzcHiHS1ok366SvbFBns02Va
MMT0R05qFLuePknrGwp+g4mGvEhKNIpvUtpvexUGOlElCeWVlT5pQOQAHxpIZ48BFGzFt7o9bg7M
RsUpDqf2cCUvPrUxezMvXf43dApghT/NzdxNT+utlEzTQi0n6PK3qbXcO8tEjPZbrAIQrn0pB+DN
NAwDG3NzlbpBPFmWRhqYgbJSqyMWS3NlQTWNM0r3o6EMkoazaom4Q01vE/El5Hd6ovjkPf2XqG6K
jvuXui2lheT4s/XBZeW9armjIL7RLLfSgJlXvEpDGHqLxLiKKLR/2et9+jtFI/2E+h4MN1iu/MWw
CZZJk1fXuDZaDxCU4ePx3+VeWDXui/WbbuDqiFHL6xWdjMUeWdrPrAkn8KtgEe+uKFca3qEai4Uj
mO/fm2xF+RI5BcQnZaRCLDreL9XUw1TTQ5pROBWAZuKgmwGGqP/rTZGw8tVHP7rmpJIDFOdyLWS3
iGH1BpDmG8KiaZH6mCClwRUxV64OSiiLuGzkzBCUMEaphMVd6k6e2FrK9uL/d9OSq5wFAu/BCUeJ
H3Ogs9rLcINQ9ISKT1esD9FuBISIQrS8KS3W5ZgH6q1CcSwBwlU+tGl6O3qNRN50KegY/+CLlLJk
wpVfd9LsH6Sovebp7glrxFuGCUanmhXniYtMHXj8pcX6FSWNrUH0PvQWGHNBpGdE2kUGc858S/Qp
IOiday2ZTtQgr3nBQShIyp/3lCRvfAy4nkwP4kLdm8lEEohEpUm/wvY6+5Bisk3S5pdhLDN7RXQf
Vz5IdXoa+xW5W6hiumpCx5T44zBn2JsE7MVwlZo+4n0IRWKJ5OhH9UemGTvv/5NX4TqxpfJVeSnQ
WCLThgTt+uOA2vs/NWgFqkcBjZxAI/guYkQWdL2vjPUJypdCcf10M6Hyv/F3mZqmu8oafCKoT6gi
/nROlsNlfm7JJ7i5nrX/TEH5kImt11w710RXsWgXBDFINABqiFr6Mr+k3iQmWIaPeab5sqUPUu/n
zksolgd15Py6Zl2Yn/mGHx8JQItm7pOVTLl2Ys7SDKNkZwF65swB6+1e7G80KmPs3MzluwJBR5hL
DA60oCWiSDwAyGgEr0BWd7v6Ts3VSPttpc7m3AgOhdV3NJ+9zokzd60tOM334gvXrKre82hVVZCj
ljZv2EEhnwoyDKOk/i9UCGzrEHShdeJtqD2VigGvyDrDqNvATg5iYx1qIsdoIumY1gfbykXfTB5Q
vAcus6OtLW49ux1UDWVthiDHb9p35A2wlHiIfj6QQqTuE95cuoueOELabKZs26kdG+pkOngLb4CK
Xdy1hWlJqxQ90sbiCulweZwGH5KAqWMfsmw4rHXB+0i06rpmLWz/w5REryv4UkugDY59ts4teBrI
y1Gey92yPfCkYamaS7hVIHBFQeW4BzPRVqusu/7YH0HxHVA+RcI8be3iW7jiaF9sZEEUz2bsuSac
hqsznDOj3EvHmoxtX5OjkTxxcb9zpLgRv1/joRHmpGbHZlUpgGjWXtXXJ7p2ftMfEhm2+AH9tMd2
NE2DHcefLyaNj9nBrY8ia3/NwzZmqI4cqJhxl2PYuSQ/w9I78Qvdx9XRfgVAWBJyHCfW8BOvEcq/
7xrr2i8pdIvDQ2yL0D45kNXmZ/7il1VSl/NaBgngYGERBjGDpzBV74D0xpNc7fQuQ8BE7Exv2bHJ
AOzx7Ww6Wvgd+DI5VzngiMw7HD8s/qquL442SdvuX+C6OcpW/nf3KEHVZbnBIUB/yzFKswbLJFd9
CDtjLpLatxD5jYj6ElWH8h32vLr0LSMYZ2aMzI3x049uL1BwwqT5QEmGD9yoky6IpWhVwkfzlvLe
4vfYfNeb4ApT9vdiQ7i4DFMsMHBqqTuRVGHeO2QOlItF1DxaQQB1TX8U8wnNW9Wk3BIoKuo2Jqy9
5/CGoqcqcBVU6piEP0gW8B31KDKjLAm6d/OhpBjKR+HqFT4HZ8bWFiYm/5UyDtfxd2bhI2lguVQI
ylr0kIlJik+xF2KP4kbLPUZ9PJjXhRw5AGkSZgBRM/v8NPljjBqS8uhfbZdhVSg9OQ7t3yAjTxhM
p+384H70OIHBUYqbwP1HP9bSNNVZoaXq56T52g6HEa2Wr/FUk9VvDwVtNs9H01drtQeBkLqBhgHR
HQ8HlDGn1UbHz4azLDePswl7siIppiVAAptLmrxE5T08qj76mMyhl0DW1VUSYhy5WiZopdFp1DIr
KW6i8cxvTsSsidXv04XNRbvEAuvTFqREerz3xCNhcVwg3i66xb/XOMT0ty9xAnl1jo1v9tbMo1h8
Uytt1DGPMhQwCQdplr0By4NPCgLXVD4jjTvrAbITRMHqCbjDsPKrUxO/Kvz7MWliYJ9v3GBr2jQL
R0tVCmtGedSQzXTNLrfjgMVkiRx42eXkD7o6wZS66+urPXkBkLx4OoQ6qtYPkULOjt2kZfe3djYV
2iUk6aQwTiZmam7mdKD7J0CUrQFod/6tfPmrT9ENeyFKPO8oucAF3x1MQD/oEC62vDpl15pUgG3R
AiYbkEleNLMUr2qfnBaNmE58o/jZk+4c+5q+bqNrSbp1OFGOx0R+AnEMYNdaqQBPAbLDjKSdRu0Z
32O6zBfGYLlw5bDtli42OyvA0jGFpyopmM31VmfdHu53NeKRupExatQUJUQs3cfwOkcVhseBnEZq
kJpFGehIiqltmH3eE7La3Ast9gBRdWr0sVqyRb69T0Coeo5n2O9n4Cx0wM8JSnal0nkC5hr4mG3G
PI/Q9MtYbvcfpQFFIaxYdZ4/XX3sp/szl4RONLysNEweXZWZebUIV6/iZOsgRFt7vOW9gRXbVhtP
kPy9TWZ/VFivZccR6RLrZbDe3j80HsD2/jpwl+QJMynUwoVaTi9MTajtwvRJbgEHcyngiNj9OZbl
BNffFDTVAZgac4IjpNx5qbw1967SIMkRdEicNIW4nI0lkuL0o5CM0RgFMME9z0NOHXwAAmbLYehj
qFsKmMBoQDYCo9PTS1pzfPkVNuIgPiSg2fSFYSrlZSo+1wkrZshJTMOjCQHCPVDWPVVXSKNSW+Ww
VJ3dMV6ZDqKid1oq0xryVTdd51BCEnwOHgI2IuhhllBpWdxTyQ5oL2+d042VF2J5NPvkzPowxyRC
j11HtfNwuBuOOKb5V3Z/Ex/ZL+3l0DonrM97jeLGq3+LUl4Z+pZYKVI89FmjAvBGDGbbfg4iSfEO
vZwbVan2R6kP0XPCpF7uCDqVmsiA+DFTcA2lROTpqgihx1LVbcFMxtYBv/puVfHqfKmO9zqYPOUL
qKmn9tuoecPEcpE2aGLy/DU7Jl55JWmH/dN3mR4sgxUN45dBRI0IMHavnmuIS3S/G2BzQ28dGgWf
g/cTs9RCUcp7ZPM2SDTTzHxMUnVt1wY/GQCdFq6aiF8wwGPh1U0YCDcWkcC7yl+pZXRgXg0uxOKv
20RlVw25GrO8W1fL2E+t6o0WCIoNb6cwgvbI+8Q7rGQ0ANdHTaFPW4gIKBxVfmy5zBV0hAqtCoD4
LFh5sDkspEQ2WEhOlJDHu+V1ougYNc02ULxs4mogdU6GG3yBV8vQslg65M33eLL2kmfoRUJIp996
4aspDao2xs/UMquAw2TpHm6rHzNIvP1x4uXHHlsfRVVaukEbuahOT6MSPqwKuBn6wIP8yH1Zni4N
5XOwzNY4mycaZ9Mx9SPJChhm8DaY6rai+ll1V8K5o3xv4XmJ9d85o0TmmfSSt4TOUVcRqE6eixVw
ry1D8RV1wxE2nZgUNkUqjBOQrzHublIJz1XARqjBxzb5Ff5V5+kDmiL+S787c+BQ6zpeCLqTinYI
C9LiyG9+Wqbl0vO7/MqpSHsQlqpo/o17lb6gVjClfAUQo1swbOQGLFoFkTSwSoirYKEQTkvDXx0j
1XbBhIzzewbElOdXuNOB4IOBeaUbsUDLWXZrmaB2sdQtHblpejGgXkd+zLQjtZ+xEfNYTnJCtEtU
LMiENTe49UyEcKcxIE426Vre1poeSU/RCmvQVZG3cqOrhqhLIQQYIy6t5MFF5Uh7EsMef4RSCM1Y
oJfdCTtz4VXmmNQESNiqgIIeSIs+pgpFFHFZ1lNqMj76kxOo/yLkmBuABWV9JpstGo9XfJbmTLzE
3kBVPwuvSSHXRlX08oh/d3SXlyH2INBRit+MXYfdTFHdLBYeYhWx8t6AbJwCQ5l0VzJKwI+bhMAv
p635JQzDuncSW+QXpWZkET05MExBC5pgbmzAah9fbB+lDAURnLQUgAqKi5VINgJFm6qNfwyEQsvQ
kmFfEVEooZ6yjIQP/92hzeKKMEAXQoycCSwb+PtemqSSY1rEO4Ye3Em6b1hZMJvrH4xgtYU4AlK3
7BY7gddZFR35wBxn9nQwRcZVo7FTmkTmFSNkI4ZKUXqefBbZxANxt6oCcn6xnenQJTNiR3P4DbCL
ihYb1qFi/bTmhwY12zDKvKvKCmxZHZRceYQaFVFhC5Ull1UKdo78REtrLpKmc2iDGGzbcCFS2QD1
dgi341L0CK3fRM0EKWkTqIFqAqyt+8hK2wrinukks4LDzKP4zssfG7whsPdRrXduB7XYIPjHeX8I
p/hb6M8XuFWE6Qmx34IM+9POt3RiKyc9Y4LMYlvHjeY9Uawiq1l7JU/ipawd/h49Ssz2nMt1ttNk
lKshATtDmvlisbwJPOKwyojuIEr+dyTtDOXPaNFtppiYuLnUbXumJAJLtOWnbaPSqz7Oq2/s2Hug
FtN6Vul52No2M6w1wJ/1q/aNifkjp1qGbaaSuH+mF+Zi+bwjesFvdZgkyHxr38TatcSLZk8Te5VO
ZC55SGwqUleac2hkD5kjWVBsm94+CZhkJX78XrmuUMJmX8B3/2xBX1OtVnIHtCpWj1VBp4xp2Qiw
MRXm5e18heWGUweWupx7W5Xe84oQfxFdDyuD6IT0Gz053O7N7fupYAQLbu7dDnTpcEUfKaNYHfro
XU8Z61KPZkI9MCRdxkBttrzid25LEzAoNWkjLFwoHo9Yb6qorE2vp/i4uvb/ukrLSGF3XrfpPQK8
6P9v26tN9Z+O9499ZDNdqgIAX4kFqK62eQKBrWngs5PPPJrIrIi9pK8WErDaUmEsEhtW8fos86oE
JoMrKe9JA2QaH25ztt92JkqIdxuTXoSyLM9sLT2bsz639KfE/Am3JzyJXaYdC4uYRoJStDMTA+6u
23drP3fpMkQXhfvpHOle4QRMwRNt2DYvzN2TpYZShTsQp/7mqWVzXFs8V5M5CX8zGGlLuM+qIgn7
rgPksi8nSvo+yssH30BzT8is34KQONFi0Rc08if9lTTMS04I1HIFFtjOxkYnU9ZRbONfkoBxirOK
4xMIRBhTKivVqi/SB5JIAUap/RoN2TCPh9Zni/9wZq8uwnVsFHyTq98DDanMWZeULWIAnuHwzDOj
AChcSyu6+EeVBJ1qONIlc2RfAsb6azYB1HSIdpgIDlhZMObn6ywOrOUt3sy+8+mUhgMqscIx6Rcs
OplnAB0cTkelhUpp9Qm1kiX+Fx9Ulv0yx3zUFzEcasd4zBfKzrrywFJeJ2lkLQFuT/3dc2M8+wR1
NJtXLVAuDPkSUlfRERh12VjGixtbEkjKMFtUwxFzaBZlBmePCFAn+GmCF3AD013RnQ4eW3LbTXnp
v0Yb3ZTQNiduvERufY/QzHrXmINCkahPZvWBqM7ZSooRUiHSG0KIAQ7ZBhVEOgzrqFkHI9m1zU4N
fiGSvdQsxTmYZ54d1yw8m90jTknX5LEMjugQzK95EX1LW4enF2OPQRzLxILTSG+Jt000DDoluBYz
hu/N/ml08z/Ht15LHC7yuu2d0KziypQBb1+lTWKw3bP2c3Qf4wxEJgMNsghqV4wB8nW7a6FOVI2K
q5+d4JrAXUHC2aVcchlfvKqcQINxaH2NDyXOToEpcj/fAHewbgl+W73fAQWI+uXly/qLYoBNuNY4
z1ExeUEO6qg8cafbKYVZugK9pNhrStbBdsdfuH4zDDW1QtOACbs6v0dlr01CToLWp2mjGA3p+Re3
5c/67oCLKDnrxmxCe+8p6/qoDSn/R6iYweqwDs4mmWTBAEVjHePp3nqhtB4ymaZ16GsYQ1OL54LL
3igIQpoptYYxEQEOxh45sXVVleNg7I4fotCnjrMu+b4xbJbfvHb6R2FHwIrfKY9bt8R5+dAobuRb
Tim+iEjhOCQ4pvmc0Dw+JweVb+z4WEfNHm17uYyfjg0ZXL5f1F/jNJfdLXkrRYEP9cr1otgdxYH2
xcmxFmvofDD3SXAeBtM6gmQeKtFXxC4WzRhEjLGxiQv9x5YPFj4k1T0W0elOQ5Y63OPeJ6Heq3F+
qAFKeunoxd3hT9bLSvclO9AZrDjOAJkP4MjQ4UqjIDgyQAcYqmvxBbSJM+dwKlp7Wn9J2C7zQsdJ
sZHrcMpfAO6c0i6elAQ2Sodmy94pymrlC79hFGsy9Vv2Mv3RgSAFE1OqI4CfCJfPx3/pdOPuKO6f
YXP5COfaQgBeTlEbgTqyhxnhETS7EMJfAExwrHVaGqwtImA6+af/dBZPkYM1GngnuY/UMDO6fiXf
52qS4XJ9VXbJ5LgFI2aEdYxUfNCfLCFJ9SDEwSWuEIufUZRqkg/4zq8oAOxX3zN5uDsLTscVriZQ
OqqosL62CHv5JJXe2DLZV1y8y49CLtutdfbuafwwJGRfDqqJCCnwr5RDzClO+FIhVXRwfMKi5xJu
yqwrGJgw0SJO+/F5qOTgvyE4Z8gSrP2GjJvts6lSQ8GfE7y/glMimm2r4yQwUgihTAN7WJ6tXYYO
7cD/OwZYLkdBNnKw6MWEsJwQ/Iu8tS2hsAjJI0J/kFyuMecoFJd7FjP1iBnudDkB1Bwgz0LcXSlX
h7vRcAdYzKBEAG1Id2cjCKpzFWmUguTu/L/lsO9qEOQJR2zr9kGmVcmR37E2Ha1KszOjeL+poS2M
7WJEldcIk9ibruoEZpBLK93IK+y6KJglzUEeoPP/HwAWZtmlaDMDqhqmMJYKUIVcDFxd81MFUAHB
lXXGU8kOQnJcCvRFQbLUH2XVxRRFULRhWbBT0ZH7tJu3Oqvghcyi2LHRdCBZSj98s7onyKVE6IM0
SXnaqXM6zvOCL7QT+0qB9Z6CmGIdyvjRNHEmg2rXKPOHZ+2buOIP0ue2oPfcT2wohLYOWQ0znC91
EzIwFGhXGgGfnAj25xuZAQJPKdK8GhP4dXbdjhmr9SdNiVKobhyNykHWZsJ8XkYFOt7bSWCJKvNR
s/+fawV3PNFdY9LXQXBx5D6Yi0WaXQoNzm5rWoK6iRI/kL1i8/lj7J7Y1fs31hdjfAB+a/sZhkem
4Ote7CNvwDQc+69wjXtgyIYyzBHDuv/ripTg3W8QJmq6dIfvsU66XNNkskL3QnZEYLuHGFB+BrXt
r5RyTk+T9H9435ir4BdguI6V80KQqDIPnjUoAcyL8Oc03I1qE9SSAOzHvs16GQljsMa6qQEVCbF9
RK+Sbu8sq4UtkYR4b+F3Yx5DK53+6A7yyJkrQYo8vHzJ6LDcg3xtx7cFApce1rjWSosx8j5kWL5w
KtQO5lPJWNUwgDoPJZg4Q7+OBS5GM0PGCSqokWIS8dW6HwJhA8KY2T8TGCOJuDpFOqQOlavmjwRC
Q//sx14TNtDVEHDzpYEcyfKp/dfvX10qUDX0NLDs4Rxnd5w/39kPU0+nUwGDup9/iwdZTKaV+F3W
5wRww9FpZzW6nCD0gw7XtWWomhSSorILyIZMTE03cDKogkjmW9fkvYN+QIE24BWY1II4ovtgc7HD
6Tz465UR2sFaWs2lcCXld8uO4AYJZAJHNY8GAUFSULxWhuqr6jgoUNswIHrQUy3Mx4FAWqH0ikA4
JAqri/IidExfNmLxPUw23jULAgi7l3dwDFAM70tvJtYs+2Ti7Izz/wzmrkdR+OXZseRpaU8zdE17
R7Q5qysrLR/tzFSdaXt2Hmka5rP0KavruV/0XER9DEKa9UI3gXmmJI89f5i6Eu8fm1ex4JFd8602
bauMY/kkG6NckXkTyP+F8VUAYIelFmtFil8VhFfoBSYsoB6OuaJge2PxoSvJErkRxJfKJI9MmNql
8a9acvE1tQrdaMlekFcUkEgaRuwroOJjWzDPyCV2iBoW40qlP6So+w4TPQSbQde934XumYM2Ry5U
g7iq+757rAOz41WcXk06N9VLw7gs0vZJ21/1XOSAGanHr98DIdbfr/YWii+W0ZmEpJAxjsDbTS16
q2nZ6iTCEsy/vyjBwi9NBRO7dC6E0zwt6HZ+zdmYtpoq3owAdrPio03x1Oa06XLatfb4y43nN3uU
2PNx+XqvcBDiG5KIx5XO9ConFl05C5hfC26faSrdt8ayN63DFYBu2RzpFlVYMvRvHpfbU4ijIkNZ
Cx1VVCY+YHaDPKAX3iixKyKQ4YjLpwQhTjcJmShr34ldPiqLA0T8c1S9a4nojM+yYDa7SexlvQL5
Er/UzIywHtxy8ba2tOCYIKLk0An++cBvlBuCNBPh+2D/St6zcakccuS/BXzFvqPrRstOcLgklAxd
LEwsRe6bYqvSOPwa2758Sh4PVlFTUPFku1TaL3/T51PCaeSbDIMiloBHv2HI8ajQLLvaWS5Xz+At
F7+hIrkSbL5QZIKG1sT4FusGfojuTJjKkDAYhhkvQ6E12cja/gY5UlArAc1vMXLryVxxj7GY+cci
CwncWtC172dpf6akZIMZ/dNiv3k/ex6EhcykzGIqEKl2YRcNaoh+u/+8I9gxpXbLYLvwliQUV0sl
DKgM63s5XbYUK0OJK+braN1rXRTAZZ7xfZIsof04zTvuqpuExAs7+DSOQ2DABwOkVUyQ0wV0Awsa
GrjZRuCOU/jQKDhQtno3LHVltB/nhvPajYq6KhnWSsu5q3p2Rg6ib6mq+/o5d1FAhw65FpswLvT9
G3898zUuso8sSQS2/q3ITb/E7XuZ/2ZeoMTEbeLE5dzCjgMY602RPNm/BwRSApPvqTXKYf161sZK
D0q43fgEUFjsFk7I4O8JJiuYaorPxXo2Wczuq5M6j8jGKakk4YmXQF3WcPi3aJL9oqb3K9l84mkY
gcrvKljIN3s0m63s7ksA7cQQkxOsZAvXeUBwCeEf6XOYRbpxIg0TFhOkU1yAo1INXM3qJwi11Bgj
VUVoQSQQLMzj2G6NVI8hlbSHEDclnK92p1mKIjUAZOrYV4l+JwDuDSudI4DWvZNZNEEdVoanvu+T
Fd4ffBMFGDSZ8Xt/iLfF3Md/nHb3iPVnPMTh7jhnSWsFKa1PZBDu96UjVx11PjqUaUPiFHBu8PTC
pBxFp1F9BivrVjYhrizC+Gqk92H9QfYOrB9r3XrGuNUmeTdRiLY5SBlI9llssyHWp04DPH+3XpWN
W4Du0uANviLI3CZjdMLIWs1HnA3vtcQat7TE0ot1zUMZIeNus8rzO/+7bU9MenrkjHsK1BAJn8ri
9AwDuUNJtIZ2+CBV2mjgVLtsOm+Hu2lmpFhZpC4H2O+2A17aQWZq3n4r5ki1urlx4N1ug2f1WML2
eRp2qeQaG2zhDccCADGDaD8HTpRHvuvREd0aWyQ0HEC10kiiXGIFryyg1tqKb+Il8rpT1GiB4pSb
g0UqtK9sxGvGsrz465K3YZCh6xPz9iWz5J62KSLjYvtDAFA+/QbTW9nUGxPD+UimOXKLWhyAp4VB
eGJ08QHmOCiIcLzAlkG/bL2Ow780rnABzBdaQuzt1d+cAKovdQp9RMxo9BNVOy4YBtCKXn6EpqLJ
Ua98/VcafiBkUBsSOIcSZ93UhCJgOgQmjU6k/aKRMa3QR0JtF7jNBKsnpyGn82xkOVAWOS7tY2oR
8ou9j+bspGC2qxPL7uDMqfAYLsS/tenSZTOGky52FbDwrbh3aDgg9g2UUwqj9jG4Aedvew77EtVr
RluyVu7HCUCyE4SfDBDVPdayxTuLfvQUeSN8kWNwBmQ6mV38NegDgn+X3NCqD5Fps28hQSfsPfIz
lj6l1GHHm+nt0xU2neQRNOSxlojDkEw0z6u3Qpk276Xz1qORjxVkHFW8olSXYntKEU8exvcfW6Pc
xDWCrVDW4fTRdlGHCn2GtMBywolTThPZGM5yJ1xJTHy4TAyMrSpMMx7xzmXHifBhurVLU5XzwyF3
tCYGtReYj7thqhW/lNat5rwNSQgQcjU35UHgSvJsli4oSV0cLDqz7vaNaOCNiUKfzOawIhdhtX2h
nX0eoYoyegJ95BHybfVPq5U/QdEy4K38t1po2MTcT4WzEyx3y+i0+irl9M+ldb+oUsGIlDuZg/Mg
zpOplmrYm9s9mu1+4Um5I9Wc/7HmSXb3J+goNE3TpMxp7piFm/Eq1u6f4ClVSxGwhEli5bV6GGjT
PiM4mVV5LD4QqnqQF1tMfClR1dolKpeFRjOzQmKQL+uRtXCAOonpL2qLkRLgqy1zpivtsa7nBezt
iT/NVUK6KLPBzxtp9HaXr6zhN0hnXecTq+mScFGAMxLssP7lGli7+eSyhShDBjVJXdjdktevNVO8
z/ACOu0y2lZrn6pxCkvgzMnqlI6dwM/BPWXPjVbjudHimguReA/vLzcUkL22B+uJFwfhIJr/EI9L
jc0y9L/YA1fay0jkMp9nPrRqmmTr7eg0janSkPAqo4bgAjefEGBzMa1ki/r2MN0hf7APEAXCefZO
g/3Zk1chKvKa4AjSAoeBABbODJccrUomq2N8IY59la+nrBQwlCTvl0sokK98RzY4VM+ux/7fIQMa
Bsj3xzyfHZZHeW+64pzdYNDU/onGRJy9fuOWMCYTcjod1rodry37hYoXXygmYq5ihyez01xYyVTf
1kjuXJwMV0RXRlDx2MDZSviB8uFBEDy0tlWviwW4CxUzKegzBBZ2r1Sms8tKcYnrP8hceXY1+hO6
P+KOeacMC5gE3+7WTqk9pNG0VWOlOdW8KmRDbT363Pr7UlHZu2qLQSzmwD8PjuHgiRL6e28Pnx7c
K2BLqubs1mVaHFnDecebgexynMyNhZ04YXpneLfgMGrWQWfK0qQemhfNwa77/nhi0xr3bpUorkxz
ltwln+WEluTOAxSkYoELQzmSfuct6HjIZP7Gp3YgfjhDCjuD71CD1+p351tJvqVV2oMfQBKxDf/C
/u2d6U77aFrS8LLzFSERI0CJFe8zDuin0kJ50Sf1Tl+LojI+PEtlZoCNnHrZIlbE3P7Jj4la7SD2
6pPAQ0YNKNSEIhFXwTBnGVSfqtP0QgIQu/67p2kmnEgNmVOKvDqYmd/xCHs5K7LCw9PW3ZKYYInt
hSWQrJgJduFBoPGmTandwmeYUWzVnUsmfMZOp4pwg+pauQSzD0M4DZS+B0RrhPlWBYGahQU5V+HE
XoGTnLpeQvzJN/GBT9/+iWqhkG6NYnO9EFm3N7MUTNlHAj/Hi1paaDJdJYwcbAw2sWbuXdjIczXw
y3iBZNAfSu/ru1m3L4yyFIJPHhlzD3aOIoT7qg+Z6kjfGlzFB2yD2SpuQjW1YMMFOFSOcIR359Tg
IKuKXq3k9gO14PDeYglC2Md09B0Rk2oFzkuPpagoXYVeZOMk0ww/xnv0WLSw6pc0iKLtaq/C3Lul
l3D5dKwhBrnNhXjOBONRsoYVT73acnni/OYrqCnKVLlytTyJ8JeTiphWLz74KXPCIK4Sy01Xrl/E
fug0P5IF0ZgxA8WiFypJ5AZFXUvMzxS7ngPGyP0D5szElfafRFKQOYCmoLCQHFnJ24cGO4gylq5U
e5U2HQXPDRRu6Jscx5sD5PU+Oax4pIGGekFH9QsPWKO2NVesa8pTkuh6M7MtZDFqo+f54209r/19
05XOzFMp7Kpwa0HfTfkxg//9z5xw8hABEpX0Nn9LoQ7ZS72OmufprM8M5HRJT4s2mvy4LsPKSGwq
qhSYx2KHIq+agARRyPJ0QilcyjP40Mxkxxbnx/kKRVmWci0LVqTMyAr82n4UPQTrLz88wndTnRtz
gs9aNMTeCaHaiWC9fnSXKbtNs9FjZgGFzeQhLIOCMJ6lMkCDeB44YQUTnxxMeazV2JnzP/heb/x2
wt29/gUHEAGtqpZYk7Z1W+wZgfkYIMLTkB3dLh/k4+Dt3rio7+6L8Vf5oaomiqivR09jwGUXa+Q/
cXbFwOy2D4ajMX3/XmFDGv8Fvu4DjbRbUhhaZe4A8OUO6PZVaKqJW1PEjz8qgDTtcUTizf+OFDwa
nC8ZBFl1npirKv954nj4X5kkzFGtv1ZDxAkN3XpkI2FEezlbR/u3Ra/kCFQEOcsyrHISuh9boAt2
l0OfLE33d0kfpShij0oAvIUgMQZWcoo0MTsF041lWR/2BoOrlmsMUIs4s2NeICLG9w62/SdqxjY+
bPpHKIGSPIGFgZ2nUgLpVFifmFbKag25hRGTlcVG1dqmQIx9Gf9xy43P45I8Pe6HwGQgnLmkc8qU
g7KT94EjdapK3+0DKYEyB7UavytSgGrYnvwfLAIAqcOAgW2qpTylMvM8jJRWM94guNoGbSivu/83
j8CBEfqC7dNGJIVVyK2zFS5aqZY+IM1RNMxptQgD4Y/xODEW+wBGeqMYhKCz1KxWTVTSVAkFwvoj
Ov49CRuqb32l/iDl1BH1cqIdUisrcsJBIydzDCd0cgtEmTDu1pM5wMHbacHOR2vBE4p+kColP9sB
U2HLu4BGTl+1CKm9FVzMbITpg7cb3yubUmIvbREat4KpeXI7o6lLOd7+jMjEqnjtN72IiJQcXdeR
UB5cb7x2ZtIkoo3yBuGzD/PMoDpXkUL1MtBtxGpqTe59rGeGZW4RAEqSnP82NLTpGk5B9vm2rqQY
g2tE3KMVt/wdRculqLWNugFi5dk4Hj465ho4yEjfj8XV6S+zj6lEjJQSJ8j3ST4aVRC/T5hHfBqf
TBD0BPzlqJ9/SDz4pQDf80k+93of4O9PPKNzIjR/7sfrMA/8G5UZh4TpcB2OeZ6PXA4mZX2LZOI3
zEeda0zpp4al0u7zO+WBmuMMZKjZIgtIPxhBD/kmyMqTKrrNeRF1IWqStLtJTG5bldbW9UGFd9XY
heIa4VvPkDLqPvgq6rB3zvFYrI88QjYwktLLQzb7TlnSSagMYabKkArQwXXRXfcSg+T1ClxX7mOy
mhoRA/iwF863Ww1a3jziG/h3LzSyWtczd/hy+u6KpSOyVouPs9IOMepzy+czJGm96ikI4Dz9cscA
4Y0ewX81MK5Qd+t9CUqmddA506rIej7q6w7tG58sBl3OEsv/6Yt+D77gukU29GygfN89v/4GJG1G
qNLO6gjMrlCrEhRZ72Bu7nYpdpY8OUXmx9H3d43Js3MmJKsVgPQzNG28jasRTG6ILylpLIZc6vBi
6DlPC10UiSsDvCTQOzKua/kZEedVBiHVKoeCxQe8Mz+uoxG0wQ87e/VbjiZ7L5qB+0WOVkoqr5j0
sY/egsB+n0bO2clGXXfGPXH1nu87yk05w32palgobfiP5yTLAh5jynD2giha8tI8LtjbvbDPapwb
7zd9HvuH9BMwnQ3EyRIA/TLbKLQ4rnsI8MC3ZadhG0d6D+s2t7aLHZqlvJF4cfl3VFp9oGfjQeDt
QAj17aLsdjg3h1BSZq5rE/w3rMfqYE+VwyZd3F5RHfsmFMnI0s318qTQQyxwrO5o2lWoXiIV3yj3
EZ7GJwMFldzH19xmPcahjb4pJrfwubSLwVT4SQsQxdgXIykZnGQMq2LiKyu9sL7W66itiCwgcGeS
kDK2J1af2n8mYC053mPj4UdCqutEPYcPlB2ttwefSRxwjJmW32jKX1l3Z269DaJAp2nLSbqm9RaI
gAlEWVE7YeCc7XKB8yME38UQMfn+TgtLFn4pxr9e2vwf2NV+YHgq0Muxa5onkvnLLvRslFhV+YLq
Fq61nRn3b2nU7Kv6miPtPKyseRpqFe71HawIhRSk5rL22O+acA67Zg3fd/avSSu4N+iCwQpBPcrP
927425vdrHY5497V4IbVO5ECIQiFY7/9NHz1uu4J+p6hApSIrWDWg9W4YcUujK797VQfSQSQlbDX
6o/THdrwrPxox1uyxp4s6frvJ45qCwaMtQGBx1Vb3E3eavd2sj9FyyUcOdHxmILJ1VJrJyxX7QNi
fOl18vHTJF9/ffU0m+t6iW7IhjAM4/aFyhQQqeVTFrbmjzSGHgBZKksqwRQ2yE6HuAv3uIObGJO7
MsaFw5aWE4A28/asedr6YMr4jjXq5oTPp6lj4i2RgwSCnZYTnkPqv+UN4TXkct+g9100jXTXblSD
IYvargU+a6YqbwnZ1CBAqTAIeKrD6ErMlCuH1SVwe4tGg4Y/bOZ9khurH+r1/CWGinoFDXyVx2Z9
s9D6q7rqQMWYi3IYOzZGRVP+okak1ej9ZEZPAiuzJQdwtQB7a8MGbBQ1WDtwVPgNrfjxlpo+w/6M
CGi4phsxnJsLTVfGyKv80Q6/BENTRgLuHDYeR0oa4Rk8YuViJ23UU2xu2LGf0NXvxbVrylubOOxA
LHqIMRaeCaNTv4JJ9b7l/DOmq5gbJVpzVziuvNmThv321ppixRH/8bqGrR47n4E1eKIkJLTcet9l
+f46WMT8m/zIxe1JQafeetqtK4dDYC2U7z/5PbHHG8HlvYQMx9MPONLBE6ICxI/sDEDVdr8cgQvQ
98QQ1KoIBm5OdgI/6IAqUhJYGrWt/wKHdGca4P3lWNKUFzDhqk0/WzgYmv8y2cM/MvA1M8RlGhCp
/Qk1wX+zqY++uvHZrh9ehewRJ/FTAKhxtOIyj4MkAd6UlvabWepbzFDOzMDFTAW1wynmbInzEHXr
puEykoVGqm4HhRxi1PxVU4YXEg/jvlVlaLL/odt5JTNmIkbcHucaCm24LRBdRtPzRr/Zkyj1KiuT
rf3lZToOEAaAnAPxUSPiUYEPm+3J6wyePi6VtTo0S6dh4gE6gO+1LHbZMelfsd7xdifXVrExSS54
8X+hsV2QXOjAjVNI4Pu6lXmurSjdyDYfF19KpP6CgjlHnnOigtQO3+7R9FMsxVSK3ATmPwvAOAq2
dTUGnXpuWmVHPBhOGPckYEwJdFbib9z0BmI05Pa8plNMFepTKn63aOg2clB+MSMI8rt+ZoDLLCrW
dNcc4Qws3yaywP16ns29yjOFSbY2/r3VFOxLbpPyGTF+oNRhI6u90sQdtk/8HTPoFPL/cUt9sfXa
91pdkstL35kKVJutNX+XiZhfdkFJytrc8WIzjPAgqYtzS/CxOrij/RQcy2+P8Ub9TtnAodJ8z7Pa
eIGs5qEhznBP5EpGVl4lAkixEvALd8EGMq1+QC/oH/rRqLM0ZBLsXpoP+26jiiHlXWfeg3Vrsyq0
0gbpNpYIFgpdJvlO7stW+eI7gmin/s3ZBImoz+N24edQQzEazpgx1qyhJ+96l3TZfl+2/5iIE6nI
fzGyqoBuRqQTOiIuM9nvcO8cgGH3uhAbRmsvc/wV8Cn0DNDTJ8tfr7R/q61oQzwN/+0Z+nMP6OcA
AoeKxUI230wkaM3s4awDzEB3kVyf3pdxjCEh/EwC5yUcS3lCAMn4FLrigE4+G1aprhS1Re2CA+fw
XeGn9jM/JI20GJLjHj3ZFZ8t/6Ac2mRdywc6e0xQuEYQRv7gbloRzRz+8qhK02Iv/8RYhqrC5siV
hN/B3I5i9ojBPHfTqgQW2v97OsLRT+eol8v8wIuuo1s18a8siekaQgNqMJKFXgIoW2+9wT9BJHp/
S27lCIuyU3PQ719G8ujfe3lRimTdu6xYh7PMH91fAutMfoCB6JpOFiNkuxifIeEnC3ipxCAckO3g
ep3pP4adSbhsWlR6fBFsdsuJXKkjyIP1wlqMba3QeLqNrxPYQidXmf1/C6PPLw6/MF4xz997hxYk
7XeYKomm6WzB9YoMnNuunzw0k7PrPQ334Z4XVSPWMR8Ony5DkjYlLjDhRLzApzVnWdO7lrK2fOY/
cu0zyici4HDJbFkwrBXD/G9a9Y5TTgEb+N071joxWuiKofLzSMmCcxfNPMDbFFHxjSFsh4K9Hl4V
tcK/uTkmk/S8ikFB8M2uEqaaSdg1NUaRWLxZmbQZOe1okXOHRklkhY8CKannlWQp60LCUwC1aMtV
l2yOu+b6znY95Wjou9gDIgiPxU8UU/2i+K03Aj/ovUR0cSlDLRB2Rz8XKwuAzQvzNZKSKIlae6un
FdmNz2fptbvfiJN9Wxlbw/0mtwVlYTzUjcUoTthB2VSqTHF804gti+yN27T6Il4VIvcTtXzrhAHH
dgSDfKzAP1RX8oH0W2jhUQYj/tvhtSXegXxK0p6jJXE6WF9SPCHD9PXAlHwDvkJnOI7HZgRDq9kJ
ZnJ6iDJ5SHEshVd6aXICPZ5UPegVOWZRGBw6KNAtHVhB84JSLMURIjbMWLRUT/8zjhy5Nv3KB1T1
eBZVtG4NUC608W56v3bL8Vbspeo8RWTWYoOLR3DY4k6ZboG3SHBo7gNN0bIVnP8asQXjqCveJQJo
886Yai+X29mWZ7kXN897lARKK0BDW2szQPA3UcTH3qefG5PBqKa7HY5u3nJCfr50w/T+leo4lmle
DjYaTLa4hfXSamvYj1kSpskvg5nD54UzWO51Q/wLYnVkf85CcPCn2f43rQT/i86a4d9dtTfCa+I6
Wqk6rZw64Cb0sclWb8U+jEbkSNAoUiwdNsBb3jaDic+VmfmP2srwI1AQjOilzSH9GJezuFLh30yE
XZ5+no/Hw7yBlpeZ6I6EwTP44o9k9IJs+Ra8++2x3GNaRMEMBYCy5oa7m3uxkGhjjHNNwE26jdgR
FYZdmVMlknSbg966WuetTkx3O7ZJZwQFqgYS0R5a2egvTs3eHeMAyHLkJxsBr77Z2xpkKvzRQoXa
ABBSMHMA+1lxapPJA4bbDC/4IBk4BMOCKNwzoSLhPF92qxlSfI2sb83Oo5Mq4pbz5fxplfevSOO/
L6OG3r6x2mhcDEg//x96o7eZ1X7Q26K7FJsPfa1vYthq8NkrARXgDkTWmdF1xVDbHhaXxCDV0Yzk
5sfWbDZd7XwgsHUKR+aEazaCD33KWpvXDj1SwOZy8jstXoUqVETk8IZpOU7ur/kd3Uz2kg0f34O3
PDIBgPyKWOhTxLBzRtWAcOnsTVjfz6Vt2dOP25UnskRAmNfrPxU+5YXhZs3ZkNZRFDcr+VJRn+E2
p9odz8hqsSBqcFbNDahnUMcg3cPIWo12ZELfDCtsjudusC3aw51CtSVrJR0vNxAtrD3OivGTABV7
I+P1dPLbkcGY+hZjoISaHTxXOD2FqM1vRGPEiZ3axlhDwmOLuARJzT13ABUa/Wb3vHx3QrXxXA8V
jZ3FCXJFoQ694lmxQPKluAm901TDyD6ShIWPgYcSp1CHvqgBuqP61BkHlTAELCGyJpxnTCpAv5UO
YebqYFuBUJIgsTdASyfij2kYw4RJJuDhOP+phxu+H1D5WhNx8T1nMRskOB89CHzxsN3fpS251gXe
OkF9gM+QPsQgrWAnMraGYoHnrJ7EWSIOmvZOXvy4Q3P1GJLXA5FPr/9H0BJwOguqDX9SjPIF2fb5
FbyPolQC7jH1GWMkvC1aVRRkTnRAcHaWVFUTsKlYm3xaaaRzn0fSeVTX0t2T7E6kggsO6UeGAKO/
8I3+34gHhPB7SWgc6DwzPtTd4DSub7umoVdzMCY6WmQaDMqRmbiFsJaovSz9xx5+snDepcZQXaj8
xa71l6umpSnjfR6E1zVXMvvJDpKLwGVd02hyLlp5/D3rOfFwT3QD0+MH/yTLxvG/6UWcbqlHzgWn
xzqR6EylDXY//UuihKBBb3egBAnZz6ISX/A3lrYZ0xoSBo4IhPPRWgfpv/dAI9bS2Ga2u11IfVnt
vCZ8Xr+IsV1JR4ZgPEE3201ZbDbY1KQV2V06YqaWhx0rfiq8VrGakk/6+xLuuUo2KRrYmEn1yBsE
FHNydxHUST5ZKPqExyfR6nW/yN4jgj3Ht3FdqWfNzXVJUjDifPa/Vc0eD/EgVRdjDlHi8gUuEX33
EZr5dDPliA7TpzEN5/+zx77XjYGJJCfvxah1XLS111i3ygfC5+wWyEnhvX9Gupwql2I6fEwkydlp
sijElYllW2tgInuxsZJTj0QXV5ifovqOMFxVLKC1clC3QPFPGiKGy1CQal9kVMP6I7Mecrh3wwcY
zZRDPtkYEt6Uf6Mj/d3IyZWGg77rMZGSG2duLErfI6pJATdWgjMWgNbo0SeZQjy5WVcMez+n0O1P
wbXiG98o1dfRDoVK8+reqBKSAQeEXNYHycMMeHyw4Yz9lVi4RinaSiB6yc+TFpN+ZxnO8XcOo/TR
A5RAHecgNnv3MJo5ICwFNEQmhoum4p7iIZp5sBopgDin/YH3SZOosJGurgxvPJlW/EN/jOZGSD7E
VLLEQWM6Ea0RSRtgOxLRDqrztkZkqakZ8N2PfgBWBslcotvsRJP8facuBMIfvA+H6sk49lVpya9z
IS+AxyQkKq7lwLQSVy49ZOQXFWfivzNXkEWOcd1qJQ7aaLTa2uWtG9/5eSaLFT+zBNZQj/INAsA/
OmNZwtOuMPdOCIOiwUFJu17mlZYHg5sOl0VCOrr56z+SwsG/W9aLtUgcHZPjeFf4YZ6q7n5CyKEI
mdKq6RYvbVOTRT5nX5QuakZKVX7ATN19PKXrmUOh3bB9/7gy/ndfQ4YmBP7m4J5LfC5+gaiQT6b5
msHUtWgSM0VsWurWibtKGvD9eEWrXmoJjaFAVTltK/w65c9I9XLgMUgnWtLfrS6dmWW77WgH6De4
sc8es0xxwNwQXAxC1u6PfWuoRHuC+XnXaB6Z3bfvYYcTdX6Pe1UaOB2tMVyTIu48QsWdxaDrG3QG
4U6afMoEQTH5D+682YwiQ7/3z1/RVe5KUDg27H8cAXQNliCe3ZgkKIL4FjJOGgu1lSBskQAnBXnG
XDscGjpqz1D1iJ4t5xpEf3GwndrmtC4EdzjqxKRh8z4qSLh5JrmoMR0lF+hb/XXDAkU9VXJi+TP/
4Y24qhvjvToB9B38TZSqo4lBnVKbhsw57u48hALT+G1bLTfAtxpjUBJ5oF5ORUl5OZidTV1tyqCQ
KH0QcDTiN9sLC+bu/mu8MOzmWuzHvBgtApLK6FJKfOjfnn7N282JtYCy+9BfcYXwKXpXa9HwIVZT
NI50L7Q4guhuD84hZQJKTU35b7d31Y6d9p+H85k4hyTBYRo+3PUOJC+EfwBfWCujqLSC5OSFLR2k
JBokxvOrMEf91LZwP+YV0JJqwMPje3Xxx6SFdUfxxh6cFJV3r5QEo/HiliR4C6xEQ+kFMy5NA1Ba
JnF9T5++b4YlY6Rllm50uu5vihVKTGiAPrGvEQXn5vLQDS86pqjYVLZNiQR8lExwh+K/iIfE/eEi
CpKq7QTRutNLdV+Zwcc7CGR+wybp7SQ00ty7zPebx7zBlcWKwCX+qOj9mTaQ5N0mSo4u0S53NJX8
4VjyNVIBV19mPHwonUIKGnu6Yy/D12DgYjhbHqhZBLiVLKTBbMOdVk8XJfnfU7+7qsnHZp52CT4+
y3iShja/5KbE2eFrvdBDpSQMF1XeFFgPaKPKpI0YHfBKZJ4ZCDeP2P9qTPrLXUlZBVsa/NyCI2DH
NDz+sW6AQNGh/zaOMbxe+FsKSEqQl5HlQaEN8mw/GObccZUHLTtB7p5opEa/5wgURmRBK2ASCwCU
cmCdZVeuwSJltkmOK68Bxd9yjjBHL1POL9i0EWDWu+0QL4+/brsKy/pbVk2CAT8dRrpJccHlmG4l
fwSgKaxjYo35LJY7Y9HRtHtNLgJYwQQ+pkLOvnF6rzeLXoz+vq1ZcQ0Un6Nb7sAbytu+y4B4mtwA
RxLZLcDYuqxkTeAiL8GD6FiCFUXZtDBKI6VQ6zhJ9bDcNjLa6b2HStB97oM+wdt0eCq4cyQPoq1g
YPcwZnjGkdrThBhcxtJUKeAqvAE2sFd7iG3DrcygJBFlZTy8YW6Wlayz+RDCy2N9qcwE+iGqj2sI
6W1zGY3NvTvR6wd+6qC4aeXq4U/dTV24EtP5QZNctDk6safK5qr8SYk9OgBobIuD0kvoOb8l19Ls
YNsGWBfkL27X0B86Au3jMpatRN/6evABUSFpV44EImdDVhp5S5RGV5wqb5MXOqpenyN1MwqJzjEA
wNiTNmnAXj31Ovs3GGbgobmbeFDRWXrFPlStj/oMCg1ZkZLpSglR23hMO+DGJBUlcEW68jvMLjLP
ZlQkff4GvU5ayglZnxb+BP1D8ScwJwCY0bBAbTN2ztQ4FhMAHIQGx8OLc7qD+vfArX/yiFmBvDZv
mxENkDduQ3MLipNg6txbZYhdT3sy0tz4If77bTy5YIWnAJGSwvfHMA8VyJKPXXjQ9wA428WKTxtv
PhfEZHQRXPgGq3W2GTllVTS9lEbV7nvo7PaaueOVUHAQLOdc5QIPW2cARjHlGn+x7ATPwvvrQf/R
oKPVpVfXyfx+RdjUfRUbgTdy0/t9DAcxTiKfeL7r1T+etZbm3eCBRhl7aCq9jZZLedhJ/1grMBE3
GCwcsRRo2AOZvOG4YYkAg/9bOrDBff4Pr+GN37rwiTi+lW0C1lQM+J2Z7VD7EoNvsJuyRFRdA6sQ
idRauBSvkV2xIe/4UGIy+4HFfddvGyPHvMK2FmBIj4Ei32Fw+lIyUgYEYOqzgExfdZvyVKnkSs9n
xNriwtQa7EkFElNPB8VE2crgms2Oh00AKQqFe1P59JKtOvcNyNLyRIJQRZL1yg1IflC3KSYtp8dr
Er+c6o8dpQc1aBcuPMgw2EZX+q8iHj/03Ad/e/UEGki44VHKy1Kc/13HBF7w3XJRQSgRRfMU+Fpx
UFP7Lh/gr2UPgdUgsSHxhHltlYR/SvTpFZS2ZahC3dCxTSaq1YfXl7WBtLs/+DooFK0rExLtF+AQ
0AW6wzVZk4c41vwJapsEwWdkA3FGm1fVR0xLzLejyy5vPxTjRfTNoKSOXavRJ0ptq3xH0afomU0m
u89o7cdFpH6TD5nd9lAfpZviDX4I8RGky6ClO8/aJnV/yRq1KX9TaNrIJ7dtXvGbR5mlPV8P4pBM
dywb/B12DXNPwmpGAL/9/NP6pI/yGl0aOcWF7B8NhTBeWhvXWgE/8pbVFQu9wZ761VsmDOIdxM/+
uoCLsaP4KJdZoLOlNt9wVETdw5wYZvPlLwdEY6ZoGk++tgUnCvDxJSBK2WkQozP1pZQjGEPKnKw0
6N2vC7M8gqIhKWIKv5Hkd5PkSeYqmCAYlLvTUAtJqzYx3xpo8ayRM1RIHj9Q8VSMyrnZ7HETou4K
1JCgz+WqxkiqLGH/BbwxRa+FJorNVjPJyzx72VR/JOGjCwKuiEaKNjRfdZknJudVLhhh7BYF39kf
XrddWNZoci9lWqxkizyTLL7rE6ljF9fjelZZYkALusSjjNgpkzL+QKy+j4uT6y/DAIH46uP+0Vun
nX6TWWUBrGoeGo8pkukf+d0hcolsJD13wqLxCNJMPVuxDzhImXdUA+Q+R8JHJqsicQRvnVzECB2m
tHr6sgpr1Z+3NKjYZPa9o1T5CWctEidUHYGfilQHMhGu1le6wlKXmDRa7AsyBOSoU+QI5cpZaAr2
DCGQV8qPSGkjGAVAvBa0u8GPlJtl+sGVqCP5u3OT95fH+1FuO9QuAL20M1MZKE8wsWrJjesHCyqC
ZBW6Zq/yv6mOn/iHiNYHu/T6Qzk/UPUlLs52NPMpb8JLZfPpYoChf+931QZ6h60naEgw2O+Vzb0y
iUiK70IenfuoV6KvAKP3gU5B9rjl4iTuz1jwJ+s1nPcSm8pyyjnyiVhKPeh3d1SpYvfCkG1FK/fx
WNAMJEunlVcJs2vNpboHTccAtCVVKwqXeXeclpfvls2PRE80v/kXk9g6UNmTVmLPUSEFQH3752kZ
OvOkAjznfy0UExSrWC5TF0EuffwldQ9H2KqKZxvtaLib2KnZIv0VMEDTAjQgjYXIgYbMk29OCjNJ
nvZIFQ8IgM0MIfNmyLRYqROj+Dq5zLMnALxxGnLshuxplZHsq4fC7MismWG9UupfAb/P7x4PvDFj
0NlU0kX1Z3yjLmUNwMy5ciTyxP+mkODQM093Yk2in1kEgT9K2EYhN3d47coZL4V0Eclr+ytANO30
DuMMysrYJf2Q48Btj7aukdUhLoFr10kj68fpmSUTCIbiWL02wE0G5KUgTFIwCtj4SAPNqTji0UCt
MQk0uKrn++1TNBcHFwlEB1PezujhN1Wz22U5TpvGyp4XV3c4P69/JuMOZ8wO2uFUOfCarn8h8VKm
8v5HmCEK2335dbY36xpo0CkcdkkssUEBBA+fFtLW+5+vFwmyrR3GD/pt14F2gBySkj8sGHqhyTbB
ZT9poBw1DJ3990ti8e0tvC5NRG+X9MxvYerTAE2RFcCvJ0SJfcgLqTskvwXGkV6WE7XOE39BFACU
B21eomiIykcwhq43vOzALL8xjivaBzdlbGIqYXJ44I1ZhITwpEb1kt9g7Vt6Z6BTVWkk+E6p31CD
LMvWYOz/rZVro4wpiHoW+7aKAiP8T+HapHEHXF11Z+Tl7tOvJ423E+qruAWG0fPP/JF3BQhZHjZb
7kIH6SfqnOmYfJLRiE9U95yB5ipBRjT0KdFfGSTpVygCp7Mt4O69Cp58uzCNHdFl0WyXQvXvdT/p
wYqoAZOD6t8LzMdJz24y6uvqaDsZNiVgWos7DXwrCDKodrdRVBZwcHXpyARDXbOVaNlEH9m00r1V
Qlikc/Ax7AkWKpfDyaRtqvYqebAvY/F3RzXMGsl1fx7YvvzQjCD1597TU+kPUS7fyu+oqLUGUYiX
6rsbxp6FW6SFxX5KX4tJGZlFwyd0uHk40IOvk0/zqe6Hcwr99IgDMRXsTlwjHjMHpcJUgaiXd215
W0y2sOv5oGTLZ5w5gKncG4a2cY04zJRj6v9kRXB0DSp3asJh62fqak1Kz59+fQTT2qaB1qETBOrl
ZjlFGF8pyBR9a5F6cZIOVv6WZjIRllp2GdliIaARh+1/h/co3XJVqcJXHfYtv0lzggZn1c+47MLx
SFUXj++e45v4Oqyn2xQu2MwcYfon5abstNveG0vN73yKK7JaT4Ee4yI23BwR+dpNgDk8BUojA9rz
RqT06QV5gssN7uns//R12pxkGk8IFOtbiyRw3sQl+FMuq/ozUZayWby0TXOEPYEn94XOMDIaNoEi
Z6CTVltzwNNiJN+fRGvQeN7saDCBInB1F7Pc/X+GJVcjrkpbed29hFlF1oYhIm7acLX93mDqtlic
TGUDUcEQuEUrsHqYv/2VIzd5p6TUvEmpM8E0TpmsgvZ5E12zS88f216p52E7tqgt9rydLul1Yhso
rCiZy+0eQgoME9dyrLSFPRo+kvebE6XIOe42wR2PiLeAxb0NI/6heusqrI4VueRk9QpJgSaz7LY0
Sxt9FtZo894RM40jpVsO68Ufg/AtQPmBrh1/vQeO3OLE5JpuDJ0nILXMQGXUSzCMDFr2irB84Jxv
5uTeZdARqUqDLgX4khCXuj9d0U3ILj2N/BYL6lsJ7DOHq6NxnYlGNLtlcM9wutbBaPKXIQYy68Ww
uRiyS3MsJApU7sw015xM3EGBeiMkkaAs5h6/sTY4U2p4ePjQ1eFMZBUG7aPQT/WHx7X+RovxHGli
0AVulNquQlKjprVI42zEn0XfLxWJnkR88brdJhii19WinzyS0lGHrx+e7TkkSFrYSd7rcWWBJzIy
c8ejEwEtHfhcnVv1Zfx77jDTYf8vWtG9N+m/och0DH5mbYnCBDQTWLWKK26HRcGBj3xMnIO3bRsy
u1aGZjMOZOdKUsEMUtcGRBp8NESBWbUnz1iq5K1KpR9OEEQDnf/RGJf7X1oE2zlZC5+jw3U9ae+G
YnBesJ2bmnHeGnXEdAmilKo2SPZEuBS7UOWOgtShlhVSrXZGRu6Ne+wZ7D0ClsKb124HVBbYhly+
2fix2AjA8QrHkmNtogpWxFCumkjXAavsIldgFIT2GrON9YGKTrJ2Ho4m5NtgN6UhhixLDf/Kazrs
6fDShYbGlt9kdJepM+koPR50xN5HGWWY3ZZV8VWdc9shVkJiDvvsga6K5TUApeh7j2k5tZzZzofx
Ks6jOF4am6fb8KyINj1Z+h40iRs8Ij0uJDgw7+J6/+l2DmFon9KQxmNDK+Tjm+Fawf452w7oiKRq
vvhKNX7VH0C7y7JUXN9dVv2B5ezgAhN+vpCBWJIFRqqnBJ7Dn8aE0MpcG7dt0I2DYL6DaEUTYMb/
znQw250ZKQ7dOJ/k7E24RWerBfIpPm5FzVDS1Gsg+BcMMlmgLZjMqDLCZ/w+9ARD9ImvwrqaG8ns
+zu1UYhsDnyqnHAKfbRWQT23pm3mZEjuRI4LKdSIE/wo67IQ1rdS3Qx/4aGJfI0kHp58Lsp4VEzd
sUd/c8qfIlQBVGExad1eh4GBqC5c8uXEndMOpcHAi82Nw29utd8RiEpkRJXVC7n6LS81M77L8pFq
lKE942ZUiPepwFHTCy7+EqAIVgLSV9lhgJ0akX6qrQcQHpKKL1DN7K2KG2xouH5WlqI1rZuoRR4l
yUDAbpDR4TrDQOYD28vF9jMnfv88v6nzNOHiQYuQzW1Ojpklq6XE33++QZ9f6ZUrNFSoMKgMxGr9
7iq/a0rWnF73P6P+svcKNRFW/3FOT4mHbg3VTi+x/rRznb0+nrkVXpNonGxBUSGABwIE/Qnyw6q0
7aZmr/ApVr5Al7SHCb5Hu3/xAI+m1e0FzK3e9P4PbekXC3PDz/EgjatLOORy3gJp7822f8a7Ooni
/9VOudE1I/Nt9q5Z9emn1FaaqRcSxVNZWEAKTaK7QTpK4emkZx2U1ux3NSAFa6xE/3EjG+fCppjV
h/EeL74lvbAqk6j25gVdiwaHtLY3ezQkttDLUsp6lKMKXhntRBU0spFWyGIBIz6WEH/M6WR0nUKQ
Ng81luHYgtXZWro1WyWn9x1eCWCeGMnK7wXIt0bk65vpTdxPNw2yNuk+vYTB7TClDzp8LYpHT94l
TGu8Iqg0C2E2ZPXKA8CcqLxkY/zoqg9Ea1A6J1a9NWtCwcJy5n848lmGf7k9UFV843wioXMhrp77
OfUJXdJCAkrb/zad3pdw8NqmpaloVmMmIwEGRFUMtg915v7ph62kvGiuJok2fY5cMv/B8UaGy0UB
RjSFpHMqzRuLDI2LmITfIfDlx+fDieDrszDwr2xZhbArruuu4/6GsUBFyuEjnuA6qUIJ6ESSayiZ
Ianjl3Srh8wMTimRyoMmSNrHklBdP4WbKwtQrDfHhRKEIo9ihHmtgfi64kdwWXzTzoTPoEhycsBt
KgEYW+V+ugm5sQ40OO4Y8JRvbva/MexO7tZasgFzMgooYKoXCbINaewxveHoe6m9us+HjkikY6zb
p/gZAUTP4nNF/uHQIkPqlq7iBNb8s4wPQDzfP7RO7P3VQjKyVXfkyKEy3+LdmeMT9a15z/8K764b
bZuwtqirUt6QcC7yl07PiFZyTd3MUuG5B/R9GFWxRd4mBqKYwBZoR4XP+bMZcL5tGpVnlhiw6+1v
WjZHROulz8FhavOrpqVVZqj6KlzPsOAldaWUYyOi8LNv68Tf6Z3tA842fIqbSNNMxJ4NgWk953KD
0S3mSDe7utrOmkldOEEWGU5GWAuPjbodThw/JTJ28FaUK9N5ZH5kh8qtKPacJPGt662nXeVYJygY
UXCf7vS094LetbQHZGnhiMPrFv+C81o5OHx6HdXQZNff+/MB0x0MpApPM4mbOiipCCVluZgfFChI
EW9A+mHZyXwZHYOdxb+Snj7trx4Gg5sEDd3H2EBHNZJerkIy4orqvZ1umoSQbiX1C4YAlkE5clOT
gFjapeBlfdQmTsU9Do0z3rS1zFLkdUr2u5Xq/8ueX0hZHLxmz86JZJIPeyjENPx3+T2EGoInubET
XmRQKt7yw4efd31ZRaHYISF5HmYdsssiP5hNdNLKv+9zW4NYxcICQY/VD7QN0s8kI85rQPaU9lL8
4eC6svBuTUJntdA7rVVlPdrRQzCMSucK9rGNcbSRb6D/vor1kBTIqCEU75cthtGkGz3l7ADfSKPP
NX75AYSrLVXUTmOO3lc2xfaD3qDzTKMmxyecH/ZY9AaBEySQM6ITYWtJD4nO6U5BYQN2c10Q9zLl
H+1jRJwc7cje2SPPltwM9/A8h/eMvqk5OHcjU/nzpp3jlcW0x1sY6WsL944YyiHW0p8D8gWzJ6GO
3VXRyMPPUQMHNRGWaW9Ys8DP/wJQ5k9IeHDtu7Srj6fIgDaVAxCyfrxp92ZXTZM6X1M1Tph30zUm
sExb6GbEVfVvkq3Xf2nES+NpJUnu9UCutxM/B4Y94pDiHWwATXgrNJX2m9kWlCgobl3zMqWP8ZCM
CiyYgCKIZSb9sXF2102yr6+ImL42Y/RDGMSRLTY+RtC7WyqOww6F9BfRvq788FklCQc4uM+ritZn
R8Bs4OLPG0q7cXXXRjWBG+z0Buqiy2m0+arm/2n/UbsWrMV06Dg8ktpqgvmLgnBSHNGHzwb9hRF3
6b+UXMB60QtNjelqqJ8AuIOxZ+12IgDIVxxlBniNOaZ7auEuMM/5q1DWzocCJHT54qpT3F22lfVY
/xZrCbXWufOKTF4mk7C3QuX+idDLRatMDdpYj1liE16WLrG2Syd4YcNh3BpuLdfUZ6s0lLoLucg4
OiB10QF96wkE9FTVo4FFW2TkJLoRl0iDZkE14ekRbSLL04TBhscvIVv7irhF3BxkCXXqMkPerCan
s4XqhgrJ3FzASG7V9iDm2ol3EcIIKl6/4moGMcG26YU/7K0YHgtpNqEKCkmFhZ9yPj0FB0nIh7JY
PMuuNt8QJqSsvZScN7ejRBlg6aOVygN3pviZ0+vTyLRYMAM4uWgkRs/XydrfoYNWt6Bn2T1JrwTO
xD+umK7uLZv5hvRjNM3goK3Z/3GAPFzr8MIQ8VbnV5w3RSRtvjw9UtPHTnYG5nyU9u/vpL7EwTdc
Ds1nM0ykswEoorMUfxapVo2BLXdwdp+rP5aoJbh/ktOuX22YBWi3ttCSY0Dh/BZkv/EulRC/bkX6
7yIGo0B5+mWpKxHLgNKnH8tpNes0kwPBPDxHunz4xzPA1ceWEhdDSOoKNSLO6udryrMF1kgG1RLG
+Ut7oF8GQOeRegmhio9YMHW/+Br9BhiSy+hyB8iFrkxxvDcPk9Bfgk4JrgzDbMR94J5vaIdCPhpH
gm2jVIvpxnV88avcoQONcD5vgUJ4gHinvMTKqtsFRw6+e5zcc/VBS/2Ga3WtyXNQ62UR76NNAj7W
V42wrArVLJmsMDTNje67VRKDeSBy9ShAMjrwrRLjR+wpzneEJba5OI4BgpefwgyCB/KBL7XnYbnj
PbTzHZKkIKd4m5/1n40fyUEt7Ljpe5O0rkPclmCCrzRHq7RkFGtZPJ0/tB8//x2mR2s/Il0ryVuU
Eg3Ix87jteSzvPXEWJon43ckU+qjBWwr94aYolAYAYDisCJrseTw+l9elY5yiUe7BkSis6GSOcBS
D2yw7YwpOQTfMkoe8bX5aYThQhR22pVzM15cH74etsfhxip4j3lQp6qUCFPRCXRINzY+Xs9/ryuu
oPUGTuOtOpzP01HJYAGQNo+n1M8NshK49cCqqG9o9hL9Db22LjYC1boelZ8Yi+4OPFjdHHc3yyzf
JX5bK3Bkco3GRbXT4sca3V8AhIMP7cSs+b0Y3oGtsWdI+YGCSzRFMftW71oHgrjl4VsVa5O2/1Si
ew7r5/ggqP7WOGV07HlRriOFz3ojZU8HcFEr62d2sJoSZn8nf7i2SS2sr1qofJJpLuQhsFaNMBEy
KoiiV5fCBoxOWb7yFZpnZjb1Lpd1Era1dZoYwA02BDZNum8yPzZMsAJrlnrXZxt6HALc03QyqqVF
luJJn+jiZznY3EBJIqnOuXLyj3oK4ribtQ90PjMg7K1Ia4H93C6MFJtwj1v0eOuooVBopvz5bR1H
yWakCswvAMUmL4hObC5M81BEW9XCmjiC+FJME6+8AeWZuRHIW/OyNLpZuaZWsQwzXMAidvx2b+/s
t/uT1Qy3222xY9GQIR6FWaWvr2HcC5X1fUeigD3aRdAAHH8JkaPz8WS8AXoPBd/eYdcwsHIU+8gS
FgHWPrT8+uHC8aI5vXte+NjUFMSf60liXlxuYnz+3WIQhW8PELSEde1ILq8Sshizh11SYdKwih+R
JGaGsM9cZwzNpOb37CwVrwrd9zQc97ZnWj464YkWIQa3ZSbeJJKc2wVs+iRgf3g+HtAJW9ETHbsL
rgzmCAQZxI3loDmWgdmwEmXthtwaiba3iZ8IYQNBVcikpHbRw3O5NjzG+Jyj6bOV8QHmqNDgRxNm
bdWZwvY9Xc8FskAUl3zWbVV/ACZhywwdr3IorCmdyUm+HwORpCfm2z80npuFQ4WqB0HpIA+HEch/
LeRIhOWxrfVDVwbJ2BcLgCUmNgirR40RvGo6wOY7QajL/cbqEHLRBqFnKzI44F9TrwLurIuiBm9A
L35UZZvniBZT/9P/JctEBCPi+QYoFtOCC745OK7zK9No3Wf/jwTezeLeCOU/vDNiE4RHrZPx0jfw
gN/W6ffOkc/jk1AQspUzQwoJs9GBRyp5NFc7wivFCg2uFCDzpAow4HweLx26Jb0iaZ5aUUaRsl3X
uiAF4Qq79g+6PH4HJF9Hkn7FDEx+c6yp0gxJ0Tp2RGQ4trcfv4xoJzV3GJAG+4iYs70+Zn9B5uSE
jjA/AFztMUqCJICuHgzaNR3BkIddgDKT2q1D45m7T3NbwSzy7YuKfMOjMI2QAZABHR9QFxXZS1Yo
GRFJEFfpjlg+UJ3bOfNoY0P4mEfftIXy+3FMIarDFTEHXM3FZmy67x6hVT6j4UPze6Ncgu+z0WaQ
yAiAy17jtx0IlyU1S0hxthW/3q0z8ZDtVD5b7uxyjCW1tNJCQQxEwcuLyyKMT3EG93DfgQNRhUIl
DggDqK2EquVRChxfS9qrns/3f5ob1sy34QBTPd8ONEpadWUy1GcsVGXFYG+O9w5R+6m2074vEKMZ
Kvl0ct7cnHbLuEEQhq3QhdhEYmd9aIAK7RFjSzHsjvoKWCRibokhr9Jae2qlfWI0py+qDolki8Gk
LsevG3RrMBGhQW/ItckPStNepziv3A+E8coiYPuhqBmefdnJyfpqKT+veKluFQZ+Xj+M2xJGKIsf
2GJJrfUdvHHW9gMmgJE45UHOy/B2rzkEoTRrrlo+2ONXis4Esgqg1fq0t/jzmSGv74y0NGsboAwY
OLShac9UIlZRdf7wBs7YMglZAvfxeAR+AdC2G29t/KXjpXNd+PSoXxauuYvF0Ehwu9njfygsALS/
7mOFTI9Bzp7CsjlUyKt0RV45J2P5ighF77Rp3DxSDJPJeDUOFpAvBPA8uqnpmwF2YkjbwBkNRF9Z
0fF0aanWQjNlQ90DwpC2OQ3R8ifuBbZZ2SsHaxdsIMf6YfC1p8zOVDVue8+DvX3E8B+1t/rd2wPd
ESMcfi8GocLbGhGC4kENlRP48t8aOPxUqcfHN+4mckGTWEhkN9FRm6/r4ULKrJpWf1DgHR+CTx7X
bHPAM5fnatJaMwMw1FM8o88bZZXb3Sg+qV3zpv3RTw9q4IBt1ffgUr39OXhTCnW2kpfFkJ0CkRTj
67/aOhKl0yrb5G1sBmz8zh39piBw2vXc9kfCdgr9jQHmQXz7R5ivNsuMkAcGcw9lo3NlT/I8Qahy
XTm7Ny4GUMlbDUpld+GBThRmqbOm40Jeq9Htdhc4tqhr/gdwkBa451Vsm6/rTCf+zgWDeSeWbkq7
fwHzTgZbnhrxQpV9ljZhzaOgFy+vaIsZgXhCVVXr3gNrYvX9py3gtYe9kFlJycK1rEmHE5Z92k/W
LQBUi5i96NFrv76WsUJaGE/IL378gvqdycCbvUlVlJcaaJ6cmjeSDobvtLtWtC/x6gbejSj68nxP
JggifGn37Zhja00BbmsRSUsvPivyOxBWbl5x6/xADI+rRm3C1r/q+oVo6BBcUQ1wkx4zm95z/H17
v+uhK4NtRawGN8AMeWj3vN+h5xCgVi3sZr0t6dAl2p40rLMtZs+3e6GAPHvO7inlpF9Q3avzREVS
L3ocCtByIjuDKP54MuFCdQ5Q7XK/YYTGqwbwbNpRIRX6Q9fVTyf6l8u9Y+7urBjni6nyJ9wbT7W3
YUNzw4CFdUMr4QaWjGivkR4nNQUteSHZ3HNTTHg8k9c72oIU23qwnVhxKUtDpRtkhxWPTYIUlIAd
oMk3sd2/UBX/7ERJcVBMmf3bF/Z3oT2Yve/RDhl8bbxeTMXGEiuAAboA7D15C+fI1Rd77RwzYc+c
lyDEM6jsL8mQixVtgIdZzYehIxxdkmCdfSmMUO5eP9+FTQai3xp65ZQrGVjFNIBRloZbAuUIG5zs
kC1EDKWWNGSpLopBXRXJP0o0dZKBg6cWdBswrpmmCYLd3BGAtPyilaKBbsS2NJFtnqofuqkVngso
zvWj/YEbjfEpPXsYCSyxSNxsEzVOM1FnD7uP679NtSCz5sNmfUl3+7A/js7x6kYyJMtIhktrX64d
yGEzTTcS3LrEVli8lRtecJ2UObtkbTOpEu+Q5e9UHOjRR6cF2i0iyjNxEv/dJjag42ZDtJZQhX6c
5CF3dyQMIEzImrXbrix3qWdiJz0xLLXspZQE/aG9HOGKUHPN1hFOz8eTL8FTe35kw3PRatJ6PQeF
rsUrZjzN0Hfa6EmYmPXpUswps2f1Ne3mlHlpbhk91QvBTnA2j3g5VNtSjBRJhQkF3MCHN/lbKtI/
6QLtSjPOEpll29tWTlAppGxe0/g+me9jNW6PC8sbf4pCIpnH6k6zIvuq+sCyMH09kcaXGc8CdxWR
/E0/BJYSdPi20SaU9TN/gvT8XnuuzyHzg9/3HS3ugj5dp8uftl8MOv107AEiIzj5PA6WpiOU1VZv
Op7r26P8V1tezfLs5Va1KuZ+kTpwPFqhQfPGjxEb1RceQqQdAa5+vsFWKmArHVJEK/AkwM/zwYh3
aPaAd20so1aEOw6hZkcIm/pGDUkAjRc9CAZs/KZkZbudfh6KVOpBTb4wVyI2MPV77guNE+WS9nXI
rgoK0MVLgxcBCKYiZ/GmokJDMIur6pKkOq+RDwmHxjfkIeeq6v1YETMGM6fIte2q2KrUhVFl6bi8
u6OLTMEGXEwrhrgzzeIwzaUwkF8MPSmaryuTJn23nelxIDN+Kzv7Ao91dUvkZPeRFrx4StzIgNQW
HfrVSHH1iDRxx360EaJ1VHEKIogegfgn22/li6KnDWBvEuL+UOYyaeSREsKel66dmy9P1aikg/Ej
yjTHEhh1meA9h0QuXkMOQ4ONFUdZ8/2HwhSzqk0YEndtrVnHifokX/3wrGN1AP5YR4OfjPFRS6DS
PGdhmKba0LUhIYg4qtADhgfvkEJ+sdi38tLUR/3/m+okF1F6H3tQQMu3RO6prVywVGVTPb1iqsvM
GIO6AnaGRtOJf6Om6HiJdIh4li/Fn5b5avpxtvcMFkpPxSqlalzA8hptT6Oip6cYQJKIRtC/tAmF
+qUGg21DaW7E7n8rFKR3pNcQ/QYoWzoV2JEhzyVx5n88S4hF0p76nTUZSnTINEjMCDIiRxu/rijr
CBwDyPW0UFtWqXDE9Ov5D9rc4osWv71BwP+2/jpT358bZEVj02meUTUqNbIxiNWSqYqqKGW9SPKL
pLQvGEdNIURYcdPTHFR3J4Wd2zgZ1FzIBGQtbn/7KRzH/RIuDmpJfFWTWehM9S5MMWn9vfClnl6s
QEUevAZlxq/VAXOXBCMPIFwzBEa2auA0DAUU01ExmhyTQkhh4c/ROz7F7I/Uljr1mu/kY98lMLFH
iIxKmn5gR5bWvPSCzdM5ML/pnm1UtCPTyQlzrzyAljg6dExeMaC31es4TibXBe2tD6QvMEG4kAUK
kT45MBrhgj1NZ6qJbJh23d1RlxhrwvPDDcW4IyXU3eHfSo702jr2z87jNBjmZBBDbzvVDVkB+D2B
yao+GefG4e2GdjMz58OPDVObGA79480W3X+zz+3s8icFcb8s2bZVMjQT2/hDz/lp2Ljl1Zu9tAVr
V4FF6CQ23FVzmQsvWVgX5X3Iig/1xLMsnsCP3Z88EcHfLIzYy8Xu19hd2G/FoUkMdNfd+mInuChS
L2Q3Hl33Uv6+lIQIEjhsHzbULoGNic8qNomKyEgVjBFwdGFpGLd/VwKauI1jfcHHKuZzufOB5HUv
iVmfhNx3etHvd4RZV/SrfJ8RWooIgOjijNyuLURyB7/XeWniQSEintyN78WHYISowEF+Bdwp/6QW
gGd1aXqHN3UeyUi3bO0/bxIGpyRkjyLXQwFcsxVcPhbjiwwO26BvFEUhwp94o4AjCiE3FG9YQag4
suj2f/7Hjg931hDMzgpxx6tlODS2xhcKj56sJ85vBR0mLUYtnnnymjJBqOpjREowAxkbxankTmzt
LgViiQ7pWvrnoaCUruLsBYe+HAMu5eG3ev1X0XiCloP7faPMjGLK/f03Jhdjtfe0UGrLpgViN0No
ZMrO0otEnFNzYkiaEhonEyMy/mIbb8fJwSzDDgjyQcTErUuZIGDe0zJpeAwvz+/yIN1s0QF14gkb
bsnF4pRUq0kDhSH2p5lInNb0sb0bmh75RgQnB3CmvvIofIPwMckr/VgtlQB4CernjpivlpDoeLRp
TQ1jJLS8MQLf4ooY7EiXNcLqb/Y/EULaKxErSpaxndepLbeC3+gxe6++YAIGm8FNUoyYm6Pl0vr1
FHnEHBLbBc9SRbBbUGyYpzA1eCTOr5aRL19QOIsyHQnTPCX2BCJVQfSb8oelHLWEEulTTFaXk1wJ
4s24QuDUEU7Ckjlifp+GI+8kpapUTpK6BFpS/Rcd/GPLr079Tf/1ShEUwDK0PsH0MZOnLK2Fsyt9
QdB0HSifFAAESJVtLi9KKLkG66CFe7bTlQiYfgxduuVOTc854UjtC+lPsrIOMuLKfvP/smzsWAva
SPyaTYrlViD2j3mMb1nzk3vkfgrkLkwCGQ1xrbkRRJW42+JdEbz2CorWtDldSpcRGRiMstRHdV0x
nFzd0pPVlH4vho+WTPAUWFEEvpvMJ++vSBCtkEVABRTsBBxeUz3Fb8HCLepnQBN7cnF4syrl7jfh
Q7ucydeqZy0erhW/VtEcq16ObFwuyzRVfi1ELJwrebC1PKYR/wZW8sTglXwH4bMznC9CjK+ceZzB
X+wRt1N4PQSgPKdaS9zb1rblr85baS7/xfcxqSW1AwnNyvFAVkA5imRPTALWM6XA5FCb3ezIg8g/
ct1HDmhjE0iAsa6Ogwr/KGHRZ6zVbcnCnQ/kOCc6+B33bFZW+CRpWvANAVv9b88JcDit0dUCCNOR
a8j1Q+80512XuRHv3X5dLUl6oTzjtquhAmU7I0IOtiMrWQZSu1pjByitARc63nkUD6ROcG+phZS1
UIfyrI6SbyXwAr94TvrMgQpiuQR2tA6HHdMcH3MApYBPZPoDcrOPDQxUCO2uKMZchEAfzutN+ajR
nJxO9tTzSs3QqRw/Q49cQxdKXlTE80OlvV1nWqIqkjyx368k04PJEEj6p+fhP70liTMYKOi7J4PG
dsJnJOXqy0sWlUwoEAAeyg+XO4NeNHt9ioIFjhhKU+YRl8O0oJV5IWO8EZ+wYwy3LbyA1R9XWMdd
r1hlseWVByx34RlLt8Kys0CeS2g64JCGxVGFRUMq3PXhXJ/wFH8e0Ry7+V4l8MFRtKwap2W5axZW
3gWcLZ2K3H02OHxJAaCP77YF9ZUt4jDcbUduOmrsBAPuf2bKdNthFAmkJMyAak2zn7J4NqS7PYTY
o5EyXJes8j784CElw85E7JnDo1dalnCerlT1fXs4Wl8jsO3S+gOKgXocQl6Y+i+qLeiF7ssCKVU8
N4U+sW/aaUgKEuDaffVyYE373/DwyrqoxfAXnlQ66ycntNqU9G5IkN5GmpZ+aKnay29r3YY2N7bp
hAug8zVYblI3IRSLhCEKq6saBqHAGLqr29jXQDMS6rZevTEGbnF8OTEtgCw/LB88lMBfwv+a4+GX
ogyPJF9pI7hvCMJlZaQwntejsK037XpVHFnF0fri7NRVAedTxyzsTYrB86rEYGYwZIFyTT4/MSME
voqIpullKkJKHJOqO2oKmIdxqfNnCIwpXsCO3WWk9P4mK7lyD4wvd96kD0xN8Aocf6NnJFkQEEwg
vAaOVms8sYOlnBqy44/KNnYb6mLyQaEfUgGos1sE73nQoQ0N2OSKrMZECBtb633Qjx5jthqXypQm
Va41aMuHovcW2E/1qoYa0bsQypPxzzX3g6T0vtwjr1CkqZlXnq8xifuGQbAhBtfD9fmTiNdICOwv
5GbZXgpiR1QP1AixL8Svge4x0NOvbNQmN7kn34x0Xy/gsq6l3vbYVU75WPIyBYllEYOKtz3U/lb8
kDDs56BmJAtSrS+FDCxUMyLrLxpv7WO1G2qPCExJMbzgZPuuaECmupolf6NECD5mloy8uDq7OseV
LxN19ry22AGb5IeLSMY8+WyH24Tyumd37qKM1gHsbUbfcjo8t+gkheXro1aeEFjsoAWhLKPPgokl
ftSuwkSczhTil25t2ZEqrzXIH4oEKRdyVSg2e+IxVyKc7CM5H1VAnc6d5rHVdqTTgyhQ02jR0Au4
++vBuNxOemnvAY5Mw+Or1RMlmKy6Qg8lBTc8qndtqyJMRPkVMpxWWwNaNiDngmthG2P3dz28kmkB
lH7snFpt8q0WdxKpjV+E8+EoE2sqDl8/1zE1u7/wKSwOWuytp1Hpe6ITQO04yhFy1PGjPe1IfZlR
roQXVaTtghfq8tn1/F1L18DeSa3gE8usfIDtNSJHGxTYvQCX308ZZdBBdGBOMyNRBDR96pMvD9WB
5nSfFLZ8nUiECOSLgBKQhx5eVJDE11qbQo9RlAhj5mH299Qn5uaOG/IKptSnd8r9Nlv9yV5Gv+JW
PGXMVCapbKcqOymyMxH7m/Ik+ofzZZC4F2iCc/o8VCzjDeJ4EWYb9mHgi8Nf944xk6yED+c7eoOf
siNDH6xF2UfLsZhKoOmIYqDrOi/GpnJn3yx6KDk2t8HBn88f8F+WJmYcYK+8diyrVOhuH7/1wJjH
7zq+16yWLM55cHy7x9RMkCKsEBRh9fPUAf1GJZOE6veQh5epx9Fpgpfyf/o5V98XQPHVniVxq6Sw
ZDcwjSpRL8amIW2kGq3skku3SGiyMIKKtXXpMhjncOShQB9pjKMe4LaLLWujL8Rgqskxi0kQjtlH
dDEWF9mh+4AoYHHAJ9falllgv/Ak1hIPgh6HgK2hmTWEZX6r7emjarU8jS8rWbwCF4wq1HcvR7mR
cxg1ejF9cbkX+RuGGtu6GHDT510b53R0pAEyd3ndm1XKi1KYiLnXo82mQmeETJDTZLkYzsZ3l22l
9DS46lJTCoSvSTKMljkWnXF9XOgHzP556T7/7eU0rCXKzUt0ek1ZmxUvxyP2y+oElhiaRNgZmY/6
txeI7cjTiG3Mg7iEI7R49NRVzwZnxCJCz8PibWoe4NGpKGjRLU17UGIfWw+84PEhvOXN0BBNNWpd
FbhsgSi2tYY7zmZFIGCBsr2P36afT1ItFrcpgv2Thd7z1KHmqoSoMesyi7tXTCaAWSN2ILZ5LVMk
d5/S9EaMi+g8Evgo47Fs+arbmWq0anQ75uNe+y5OgInkzTD3c44YRfH54ObPj0L96tTe+SRslORa
8Q3WM5i2mVY5A9h77dtEk1cYBFcG2oLFVuXCjOMgd9HiJH/eHMI+8g/Aa8yGQ1Uh5zjmQJohNHkS
ldcna9SMP5het+EysRhvyrWWxk6iRzQg5VAYuh64LP6wxLrlVX9k9eo5tSFwtaYUn0K2Io6/j4uy
PNvFPsXGoAQt3IZqvjwXbxYDhSRfpdgTvNFnSBlQi/EGc5/wzIiR9BDNisK6nRcvRyY+vfd7oMs+
tWDHjYx4WA43iO/pULoynCOe/+ItKObj9sZteuXPtXEPedCJprqMprdi6BunMzq9B3eT5udiPfq6
MNdf96e+EjcOrw9qEBAe/4bUow0LoBQuBrFP7XOOGQom8v3LbOcb6A8fWnHglwhxrhfZgJb0FbAo
atR1hoCpGEfRDA4tzw0403CVZvehLJEt8MkyqBCWqOXSp/Pl1CcTGlo8LgJB1gjrS0kVHRPWrxos
LzL1x36ny6cfZJinHnI7OGqG6ysVfp0i2flkwySseN9lHrv3N1EJkxNfb8RqPvTYwbakU0EO/F4y
a1HeWdoTWMR09hxVEYv/mTrTscMafz7tRv4pfV3G6mxlpr8yJBBszGF/5xbqgjo1Z8jGr8DUmagm
XS6pGIau31JNEfb3GiHiMeyme+kRfewf8uuZPP14rEHQ/1S1cx9NeX5sL4ydQoQRYpLHb1xXUk6S
B53gfP+g/hRrEVGdFsY2LmzcNL6WH8MtKH9TlOzNOAZRF4HyXaSZIkEywtY6d96B3upkj6O2qy36
kvhJgFbF42tWvNaBTg5tSc/bctP7O1EK2HHA3yNun5LWRHfOujgrSLEGq/HK2DPPTQPzFDD4xmVh
d0s8KuWVf6HWwy27znX+9YXWLh6e+iqKE1aQ+uuVZJet3uoqpzTYU+9LFXOut7lP8NFrV5jMNAgy
9qjuzxc8+FhxSbDcD9zDX2W8wficQ/K4jvPWy3jYfJEvZzWPyevcC8irEVTZfXQWcy+DybYAj7Tw
Bog0r67YjxbNCPAIf2w1rT8tl90TOo0lSumuaJHWJmc/CqmWqK5K7xlfHl2VWvm2/eFOAGQqmPop
c3+dAqcicPUXXViTHIZm++ji9XpD5LdMo3b7zXLdtoq8mlRp22wloJV+wTOIJu/BPSywg9DDXwmA
mv8mfTfKwE4XzG2RUPkhsVKwZ8U1eiqTozI2XFkq2UYg/TJvpxbnc20trp3xj5w3QjDI32y4vk2K
wY8Zsrh3lC7cBifEsud0Fv3DGZoaom4/Cv6RHMbis1WOd2Nph+/Pphqsm3PzFqfa4h34Rg2ioB+6
k0Btc2V22gP9P84pEpXtex+X2ELJ7lXxMAzvQzqYLk25XWZzDenKlxv0X+/zW+ASWWMAwRGp1yL6
cBcMRGLgw9fjFvz8O+ntQnCGPGFGiUfxxaxhOw8kcx4vazqkJsRpQhgbYxFGWjMzeC3x47KqjT+v
RKh13WrA6WWx4IC1GhLbZlYZe1hwnpWkiwD07YaQ3Zbk57dISzZwPPL+mpdq/NKEL/dFHHbYcWB2
7kWEsJtzmG9n+9aGd/9UbjGGhWE1ybSnI+mObT8IEMSSzBEhIlYaQLNulrlhmt+DnfdV7S/YqS8k
MStdkLZOL1l3VcwHr0/hgWEG2CbGbW4pdfMqdtzP8Ygz00b0entwk/qNdDZEPwntqk1wSW0f0/Vc
hAHrdP8qYCI6lD2vjPskxnS4vbzwAOlaQK+J4tqoRXXYK/w624fzZdWHIH8k4NEBXAYL2joOrpYo
EkVvqOLmQ0Ko8lwQ1Q2H5bnX4fz1NcFbQUgYD3jmTPS8mKlx9D1bhABxBlUhyfg+glPImq+DFOe2
E8tXG9YBi/w3RIp+ut9DLYPPBHY0QFkdpTvYRO3yTNHOync4n9a2iSO1Fq9rQscAPf/F49YdixYj
1riy8MBxjLSPjBR9ZhR3BM1rEe9qNaK/aRGmQQeNJ12UkSvVznT5P+t89Dih3CW5uesuPL1Pda02
OjMY8JdmsOttkETxvSSj6ki8wpafFhx+LWLc5mCA6k21l1C2npWMSzKEW9JZDwQllk9PsJaLecBt
P2NB1ALl3pXoISFuudBnJPNI88ShbcBNXJKzh8+e44KSHOe7eNEPPjy+Zf2eUETDgL6YGc41UTJi
TeV8vNTYMfkm2pprzQRr82OqFNbvqc+w3+TBe0DK0jX4RDoOMynIs1cyzWs3EOv6xEL1BRm6WPy1
ZLXrz485PsR5Atb99SoJa3JagkZ1rbuei/YsJDHUAFdO+ISv+jr8SrRPzVrNYpNA6CI6YlFzebA+
27CCZWQcFEdmUk9tFa2MhZF8o9jMIpzghTsQpecxZZQF16CYVLPdiberQE7YVPj/w9AS0zHtTJH8
EUn9AKVJFu3X05TeMTGEsHvJ9ioKL/U0idvK0Mkq5ovj2dPq7q2hlheYcGk9d5nzobXExyJfvXyD
5xfVWq8sacqNXiE3wsGHKYfW8Eg6NyMfnUDm2MNkQh446vmC8YoVAMZVf7RCykUPpkqDITjrKIOw
6qtDDonvotkF1Qta0sd/kW8wCToJ/xwuFXY8QUKTDs3GvJWTaIintWPZdm1lSdZj9/6mZj4S3VQ/
xTKw9Osi+SPvobKiSlslXyl/TgFzsPGbIt85cP85NgWQlDnsnoWyqmZXBf5s0R9M/jW2ulxe8kjC
ibncj1RuDVVsLrB2pVWCFw56ARCZSSbYisMueh5for4j0jwxHNNoZOGBguGeEK5RuyTHFn2dYSjw
CcnLyO14Ci7ZE0JQ50D58XoFo9DXab2en6XH/CYPS+SioaB/dwASCjbcTXNls/H63v7+TOxJ/uJl
jpJonsBOoCeXrpXpzoefjRiweBo3E3UBMIkUqorgBwF7aTEAw91rZhEL42Tj5y65jqWPM6jR5Eai
JXbT8G251PYTAYzVY6BobbHlBEbowKUe1XLVFtwaq9CcIGF6MQ3TQUPgO9XHl93jda1TsEIdEfOz
qt3Q7KwAg8i+AJUOrA+vxiCrJ+24x9++z1OdtEXFcUcluCi7shFkFlGWcao8cXiA/nhLNReOD9bW
VwT4Zh6na9IazfUO0A33wougy04o3G2Gl1LtCPR7O8hQKG0//F5mH313/8PiLgqZWAZbw30Ad64A
As1fvTjUjrtFmLPce8jfhLED2cTSi8GzVu3vitwmVDA5e9MTQHD/Dnb36Evm7rxUVPx+rcDTK04X
jR7kbgIF9xsxjzxZpDiBGgG0rq+vjr3jr0YcJHiU/oyqQ8bROleDOdW/0ad9kpM+NDfmh8sHVzeu
aNF1qTNv+6jEbzSLa6XN+O79mzeXDjNecBm1nnxyATiRuZWyM47iwdDGHBTl199r3vNeuxupOuT6
hJR3taEgEjDCwE4YlitZD9LwlN4Pm/JL0frB7gRQo3dc84VTUMFtaubsDBG4uNfdPLSy7r3LM34v
drUuH4VfMxsRufSlbyI3YU+C/T+wSH/wt3XVD1bRbqgp5fT8SvLFAkJr1NayySuG8JLuNfvWAlGK
GrQV5NZpp8AgeN2wCIRx04iePN5CPMOaPDubN803aM/NOvWENksJQgTqvsBudaDap+T4ZUiefAcB
iFNEddANVkqZXK56LGPzzdrk3+CH2JtKoRkWN7eOBvRXdUC13PUTfFvMxc1UPLs/ZSJ8OV+4RxOa
fFbDgPhx2VFJpRCGwBr0wK2oTtYABRRZIY8v9FkywBbgIXwGorUkGEOChp+u/zfzlZipmAo1rT4q
nXmow6xyRXAARwdkIscPY/w6auPRAabZO0O97bDehIfYtYsfsG5VWs3LTNjjlI2eqSlEwzZwAIjV
82X4GJCk9kJo7CNBpFe0xDrPDKijKN1OpP4eHlDwQiDRpiWtd+ksv01iqvk3qfKHkXmtB3zkWfND
/gG3K6CJEyBNF81Tb3pWYa7unODsayKbCr6x/DtbLClvgiAmPTI8bftq2ZA69agJW18CAFJ3hh5r
kjbWI/KBr0VHa++QzJhthWHeUdYDEh5SiqvtorQxzMjvFdgcKvXsqHsueFuiyrcqSil97a5Rb7kv
TaEBBw5jTn1tkHl5WZVbfuOopL/bn/0qBDBbVA8JHXfR1yrfbBqhWVmEZHaboWJD2/jn9i5dj56z
PxNF+ADAHfkZIvFkKmtkoCLmEsFEgGbunrjHEISXc/AvJAqjDY+NAu5E8D8K7cM/ogneA3oSyqiL
PQobJeAFVWIiuftK0YVDhGuPmP4gyfAbSRsDvOE6Pj+xuyBql4+2L15EmkgCYiPNGPnwhNaLW6kj
/4UsgiIt6+Vx3ZM5dowywTRWkh5sBg7DDrLNvgnn5pAO9DgHoZoSmXq4bR0wc0zcJE6X45F20NYy
xsy0RTBnPA2BoaIZceOH0oeIzFyENZ0FjciGzpsEF1G7VDoFKCMOe1luteo/0/LNEuXZT6n+GoyO
F/RQc2jQZKlVzwRMx9Kwp/wmSV0AVJ1G7m8b9LJXXVfZDGlXR20izbpiEfsG6rRGnETocr5gKDBa
y07MJ0uyDw2ILM+Lcir6asW+2JaN7cZrHkzE0Ve5jq/VC26s+dVk+AH9mrorxgTFpSAzAGuGKyeP
CrAJAyPUsvCQkQZEBI/pBd1ztrTnIW/7Hw++o5Q3/UYTDEEeh1LuG17904jxd22b7oTDASjP+eTm
gbkJGuVLpe2ON8/gpikBzrCz+BH9m1YrYFuBYRSDwqGt4ZIhpZmSSlCccAJ1WqsPOtbLMXjjTaZc
chgqDNPEZ+yN+cXP4VD82J/Yxa1+Cc9jPPslRjQ+kxdu/9ARM1M5DrqsxVOXMJClGv3hwMCrj8HN
pfSVWhkzEBHZN9bvacDyKGYQIjbVlFoqFuaBR/j/4A0tU4wQOaIAmFZ7lO/UDTh80b1oqCC3xHbi
Mib6/kZHnzA4U8ysbq2tB23AM4CLTK72tup5r7xqh1wTIvuACc9P0NyNl7uqKm2riL3sG2G5Rapr
vkMdLIZuUxBulNBfdXwEArMwTAGotwEcvVHfDTpJ/nB8l1oA8E1cWhKnvVkK7B0qghp6VZPIexwB
xMKEh9hntvbZCdtC72z1Gg0m+ZIXESsdRXIFqJsjap9xv+OuF2cKsMPYY4jzLk+1t1s+HO6Zg3RJ
h3E14MQGPSntyq5tZw7VHoxXMmAsFCU/6sV9efGCqbKUTExdc4zScMPi3ItrVZs9+OxHWaN9IiqD
ncDDKwVEM4PJXvvJvVcA8KC1kRG5SJzzk8H/HEmL9IorPer3lLoksnG8OceqwbNPpFsOruU0zqhc
nJEF1EZJV9CwQBVSITfQ0VE+FjVdrc2yPfOCS7+og0kB7xdMWZ1hTW/QkXy559ACrrFDyDiD7rmE
hBXCiIPok0y75vTL+kz8xu0pAr8DJhztsAUel4mMPB3zC1n5RXjXrzw/o4rCf24g93LMl7rP+mZB
rbwaoc9oCxBbpzYIdK2Qa++cyITglTSFt2fpUa8NLN7a42jZ/i/T+O0CsWsu7OxPLX9dno/m4New
dSg/nG93srHtyLY2SvtZkRk/XL4lWaiWyElRiMDBAvrgyfcu853kHL3ZyHCyjoWAVLbFRatDe8d5
UtwoazHP4gW/k0BRpErwc2PsMTzO0rKT7GOptqjXdnNttewP5NOztEC/umjNc9wHlyLJ1gxZtPMz
x4M1DVpFnfDWRaUu7jkZY91t/Dg75ZoMw2kRQD8dXOc9irOOVCRnM4P4FyhIiQGyjQkFlSejlJpE
r8j0xWkZ2PNTZjGGwESw50BOFEPE/ze4bnaRt1tOeWLwjqgMnlPDEzrkFdQF7Hz6Hby+qbcBu+/i
Y8JfD86T1AeEZXkJRXUTGRdfPPahHHhVlQI/fyDbaJQHHohOgU4F4sXtdoe2zZpHi9bjaV2ZX4at
SN3xHA/IrEhQ8WiMJXKMbpCNZwCQG9RiupzGnan5LXn/iajj3O6WHzqjonQBK9Uwv9XsM/8sxCHH
2nrRqEOFs8xBDuZ/K3KwnVjXaj5FDW4ybXrLU9fERdeGI/vn8IBbkdSZZKRAH6Yb7c7yjDCrGHU6
4qQqyy7+AJffOVKF7oeKyYyCOjIR1QEyp0DriZgfQnA/68oRlsfD/tk/V/WDFTGli5a70MRcVtrU
KVmAsfdT+/9G9CKk1YbO2M19Yc66b/kaBDr9B/FGOI5SfSsuW0u4eqewZHmHTorsuwofNIvk0Ply
k5HOw1qGHdN/XBZvZOP3wfsu3GxoPKu6zCapkJRmBhYqzNZ4NMLmBxIbBZ4ycrvL9N9R/J3UHTvI
b4qpnelsWlqJOmzX/XFUx8jFNpygqubtU0twtMoBE2h8E8dJT1UZxIV2MSsn6d93dcbvRPtPD9xY
EJLoDC/6dn7tbxMzm7MBC5kMjteEXoUYTtWDVz1KElOhGRer62ApP5ylFh5aNY0RYocnfgMCfM2M
CsVsoncJWzPo8LW8+wDJ9iJjWGw5MPQli69/boiGxyqIoOQ6RM2GkOSZ5N5H1YT218V7BDIgVLmd
a4+2Oahx4eIBYFTNorqEqDTqGaJtFCealulWbNtiPXcfdFSmy76R0Ge9FJmvsNZ3SqAnM3GkCToZ
mXT1RDDMk79Uq3nE6kqiu4+IWP897MNPluQ4Vwc1A9lXCh2ugKFXEwqx9jvPvghZUSEVdz3z/onc
2akWX/vaP9h32qhXIrRKkUCh5J5t9Wq63vvj2r3CrpCm3XDwq92xz1HFyK/n5oyviKRz2ebVkiQg
TmcE/kpdJn+ha1UgBdNOmpMcKekYHvzQTsdfMvG+57YLKeJv0n9vFiQrJvYQH4H4RWMAONthEPGN
vZVr90TooCBkjC2zRA4BeJFI6rykq1F4jnfCSLQCIhLd46JIPlxLWwUyYdi1qXWQnwx0jdiFvxiw
5990W2xU8ajY5T7BCJsMQ5Qj++nBAINwWfyAKCFw9xtqY4byTW5zwDFO9gNFLF8mAtHPAmty+uQn
105Fg6j7zS06qY9Sz8DVbEbPTr+zhzWm+4odYsqI5QAO4I5nB/SS+J9GrPTSuf8z+8tM2QHlV/NM
l3M5zh/cfL+YKKKvQbkE3wRoRWjdfwLAasRt64s9xRudxVzIq+Q7/oEPOEDRahavFjPef6CSnQjk
racdVWbdkH6SM/keqmeot7dbPB+ESqfyXqKyQQFhw+AeX1k1QbZsHYxxdDIC2ykW0CZC2jluddSY
6PrkrCtc1u9XG/SUGz4dRRTAkZNQSTXENRC39jrnIH9/RPqjfi0locwC+2tKLpJM/NH6ucVoFbUp
qpzJBJoYbqlmuTEVgokryGehBk+mYBMki1VW2i7AZuNawKItBTRSNh1u6XWlTUd/J8VN8IT+Fo2T
zA/nrtBjIboNj26HPk0IcVEJsGWrj6cEL3Hias/zrKwIjWrVoDdwVkJETZg9zo2x63DTwBtgyn1e
2Tnr/O4DAZzlwDtkbKIIAgdsGegbiTA1gdq7EIxPfI0OYod9WGV7XE54wlmVnt7rZmtcTeqewfCS
28q+l15ID5bfbGAX/93EgQK6FlvSpAZ0L6aEWc1QhQLCQ374T1MxG6PE/rkq0gJ89BtiQhMLo6Ai
sMd40eiDRro+NjPnQb7F+o/jLCxOgOUrsPqtPi5Idoy+f0lWFkheYCBlRY23XtlTzh0t6ZSxmPQM
v3LCOroRlycIFeGpgpNqOxlO9GQ2/h3eLd5wowN0C94WIsIGjE2ZwubBwvmQig8rsQB4aNv9URz9
XGBuoIjCBk0wMMaoFiuYt+bkB9EWoL1kWBuKvyjrPPu69hHXzcBNLlFmuNwFm+sWFjonjXbFcAU4
3BpdkwhI8vxw1pBHMV1rcmt5zUdwmiXRx55zttWOQGSPsOBoS4e655X/vtqWYLu2ou0HM6AVEDE5
PNciWeEZyq05ZSxLPKOQ/cBEMgzTcKRogWE2ve7zr/bQ/o0C3zRfmdeHpANvd9PqHDHX87VYf/ab
t0V700YahQs3kFiHVPN1jmIQLeux3OVK8tvZpU3d+BT6dMAlm0XoIDUJ410A0SdBRPkS1WHBPliO
91GyVPoDSctlovk2/ivJ13CHaNSEEFr9hsNmxxKpGyg1N5LOnjNBQtrQ/lRQ6NtTGqv2aNqifEK2
0A82SX+vdchS6Dvu5Vaa05lc5ewZcA/79E1XVCKO4IYEzVsgrW06mANpMP7HehFRGcnpwfvmP5Ff
0nyhE+EMEI1ynpwMP6bVspjEiT7ByUdFP4jNG0OE361q38YbPFSCAjtjov0x+IDBL6SRSSwSbDZu
LB7yn4e0654Lx+npb93wS+tuW1ga0WjQ6Kp9C7Qwqye+7gUHup+3ejPGjeNfQN91bFAjrXSFuGjj
1kKc2cvhAhJvla409Fgr+Y/E2rTPVGoC1CPhTPloNNNd3DNva4FH0ny2ZlE/hgcJNG/SsdKfQGJi
56tz9C/rwQJ7lnsTRj0L/Kd1QmRaTkA9cRX26SEoZTNmBBG37USyT7Hel/K6xSpk+o9+QliSqCBS
Ln7JC7gBn4EJCg+3ZyMrzyi7w+QqRHt2dbnXiNA3xrzltkLGi6dZI/mPXCmUNmz/OJ0imaHTQIqW
ogI0kmpkW254j5hyt0KWUwi67PCEAJ+ZeBM0SBKB376mGr6dH8rwFV3Q5iQasIVohg7biCUFW/Mr
zNxSU2NIne9CclKEd/QKAdsTtywm1Zei+gT7r5roziXEJHODMRMPw2fgs1W+cXqz9bFQ49YW8Dni
C9MCM4wtuC1zjxC0/zk9iOXdhHmOGMvCKwpLSEAE1R3V0iSL8sp/mwpkos70XP4tnnKYuUFsCra9
9HTIz3uT7HKdrOZGEOx77Y4aHVofNf2ob/yA0H0sQl2yRfGewi6Z0SxiyhD782ycBYvki90ZRRYV
wcUG9sFgZn1Saa8hO0nTVeFA2X4uIjfomvTUoV8IrmSM4m8x7NW4BzKCBlP91Dt4ClEh8n12rapC
2ltwlVKHXq4KTZOmZobP0QXD7xmarw1YHAgOmffkhhNLRLE9ZjS2uGp1MR2QO8CYt10ET/9a0Den
By6YAJzk31OtrlbuvCHbXf8LjboXhDKbn3AnJtWp/2XVS1ClWv0YwWg+flSULU3BiMbD1xulHqHU
yPTKPBK7ok6NOgpWaTdhT/gv0Lbf6vVGr2QbSeoiJv1j/6AM2XQQ5uKziFE5VaUecb0Okk+MpTiF
iQfMHxxmv/yZQYorNHklIUPINgcKkIl68TfJ9gA2nNyCPjoAds3ssj43st/+WIlFV1bGFMBS6+cE
5D6l2ejtob6xHPRBf7r1GzYQ3bJoA+OIJBACoDjXDgITTBVKvog4ff9lNETO+1nnBhVZQdhnO+Yv
Iu/nCJPMDwD4KVZ+H6jC5+fjn53xIDBsjpxYGYqOEzx4aV2B84H4HXpn+bFzolMAYjA2kLa8hYCp
1eoN22gR6oOt1fCGTDdVusggSsWSzLuLbasH9WxK16kxgdkrlMdJYCFD3k/faYaB2m/Fwu5CgYkO
bUDYC9QZw2T6foh7UeFZ1xoypUYXdvGNisya5/F/haHgzXJcnkg4XRQy9IejSsZX7oNwvWgUCpzi
BXDt67PPxRTMKbizwKXwmEP0mAHfdGXIR669jGbfm6Y5a6Sj+sMV4QSw9yAlKzpzFUZMv163UPtx
sJzo1I0nZELfJU85atP6+S1lJUmqqL3JhiYEH9Tm6M7+OEcIMNULGieNKj3nGDGEjSdUkn0qD9hN
NZGrQ3wJQukzbp2UsGqSPa+6K8b+lgZxsGQEBwzpKj4dCAMGvDWg9aVFLgbwwNLtNL+W3YXVCYFB
7WjyZwLy1JCLaxrqs1DNMW0CcDMjvhlEw8cjEW9whlhcaADbZSbzt+s465juqVtkkTCILHw4dXlm
GnXx5/7B0OIOM6qnJ94XXiZAzto8E0gmTnUtECei/Opx2Jtp73KgaLQumTE4xC9CjOUndm6t+D8T
qMty9HSRFej5315Ajl+lOjWeaHg3YfWQK378wncKwaqQxf9V9SUtlRUcLtVVjyCxzen5qcVrmm5N
abDds3rmRKq+VO2gcLqopaG6PUnVuM+Co1whOSdqg/2jmxJWxE4856L+1tc2v5FDzBSSva7F7e80
QPIWtDwvt/Xhwg2PO20+9ECHpECdjsgg0x16NEKwLKn4TLHWYPUlT7w8jddPZC+OWfUaML5jwn0y
03ER4tDUAMbudRGDqkH13vicXasnchF06fnYsK6MDem/Ci6Ipc89sJENWwfMXzFjbQIvJelpPsRM
1YXPoDfvljHCGKF9hsqSvpnTMGAiK210mwo/DprlhTgAjQ2YpYrfx562QSUpqQ+5w65gYGJso0aQ
2+1L5Oscli3+BYw6DqmPpnUfwUp+p29HTt06xoOIQcL3cq83N8PVAq5yv0Zq2DrQfkD3Sc4pLTzF
75XYjOKNmNsbM/BdKUI+4AetS+w74mnq881sVWuM3TuDkPyp+s6NPmo9M+ij3ZaBQ4N2RxrtHy+/
QVNRop24t2g8OycJg6dbq64sa4IfRNKdwGYcJFufaR/U+1IBps/w4ly2xJjGYLoEAFQM/sogNqsI
RU7Zf6TA0X4UY+yAHt08BSw0huF28wNlZ6y+R31thihNRfPDBOf24gDZvLbKPSLR6B5WLjiKqqy6
wuZRg0k2Bx653NUXdygCgNhqQSkwGKaQiKobMEW4TxOI5X2wjhs2W35VdPv8jwTb3t1rZClmZhfd
W6OojBdTsFtRCLoAB5VlupSSYpBe7ekUXwS2U1nayhK5TWQXbiqRqZyNoM8aJq8iDdU4jZ1gakqe
tOXwvdHo0qU1Cs6iPM6jgMppw2Sxg/Wgokxw2eWqfYEK+d4iSfVuX5/pbCq2bxuhvns/M4YJARgX
Av3UsksKtFeoSFaHRwDcI7iYlGYeeeZJXGTaaEraiKfXxlZuqbAcz3/9g4Ms+5FEUafOeg6XjHY+
w/k0LE9y47iVSdSi2GW+LVanXUBMBvGxk0eNnQLhL71AKV0ZhuzuhgMKl9stBVU4EFPNxoVDjSFs
hLTTc+Mdpqezsf+QyyXTEMCrxEQJIQMBI3v0cLg4Q5Kc8eqVn+nefpZs2OXfJvEdPpaGczf1Bwcc
akf3Gtf7JkczTsUeUQ35tTwZmP4jFDkuB8XMVzfvPC0aMxRkm9K5oK5UezFPzEmXwjZEfK8O/4/M
cAM1k3C2jhIdG+hQrCElv/D+srYUyehxUzQ5I8IcGDMCkPDw8+N1qbSLLlS7OMdxsHLKbSN4vjL5
g3udtyjzedrm8oR7eov+NlAVzvNbidgaJ8ngXUFI/4kSMBiQdeSxP9dZ4Xw/tsPPfQPSNxNr7Kxs
QTWV2Vb/+gfT/Jb0y6QilfKfjjZD94zZhzk8wUqq6h58uMOhO4ul0bvuKSvvyeT5UzZSYnAkfO8u
F8iBIDmKVXUVGfCiZ8DlAug3trwgmSNgxop7gfA7UNUhjp+3LgRbOgxJ0LC3RBPLDh1GVl+l4qdJ
e0Oij+6xLuoIl67gs8E92o2+5YapLD4mGZ3hduooKerUkPU6b01LjwcWsaElltIb/k2JCzL1neCj
Dfzr5EvMr8ZbvWSAapHnkVV4Vqmy1MN9HUPFOc7w/ygKKrq1SEGb4urhwFCdFAdSTElnyVGtVF9e
vQ3dIP+BvS19nU7UEAo6ANRwxbtHQcwrABVisruGsh6P6IVU1fXvXXhZlQ7p6V8WF2HVoPURTEUj
XJmW7xcdHZzBxj6ZRuygqOO3QhC3NEJ+rhkG4OTeBixfNwQbcELJeRnFNVALM5E3v/7XnkS5D0TE
Gbq4TkA1EMz9K0MmSVDX4rv0hjyFhkWKRTIq3f8kNrWupWOBgWEMyswhf8xRh52qRs9OT42jpM5S
uDGOjtky6UNzGGIZp4yf9WYN8jD/mKsGJ7B6qs43Z+vOA1J/LZHGQB9Dm+KoiaB1tTyH5en8z9Z9
swrzHGmhyV4+KazpjnwOay+jQtqvgcgB5mAU04qtiUykNm+7hn2wS9npy8t9ofpOSebfPAT0RjzJ
YpZgPuDbDRAiW2yNXrvLAu1T2LYR54RWI8z9akj6Hr3KRNJ1TBvarprdR/khZ+q13A+XJ/ebAW0h
nPTbQq1FGVOgKt6kqUXRMpq7uZ3vHAXeqTfptBctdschqVLcM/oKlppHPmeRVZpoaw/zT9E6vBCJ
w+RtRDPvhFifZZNqgFjR/jHyXnr/KFDqHDt/A+nNMRIQCv8SrVXHtVGGBMwt/4fcFl15izw6XzPX
n9nTX3qrKE6wEzZ52/khFZqZA1Vg7GL2XItcyEd8DSbrE+yznPOL3tkkAsSo6ZcEgJnOMvod+WIU
2DK42DX2F38j9cFtzjB31VIMmqhfBoJQpYK6Nku6+ptKohnpkFrjB0lUbkTSxwEzzd9T4+7Pjz4o
AvViKX691QAnO1S3QOdhenQsOWKNE+6gXsdkiARn+4BnichhQref9lvgLEtp2gO4H3bdqF4MEhkP
yxZsQHi9TPXG6XKOIvbznEJdQq25lxMVErWasgCDRFaQj+jfPmZEl+NaKubSjq5maZ5mSubEpNLS
2r/T0zwhpbjLrALWmNRpDk1R3PYQgVRDRf7xxBkejPtYE1UOiOusQlNNbwNbhhoMucOF1xTf4sVT
X7zb7504RgxZ5mrynkBNO+n3t8Dh2V5FAf/u7cN6T3RqJnIBMXhlxnKixoywM4YBHhas/7cZACpZ
njmXwibdqX/fO1E9xszH3Ep9gGKgh0pc19Vov4tzaMyeYCeeTQeXa6LNmVRlUvdLnbIs06H0yTvC
X60M/sHDA66cdPRwZdDs5R7XSNaY7NxLwYXgg5TIAe58FtHrCwC4HyXmfVRPD5RBTl7BHSUv/VB1
fZkLCljAenA3AxSTL22Nx2Elkhi1Xqd2/8DIzmOXWPOs7yrNUwfP1fukGas2Y9DlbU0SIa6G5guu
yGCeyYex8bm1B4HbZeglzFrg2TzFhHMW1tVMrVFnmE2JKJTJCvHkgDU0KRN3cx9f7iFGApIopvjo
4lkmjKiOjdBkbWfpKSuBLIncWSeHIHFsLLxFdDy+dJdxzPeZ7TK+2xzIdmL5V+Givkpg7XVKOl98
vDAZvikoq6AtowXH/vI7x7Bpqw4U7uvozaM2lpNhC7Wu22Lgzp8akaWmuvX8rgVNI1w49q9X7cwb
MbEoKGaOLAvvMpZrTA9sZzTMok/mBmQgECU3QyGAhJbTaeuNr/RnfqZVN2Knmba7MsXObWYycvHB
J779Pq6a6mVJIOldVkCPaRH9CJ8y0SwRiTOExLPvrJK/3O4go3ZzZYcmbI6BiVgCQJtET/QGq0AP
tOgJoInDxQcyUe/fHWcJ5xZCogUvYlTzQ476JObNJUBaMuhYZn5HxvOt+AQXtf6GiiMRxq8HBX40
rtCW8zQ3uUG4Ilk+zkhMgnURU81K6nammWn0Ai4wAFu9Y1fuMtSXeSh3+4GBmN4MVeBw4EL8hHcY
Sa1SyrkjurbeupFK4nFhvAEGxIQnhHkViN6w+dYyvB8kcy+NY0F27VP8dB26nTAbnRJ53nAMh/vG
frEQQq2dRTz5dkVptVfi9NWG1E0+8pl6I5zHF/CZ538Jh/1395pBfUVOOyx/dQ1oIdSq0suBTUqX
vFBq+bETdNvMri0tMqR2ibu16D+3dLeoqzkqwsQMTgwHm8t90iGpz7aA1+RrNq6vaSHyCewxt4uf
hBUZdFiul/3AVWqdN0f7N8MQ61b13jnvPh0GfGm4WP5/fZnmsRuZvoIvJHt70q78iqa3u0gciXHh
vbCfZFrn5fwafXqpwF90ERFzoQyYoPFP4sy0dzE0gORGlMYP1uKhKpRogfdFh/IkPOtRg+dEOz64
LL9nNolv6iPdTivNfhOabUolR0pCVyO6PB+PCgdlkwZorscd6af+o008kE2wVP0AHMIfgeEtHi1N
9QO2YN2wb7OHKACAUL3t2WdWhuvhsj31WwMCd+EahlMlda8PlkyGrWUIwEet4VmfDCrDbhfyXy9i
n+wMQy80I0hgLlKuZiTo8j7Y9indm38iPf2pmmN58i6djm+loPmYkI9MHK4z8OeyGQRXT5yr50rX
Jt+0SoBb84BBe73bEXkPrsMnt+076hHNoBPVr5HMR5itiZEhEeSzQRgp8rWowyfSon9DVjYxR6rb
5Umk8WzTIq8QCagO50MUhGS9dl+gJ30Y1Scdm9OstZi7rhyw9jcVFjhS7Xocb1XyduayS4N7Tmgh
mIusFEHNDg3pM+wA+6nuNX+mOa80lVQliM2crzkJIZ1qLfjUDS3B0HgTLSIiTqYcLTF7P7yJx8+9
8Je5fIZCB5dzwuzn18fV8X52C0tIm8QjxHajtCGRCS/pyLJd8NqrvXzuY33kvXQZPtRm5JlOEfsT
p08ww3BUlTF78IvdmECi6JPj4AY1OH1Up2asbmlnk8rzzFCom7civu7vYKVRoLiUuHJKql+itTpD
9MhSENpoOnt6nxQLQbjAC84Z1eXhEt9pLkLwL/M1FGVM5C6Q2jm/n1cy6Pkyvb9eqsxJm55oMExi
Khq3VnOkKVpY5anvfPlTOCSu3wzZvB+Zq8udsacHzUYC83su/mQDy9qjAq8iyU5Ykas5BYgFgBJ1
ixaQA7aMt+PA+cxoq2aJK8AQrOaFqqqyTC8NMtAcjHrd4bEC1F6ZgSq0LAh8SEZAjRQy68FGVY4n
R+yWrOPcS8gMY7wD+ehQTm2hJ2sHxjh5hQEs/lUrdQTpwjFhYMu3xj/dVHboxvIHNMY1c+4G2TfE
HHqIs6d1mbsTB4fyVdYVC61VMR7crW4sAzdWot/7Sr0tyIPTlc+X9Uc+OMGkKNWD1uHhNQnhQUnX
4HSL5HUHNEH5GJC/csXguPjmNU8TOpiLZOclFoZgR3oSJRdYZizelRIvRO1CoY4Q30rZ1U203Jne
dNcALzumRCTc3rQsgGLeDrFnPAXvxFX+wEL2eo3tzO94Gd0QU6rNEU2kcTD8iXHnJ7neKlGd0mri
93CPApAp+03RMjMPNG5/l2AztE7j+1d8APnKFVmjbeIFqdI8RXKT2eHcazNjDYG8zjZdb/ZCP0ce
2Mb6TeLmrBBx/KAkToXblMQwgNuMhhYpu5DlRLk99pOOXjsARje2PHn5GcSxK9HEwoYIVWWpaxTU
ub0Y9N37fQ/OVOumOqhv2NnkW1N8kl/bMyooGf14A8Ckpk0NqHvb3Q+LP+g+mP0qxRBWYhoFKkL0
jwBNWuKZKGYkapaK4ccsCScGBaf+KFIC9vOy0B6J2aWS6pD1/rGb4zZA+zow33/+fsgN0D2FWgKQ
MkTBdoylnfiiRD2VPPSLYIfMZI3zYtaxj7sY1mtBaWq2mSPUIyS+z7p0ClpksDbYfNcjidvf9S/b
WsuQdnmoDptZhjMMGRcBHRcsbw8JOgNbQCSqTze540yba/otpwCjEzG4i+wAxsX4KriPCTuxz+02
M0ox3YF2WHm6M57fR9Q0+bOoby0qRvVmztQvfy/jIRspYlf8eSMDtyPnwpFJtoQ33INjALb4xfPB
/sMm11YiauvLlUzv8sNgAJ+bP3CY7OZBypOsNHh4xYnk7oJU/vbNa4/NCyjAlCH3Y++AStG81/4o
iNSJaJYhCBBrcrqufDGZ60owNAIezASo9rcuxL3p5i54U99qsr+bEdqjqx0lTs4PI/urCLdoKvzM
NppyfcycNLRaKiJeJa/0a9eaaZR5mcD+v49MxoNU8veDKBlYuRBa8Gkra4C4rscgDGdoC7ndmoZK
dmy+uaAK4uCACvt57vo4uziMnGvPisbk4DQgPPAdzz+pEbhQ+So+oP7X7cSENlB+pQkxrmfaEW7j
6MCg5VYlQjd82S+guvB1Q1OZeuESWr2T8mv0V9VI6Wmo6KkZa//WCpr2xTlGhrR2CvVq373pH12N
TqrdFhvRWubPY+6oXeJmgOmVOXoCSXl+NVlFDPEXdE2zIDwwrIWRZlL/uDQM+AMONWUUMtz98MM2
f/Jrqn3+FGBokJ7Z5puMsdmCR7AnOY5mCjjbM0Ks/OHmjzVhx/N0f+grM1kWE7isdXz/pElhF28U
v+99W6Q7CC5Aua0TcoL3JAxD/Jc2wxwpIrrQifhZsY8JrlJ434PaqRCU6Y34OP5BA+uxSWLM6Q9n
Eh3QDl5g9RO+3T3E16wYEoNgalO/LYitA3jKrqn+TXmt9Nb4P0I7PDjaTadYLwe9EKtl/ceXXE95
5lxRo2DLLmevid6alXm29FUaX+WDvWkMfAdy49zElQcXV3PkqV/IzFDfFj1ynK6kzRikwCDIjxyQ
oQ8nk9eDJ4a3txB0V2H3xKzoSxePtOFIhk35h693FP07gY4rCFkLT9PpcnizrwNOQRLuxUsmNgbn
m3SOU6Prje2Wfz/Uma/Y/uWDKnKvHP+yUWFWefNg+4ztr5l3seFVnvceSxwyubFM6THpR/Bo94dF
fxMvP8x2PZZuq0JvtNJY7goWH0zfoyEzuiFX1dhhwt9fuPbRXDwpIzMrU0tgd5o3zwgOAjmVVi3E
Tn1d6fdshom0eyOdyY6u6LmuPeBVTeNXNsUGHZM34dsSzWMhAsm69rN4SEaiJ0nMPzqZFUouVVLH
WaEAqwq+7G9DQ7wDWigcUiKx/sjAe9T7gzOBmwXh+xIB2aBUY7AJB3iGlLiSItJyrkkqTKuwBFFe
fnDJKQi3vsK34/dKOql2uxuTQE/rI/tI2Z+CuFDDiV2Z3XvMi8u/vI2UNPkDmhr/uMH19xUQtfWt
tFT8a+F5Hb3AhWSCbwgYVKwrigvEnFAptC9uNNEwf74kXvBVPVi24KzZBgrx76+ARXZ75FKHeQyh
ob9cbe9xJ+0hPbX0Qp3ao+DTfSOsk5i7EYr+OjptdFRfSJV7QPrMe4aDiv1KRmxfbNLZf5JuP1M2
e6n6QusnBQWn9jjUcFbvms508nkOwNYscOWR14Q9nb6cJgRbESCoEzvCYWji/wAoluY1pZIP6eDw
9icrGFsxyrmcobAGicvGu+ZAEPfl4w+qsSuZVEuOed9AJ4OBwfYji2GSpXA5MPIEWKjb65RzZRlj
bucQKzcn5JTkI1kMd42xcujQLwcb6vCpt8hRVz/vUvs16USfBVciHBxFAZZOWbxQQXWij3T9FHty
yWUX9fJlYdlv7lBKnkbjx1u66qvRsuRHUhnFUCgYqtBH3E49ECAvwK5pVzAYBIigSzjRPBAbsqQZ
yOMbx2YynF8+w6m+PTnibulKpdQRSGmFdGZQ6Fg0V5B9/kvm7adgMNn/AayctpoCwnuMDS+/jG9c
cmnfEC5l+yFLfhhUeQR7W7O4IXRbsen/cdHdaS/KbqlfiwqWUvIvluRzsDvbbobWLqQZXYMKzBhh
JANqlylJB5YV/w5iFeclGUjiK3SFw6WbxXiJrxwBXJl78Si2Ba8BeavuSPD+h1TDNIr/D7mIsUQI
takYN2SlE97WvDK99PRfeyunEjRlXoDISGN9tLWbwMkK+yrDQndhEVYxfGvv46XlaGevnC/x/b/w
uHe7bDqqvWDTlh04FeSdr4srQUJWI4f+YmMT2I0QrYjkV6SckbN8q54yoGsmrJmem/PEcDlWkmgr
OaR1Y0kQ/jtEwO6as+mJFHsyLE1e82Zdatj16CeieDP5cLplHKpRu7qfd7TsikC4F0jcpsYnTeHm
68cEX0CY3fA0r+D2a6B3OMzF8yF43db6C5c4GddXKTmZDC+610MjUSndc24dK8bq2EWWdhWXLTEq
XkXNobnvLrYX/BwQ+GCQnl4Ictmt2PrghB4LAUPf2e4uwDMGEGhYH3RMhWVoie/wB6e+vAlzst/5
lcYdHuri/97upYj+a+yI37GYcQI+QM5F4X+kFRB9TnQI2/0YkepadvP7LRBpVumFmle+o5fq6y7S
CWcDeX5P7wdgApIHLnMo3KcLSM90CuPQpscJithwZc+PDGK8BgcXdzfSpX8Kx+RM2aB7lOobkGCZ
mRn7t6gRNWTcAol80FsaRArwhNzHmvbqHQLRPbqKRsZnrxlRplrYeuXKOxHqY/tOcWyv6AZKdCSs
ze3PHdqXTPbsVbH67Xy8/SlvNnxNlbXdA8mxhHC/KM+m9eM5rkD5piA3wv5zPGAMyFVJMeij1XUi
XeYClJthG1Va7Cb1Cpn7Hv9imqLAym3tvgvooDQ2mwW0JrJLD8grJPIqcLh0rbxepHVcIVu5x93s
9enqBvbbvtZ9lGbA1VJ/7O6JuLJihqWJ02OTwVCCXo1xThSjxTaA9CgR7kF3zwI/dmqzd2fjmoZ0
BnR5vePUmWVkqc8AmfnbxnqnjPtZJQ6NA1jrn1Pz1lwmXUsVhSSRLugPqvueI334JDbVN76hk9W0
nDOt/r4f6k3kHqjf4SK8WYe0jCGJ5ZWY05jW0fH0cJVfvtLsmYzaWC+9puG/qUKsJv1EEj1P9sky
M2D0Iwxpv159SQdMlJaqNxn/0p8+zfhI0hTthnbyJnaKqiWi72PW+uwIEken72fihIA3xvfL+CZw
2AU3NQpg1DT0TdAqoBCGTh1j+z+9E2GiWFAmWTbGh+wA5q1M83p4yQUla9G82iDvOgKYiWoibm7p
YqvyCTRZROp5ELANtE+uLTOlmj4cYTksbH0lnlF618NrCuiTVKSLfGKmyPGC+/RgeDqL1qDymNzn
Y2n6d3USKAUyCMbz6ozKRzFM6Tb0EMrG8KSDpC48g/2hqLsUgNJgExJmwJG0Vcs6PjN24A4M8Ni3
bGm8el2A+MXVDx731pVVW6S7/OuDrqg2vmHon7ZysrkdyMrUTyOh8JvSNM4mFCPtu98jGdj9xV91
CEjwKfeqWBt/7crI0sZdmgEIrjjcz0B6WFNM1IKZTcsOjrBqjoIMw316TdyZaqPf5bg2tmmFllnR
eVU4kbtwZJVwXyCmiNuoRve/ANHSBD9CClQYUhx284BkT7ee7iCs6vjBY3j9WVJa2EfP5LixaCDo
oU1j+DijxJ/REsLB9Zxtie++zCbUDqX2SW7GS4RvUu6VI8/LgHNV4DERlI5Asq/fJQ5Yo8UWbt1V
4SvPywqHcsAFDeFU9SQ1QJGJbfDRMn6N7iZwZCym6uZJ5eOM6Bvq2020I+Cx8orkiFWbY4sB/m+Z
W8aJn0VwyvnGP4dKyWlzeL0PnzUL9fj0UlWTUsWF+jNrGoev0UKrj1EtZre60zqeZJgn86ToVDPR
LLhScYbxA4jhpiCoewcSqiRVnH0sCXlwwwF9uX8/smL3VE3OUuk63gZfmgJJG6pwzm8gIIYo7Dgd
3eWBMmZJOO0tjw2fqsxnrX7rDdZGtRzIgXyjzHIOm+608ALBec7bWHOt+lKM3Y5/wEb7eHObYfJS
m5yr/wh24ixPefG4UzHCfi5V+HkFjRgvol9Eku8E2qzPtbtcfz1GhlrZZYqLdd3N6RXRS0xxahTn
0u2CEos1ywUonYMsFpTDd5qxVMN7rOT/NRERPUKVorukzMxTC26M1lQLkuBy/4/YLKPjByy4YJiI
7OPOxd6LB3YPwGLQVbkFNit3KZx1IcjQ0jLg/dPll72/x0CzOxe/qyp+reBclvZkH1bsTprf6ZtZ
cqOWMtp95EkReT0VOGhYTaNDKi0HSUj2Wr4gdyEeR93m4BEWVxXSeWdJ+TtTN3CwiOu/+0rePP4B
y4YiJn0N6AevaJ9ywJ59pvq/YlQqhdTQ7A1joqAwzYFxP2NH/bH9/PgJ9b4M70zMh3xN3nJmXykX
dn6HlaE2r0CzOM2UNqkuYIBS2+UJxAt4xqLm2K169MnbVG3A0apwiAcSG0Qwb0NKBnr0YOmfZ++G
n+Uofnok0sdoP/oGRKO8Eo9suH6tFPFPif8mgCSGs+p7LYMD0Ona4YclRxrI2rDc4OQpLL/1ENFX
fdRKlI1XYwrNiADSP1LU1rpTuzIyBCHOSxvsSVmYtqRfHOfuiSmeK5fFKmZDx52B6b1SOA+AYOkE
fP0OuiA2QULhqxDYrj4wHCClkvSYB3KVLdcDuKPn12vn6MLNDM+khiitbcxtjr6h2aPfZx3aOGgX
zdH/BtKk6OMGOlgghfTrAk/2bJmJWuQ/FS1v2DWTvpUgpRX2gPi4aZTO6CXKTJrEvk4t/X6BYH6n
CRLTsHAAcIS/rhW8DU2RruMqMZgdLgL2EZMAbiAqpTf0A+GXQ+DiLkBM9EiSs7G8kD//Yjzs4r0K
vXLXkDxznCtqcNfoNlAQnl+4M+FO7s2V5dDXrKAWU43LrbGxR8OTszllyN0UHOrqWrk5fM0WDLNi
KZFfVOJNc1dm4zN3LThSTHq2GJ9VlWzuYyvTpIemriXWgX5fn2v/PZnGyHv12W120fBKYv7je/dG
yX6LMjNd8KbLm5sbEh7nwWwfRgj7rL4jfi+AfdgREswdkXwLAeD8KByiMHtIINFwWSaf9tDJQsWh
iAWAkmpe23bqaI+sBBEJc7NhDaMWfElbc5xFZ/dOlr6Gad3DboCM/xiPW1Q2ePSCDMWqx9PoQg+F
pBlHHXx6eQM0h1+Cm3ttJrBqx8dOBEX1BU3R1g1DViP1vAS2SgASjz3KhxOcMM7Z4PS2dt/o6g8f
rUswJRNVi8mIy2ogv3nxx8mgnaBoE6DypXPJ2Of0F6QTwBoQoYOA83UrXwaESOfgd4N8lfthuY3u
TflfkeoscoeHGHl4xiFkDnnSXTG+qiHqUD5GSLZO2UrDbrmhbzEmhbhgxeAP4UsDDsaHe9tICUy3
eJY4Gji0RtIPVKqmwPKeFW4G70DwprYmGtbXvofFsYnuZO/j4D4e4oVLgSC/aQcpZeFNlV09JzEd
9tb5dF7d8cOPUqVtYLk2mt9nC0lMdciCrhZ3rh/oGl5aWptyVcBzFU850FNHj/4odbRy5GwmMGQ9
94flcXHbgU3J7W83dKgLEmcxYtCekjPRfz71l741G/gE7sF69Ya+yk/QLXU4nrvmqkYSiZbSPtZi
+kK/zFDERXvO8QsQ087tMN7E+EUaLaynIPqaMa3BnPsvnjGT5kBCe7Ejw+0q5EkTddvKKsSvtPKS
mOs4rvqyKyg9bl/nvQBFU0jgNUWOxiy7tHyPFjxmC+yRU7dfyz9Y2kHawdCLfDTby9XkdLoAoLL/
UqRkarfZkfoexYfFxBaHOcPaclsbMFJvtYUzBCv+EvyiyvT8tfC+Fk0rzVzPUuFrTcdTTzsgY6mC
OMFB5RXPI7zy0OptA5dlPiW9WQez0OlRbPlrYaoBBtibZTgQLdQCv05p+z/xEFzrNT/51AZJroAw
BOSFTZzl+1hJi50RhXyGmdNXHzRmm1StDKQoBmLxUycOm1cC4BZIXlAMKGnMCKmzjQvlds1NBheV
SH0ypct4Mrhik9ZMNqGCqWDHwqjE6citVNOnkqCNLASYI/r7BLo0tBGt1BJSxeFzQGl7pY9CbQI7
h9cTvaPcyRk439ULX6aX2hNha8n01u2AoMbO8FiUzsCLbApc3xB7JaeZW74bmweHBiX0VMM/eUbr
K6/+C/WbOqZ9ubLWAAiTn5ltIbd9hWcLTG6UygScfoqZRgAckHblpMuwkn0ce2nZTTqFLmYbPMIR
5DKKz794oiWXvQuExchdMl/Bv1E6/BriRqY1OK4aSjerbzkGaUtPLrqJ5rX6LXwNiCoBpFSfc4JU
h/EsucqrwXMniScq7gGP9nUt2DIOS9SIh+er5E+hIlmWZZBZSZGRhAuo3P3IRn+dJciiPIOlnq7x
EbJNe5lt4c7oYGYi4DiRXyReAYQd8Q1coC66h+bEiuGZXPqAYQzLtOgUPdNRlAze1Tl57UHTfSHJ
w3s6aCOhq+fOweCSFJdsoLaPSouK0/u7q1/sS36CHMgf3czIp9htTo6LrAwcN6WCSFtLWA2+VPfv
Bm9CZdDFg8+00YFWbNR0gFKUgbbTEI20LDesNWkgjW1I1g+6SOjM2Hf4dTTEinXaC6xQxrm0YSql
EWUTIhyOg5VNjJqQWJU+YMop2L03q3fNlEhowweGG1FpWU5yxuUjmyfaTquuPKz8pxzUVFc7h3aM
Jjp8d+ccS9oRErrka8VIMhg81AuRoZ0nqcEcyYkXHood4xZoVcrNwFJhmKFmd5+EdH5mjILGvqlZ
ecHkKte829KAZxabA2dAORhJSUqS6DGwPG2jo4nWM/HX1k1I9+yeKLt2ZMwmklwyJ8y422emqodR
K5Sz6EkFua6W+6MuwxdwV9mVlYFQ10RnFGRjDQ1af9du9b782bh4vgcPD90r5oh1euxXtlL4HZbx
j2yBpIcgQdgveBUVnbzq3HeMW4jHqeutJOX2RDJJKwt70qu5lOJX+pZ6nxVyvlCHt3cuncFZYwUU
jBBINdAJw4dKyPiOOhoEY+91d5hoGc/3BPAFRuz11NXmNXk/JE5lKXYGamYh8/DatVRZkrYe+7w/
6hzXGgRW3ckz4QS+EVOI9gK8sY2I73HhwWOn9Y5V/jDfjfLoD7fuVift6jErEy3uhyP0krtYeopn
gtvwQTbwfLDjh+bMIbKM+PRe3xC/blaWB4hLSx01xUnENryKb5sfcBjZTWI4vumihBEFG3rMeXLm
inyxQGrgjQAQhDAt7d8va1SGMdAo719EyhJ0oIP77dQyNFjYPZW+FoV9Syq68h5HzDox21Ry3ZFs
UARrtRlsUR4QnnekigYdeXC8GlwaUFJ2nJFiaI34p61uvOLw/SqLZp7nI52E74BrfoUJomNuCddP
eKUPHIAAMs1zz+Aipq2lW9ofU5UZJB279cIrijnYv0LUDATvq6VB3BCKlshKZ5Av0KL18nJZTH3o
vx1wXf213PgN0qZhjgZ9paLUxlx2gpNBH40lgIS14zXYF7e8F8iIY3xZP8aOAMD0asjSObcqJl5h
yRm1anohlLwVdbIOgTJKwg5UrKeZIyKh08P71KX9kMGi75LBGLc0VUpvkQ4gq2pzSJHTFeZEyhLt
cJ8y/88ryE3USMlgwum50dcC4Ok4Jg1oQZMJFabEtos49nvtLIRPfc/Bwb8H80NeHCkAuoQtqgZR
kvo41l1y7pmS4//BaR0DX46jF/92Jjsk/9iLagytv2rSDbSXNxp2NHcF/F0BhD4Z6LQ+Vn2RYl9J
N3+okp8z7daziQfCMoBKWeooW0lAtWyMbFCxCeMM5E8gPQ75Ac/1+rcUSncLfKBStlmq6jIhOPog
FoxuhOmKOQXNU45NzjcBrsLw/UQPZ9TDGe8tWpc2+s27NT8vk/Cv0AsL6drZUEPhmLUWeGm7FC8f
s+2HBTDQJnKbxSUz6uUD6F8HPqihnTl/aoor5FYIrXyGz0N8sCT62l66TffOVUIIQJY52ZmDQLRl
MuGndiDVtIDYuOUO0PcgF59uCMPDJ3usDQAO/9f2VnTLsGo4l7YGrv5qyU7nacYWt6BAFHt2He83
5zqZBdCYbD8ervNzy4dx+DwSvYUhaqK9oNonxLJ7Oz0ktreAvyFHdED8ksC8FkQfoS2WngHztCFa
06YjF0iH2Puj7V9sKHQ3FDcsCMstCnz2qQ+VScb0VWfr8WyvN3DvpGcAiZ2DDH9YOzudQkEdT2Ym
GceEeUYzLrBBf5nxLEXfYerXCK4PylsEfdmtOxqbtGCuJntk04Q3vw3eP/atz+kJDWNQKGFREFlH
SZUZKczqnpqn8VmvKPT+jRSi3DKcr2ozH1jUGaVHV44aUkYW24JMjQYtzwKwF4bFee7PluOOuUuM
QyfhrUdUHXzZefn1xRyCZtc6sef0VL8MjVXOnZubJ2G1kYNu56AaghCcQoYYrA1FwZUGidbBZTOz
b9shShpGJl1WAZPXg9fGrTzHRRtdbQ2UPGziAZ+ddUXE8l5+i3fsbe16pADoIwZCCE+/it6VTpW9
BSoNBxw5FPxnehxSET+YMUD0y36iZKU40eM5em4Kdyi6jvUJCKv40IqA92nGC6EbIb3Kv6T7ycbO
MGu74p4XNCFhjuapQbdcE/JDmUpI1LKPpvZNIb/N8cMK77yq1bbeybvEDA3B1SBwBsKzFkRScH7Z
RXGdhYl8Tx/QPH3KWj/8cP9NELdXEiv4r2QWSEV4JjopAFMvA5yetYVBW7MRdpX8jFRMtqlljiLM
NvaXJ2TcPx81HUZqE31M4F4SRB8d0g0cG3MDA//g3Dm/a6QAmCfhQPwAbEacGBLzb/P9taaetsZU
lknT3x7RAHhNJAQ+jXVhe8N1pLr2Rvv02G975YKGrnouLg/C6O2k0ys/PZ6/vwqO3tb4PxiaKIuO
E7NLZu5Qok1srE+bg1y9uTaR8VopS2Hh1+L3rPBKt9Vcdg6HJVo04izqre6FcjJx+F8xWAEko7zT
/Cqkk4VqH3KvHZg5b9iNb3laUZNbTFSPPs8XCxs499Tp5o4yDz+TXaJlm3Q0fLx6I/55H5bSFiQs
0pvhFl9yn5SXPKXeWxhzSqAG7Z8Ct90A3ngb78N9wqt9ZCG1UB6rMaUXSQ/O2SpKthhRVhwinqzT
D/nw0ndei+IFaXr45GlbK/ZxPmfuqwPG7anw/ckhSRQb0lmxaEchwbDxI7Zv3ibf9ASbEkuQKuhC
h/aYvKPwZZqF2Wm7oTy4RC2lPzPpgI8fBO4ja/pyhXpLx5rqVnEV88FwMK4tnAyUkD+7rXrcT/SF
Vk+GQc3hbTWRVVvgcYtIRWIsYLNxZ/Yt9hUPoXcx29UVbinzZP4TEWihz9LKMIyBMA5UNCsJFeBN
nNWOjqMKhCzw9NTmMTrCCMBWOEoowEOLwSlAlFXtQRc1QsgyZGQoO2BefsjWJyR/g9kgXdzJIhYN
mIdc6wx+Jfm+7me8H5syDmX+3DNYaVB2YIypNNl1HDspFwzMY8yOa221otyL68SzVyKHSAemABtA
jVDHFKoRDBdd8A1KTE+UipvprfNiaZ8xFbFJ2XytfxvAVlKybcYHUiCZSe6Zk8fJfWHPforW6sTL
9Va6Jf3DiMXKAj3U9ReEzUvqBYXSqm/rOwMmpjEoDmJ6kOoUYZkxggBuCkBjuhVtyBrTCn/WXgo3
viuut1uRAgD26rrZ5C1clYWawzSt8r6Fnk2YhxbG3RsXaomsa2w6RPG8hP81afQsvHt5NwmwZPg2
19TrXliJ12sRjuaAo0wKfzGhK5B4Af1IIHLJmcBxigW7+AlYkrOMXXbHhypnb5r+l1QlhdOtH1kg
+C47ilLOtgO5JX63WMqt3vmV/Fm5h/3JpuLHrms7Fss0pN4CqbThpC0DKhoxbZMbjHzRGMXRmWci
T+Jb6LdmNjIvyvB50iL6xewpHOruHEXAMufEGat7/IVDFjt4o8EcQefNlEL2M5xYUJ9Yt0r8Rm+H
8gu0ytGVYqaUybZhref8MfMPK3PpwEgCPrgAqimxnMVBSQ705VPZ/Hw+pseNZ9X7TWPs96QTrBzC
WGPlvgnXt7pioalpiszbP8Qc+gnbihkCPL6WnDwgF6h32QOmqoU86P54XH15ss3Q9628w4uiF7N7
SNJHdj/SyRFhhrMzOJKur5kw9lVEwr21bWXpgPrOLQvYBl7SuHOJcvvRhGw40Z6HKPpRjbKshW83
zrIT2M9zkSZa9DbcnfxgoPVhwWTry8ki8B5xuRRPqN9AMRX9Rl0qfsLDy5t9ktRE0D3BthZl3mJM
pqRdo/yU97TP0KTag+kil6anH1SB1iKW0bzkubEjsYRYTULTEM7t5DdA1OkA3iyiNHZvl2zMc7O7
StnTjxubAhSvmLqGelviukQzWFybeHuXWVbEVZFSIcTsRtmZHjpbUzzQQiv1lPrqRLCrlq1odxdC
hB4o+tc3gZ9AIiAp5TZIJ0Oh290sGyyRS6UQVPWhwd1Q60x+nrlBb1R8FsayNN/UNld36I6x42sr
cCOU9zGSYMUy/I4npM4qqZe/6iTVepmBNdyUHhZx6EImeys2ZAvYYUTLodXhwC0SqktUzP1JDz3w
5F4MX1Fx0CX7nUMgbFTYK2+JtVity8IDtPjBW2Qxeo1lOcDUxtN6uulFKBatPrIAs6oC22Ul/qmf
fJeCBZ6VYKZMcA6F+80zEJ2cxyXKxSZFLXah/pRZJ0jJkjRJcz4qvBQ/oMHg/kkwtv+qrnl+KOLC
dr3UFgrLJsf6I+EJgFdv9Sv3D/lZ/4eksOszcSZkcu2TLU8GyHbFmDk2ARphFReOoBfl7BDq39+t
Ypa47eE4gFgLFNFSqaJMzT/gFcICGRp10gzQYlqWw1ZC1j+cJGHA27yv60TavVUk50n1FSMFKNEG
1BZ++zgJ1m4z/FBNjuD+A/XakQN9d4dklBA2D9W0byDA8B2fH62LJVWgQqf7xJ1g6lee7XNjzg97
PqCS2nwUjyyiJ/SkJl3JynX/dHc4d1sBxzlvqP3jXHMkqcgZvw7RyKnzcFWAzlTD3eobFcpYKJFI
ZN6B9O/8iLPFjJgkR85RN4ltwnDZRQlhHkYCpI9VAVbg+X3A2L7mK2DN50SOmyi9CHkE9saYJuoH
cxyOid+VYdFczLUBCKsGHRNmHfftKgwHiJoKZPzlHFeqRCQU3e5YDu9AoiIdFVAzV/NVMHZeiAcE
QB4APJP1fOENlnXZDNRx44HJPTl/BjZIbyKRPTI0m6D1ezLdfOy8gvV0RLcC4IHuQRlJa7YHsJb4
yFug5TICih3cjliflcs6m0YXCagYKGx0mVE9f1/zfXIsE+ry/MHwR+Djtinmqp7yVOApmug8IbrJ
uO+1WpV0U6hSnbBXwLWB9UC5spo8CCa+oNq7+JlNuAV9lnrde8lgBiUm/Gu8EpNPbNIK+AxUTGEh
mHGB38FUPS0pgfkkEEyvKCOjyS+fDlYajg+EzWSKYaw+XhDEzx3vYkm5xoq8D862rKeAAYentem8
KBVUCy3Xqh8sDP7zUYbfisKPsd/aB5V9cpjY9ALUPq7u3PWOMYGbVXZCe7CNh1bSBjP7k8/Y1WJb
RUF1lRAzusJOUe/W6LppOzqJJ+DIK7cLT/wvH9/ShwOoYNo4eBq+ExnkaKurA0zuewkkx3r/VBa7
sM5fO5gBncoyfrjeuLvrNCwmD4a3SGk3fciGKUxKgMH/sLIBECf3ufD/Ubid+M+uOA0XG5IBp8PZ
U8tv1vtnFXbDgsWtzNlM1cfnMxXfWJST+3I0LoCw8R+YyH0bK9XiaRUsxfa48V4F2G+P025LADEC
O9j7I8yv8FEkSEW5SxtlFF4kKTpci+DQA97+sQhwu4wuwE6k0kAtrL1rzkU/S4e96g2GDdnqN5jZ
Sm8/rwtuIl1UGgtCQqTAXWptZgXK7s6rfHJ19RPjVB8AHBpo9qFsaswewnjh2PNvLp33MAGEwOc9
5JxJq8YHLt1utNfGB0yLvDIXgHQ4QvH4hklp9l5dXU0JmH5/Xc7wK97R6b5ao/4DAAzF7FAPsrtZ
P219+yMiUIS1MkU46K8FDd/8WQUG/Iz39CpL0qZy4YybU1VZbCY63W5Fygz98wYatY18inci9aSF
4TMr6OPbixjBhL+l9eDE2AHbd3/Ead66zH28d6hMJUxwpGv3+68R4V4sIsA3IR63CmEx20g605NJ
wIJfSaSRkeodXMFF8VWzThw+psOk8oybdkyutc7uYmUATMnx0vTZPsa+rE84yeO/W4PnP3Q86p2Z
iwmJfMZikAQjUJjBwc19fz4JX4HmR+HbOLREm9ggaQzucxIxW6HvtWe44pXRHqqcIf4Wc8Cm9iC3
UE8dO/tm7vR3oTDxIEFLD98Me9mZZowXkewGBeyphWd5E2uaPfHiy0NU7I9OSE0VnRLbLXp9EzPv
Bh0wStzM+KXxJ6FvJxRgqVbbYD10mV5mQiOioaN4YFcWq7thJaeV6CqvBy8neje6yhB6moM7mPjA
JVPwYLXUxWLijmSgD1lTbsQHAjmIqvFwtQ0gmowry15WdYv8C9JdWnqK/3g/yGRQxfOuWyEiiNSG
ZklHY/AyjQsDf5FzOc1/lvlpI3RJ5xGp9Gzp7OMocctKqaI4Zeade8Cy5BaAIaVFop4jFhVQ8PAQ
WBKOfJaONDRz2gJJ+FbBkvpJUXw61hIQO+Jp2UMaeuvj4Wkau9DlilPn+I03IQI6p1XVwRw0pn/R
phImoNvyNSozYMXfyhG4DnhqEt34Tz45OJmi9wivvtvq5Gz2kAlOGCEwByqtwrKjwW3MChhcENyt
3c4cr4QZd3okiZOqv1sV+uaweAl2gSDNhZmHC1L0w7RbTVYrj4j+htKQULjGTaGzn9sqinzyUGx/
MiRpvRYmDH+2CAJuUaVVlVK8sefgTpG/4dHAhAB7MA2aCmIlKCrakBzgAHkeoGhp61cIh2PwpDob
vEawlwaDSCnruwkUApAZrsIbfdQi+qtSkPvPwZ712rxUi9EFJjaa8Wc9wQhgieupUlpBuTLeFOCq
mqtXSXHKsRo9zQSUHLeGt7hcCVr/QE/PHZNDSQWVL7HV39KaSNkJRYq7X6RtIUzMgk4FfNrwASiz
FosZy6EZEFcGeZJwuxIXAlV2o9qRNOU5pGij+nL78XOkjfweBC8wIOGzMD6FW1ubOTpzCaXPmgFb
aRyJjsb1FdqwNjXtJsK0/I4tUtrQXsgs9Yqx+wx05IDMiSV38yz/IAT/i7BefAoQD5ZR2Y3TUh3b
7TCNYWsrSQlVUASzq7vPkEaTP9WmsL9SqH5t5xPR0yxqrNS40W5OvpoSfJM0ap/CqsIlK5hnD19W
KpABGTELYTNQdg4TzhssdqYpi/04SH6bPT/LPtyuj89zGt8o69nTqTQsECuNQGXnaek4h8xB63RN
ozLYfc8ziP/XRH6z9dQXeLyu/vtzIc439I1cfqporq2e+uM8rloTSpuAnVJHrqog/X0mM4niN82D
wUkRyV5qq/EeSpLeRxNEGGBJu/3W5mxI6TZNh6IHilh56SMJTdeEawzseGlIOAkjv/Cq8buXHAoP
WKo7L7XlfSvKZckd43WiZ7fB6sxc/tHvg+TJtYOmytHQYYinbNnIrtDlwORGYfSSGibpAP8o1koZ
1fdsrgdqOedXZ5qB66xV60c6Geex/vCzgP5lUsob9mnFAuiGd6ofk6OQjvMrY/ompSWz6dwoC/xv
sUVRvosaU2x90aH7EQI63ovl2HjAgU9oGqJj/5CuwAl3+VN2E/+w52zafGXFa7U6IKN/ZfPXvu1t
gvBhnz+aL+zkYayHlrJ9aRXjMTije7BjFk8sRhO4H4WwuGnE9rn5nKXVtuFc5+bw9pijIXDo8yyo
cZd54iuct33vjlrMQKowcxL2BNs+fME9mS4JO063EMGdwvWaA1CL+RL6PjE0SzPs2RZT0gZzIviE
5q8zJx2ViDAppRUjk73+zfnxDri8v1SDMPmC5H6MGnwvOA/HUmipGLdnNJZDobXpM9gf22DL9Xi+
eA6+abnPtk4CbvkIadtCNmKXQPh9YMAU+R6b4A9iDapamQAfxD/g+QDpnTjVr7J05pYpCZiWP7Z+
1dsoFmCqFlewC5JIOxFHwESfkmzSIywFI1qBNpwrWyMF9upaK/y1QV6PCLIOmUxInHKF9uHoUWcK
+2bTjuJK61d6O5Pm3H6DTGA16Z0kdS5N+wcBn5VDQr7rhlE29qpB/eG/r6Y1zESN3h0EXfhbBdA8
bISZ4DhsLnPk6jAEpDlJvZSYx+VzpnQZThCPnUe/G+ExM3asGZqWkKnMxuGlr55KyS8Z+ch+Urwf
Ud8ensx+zgc1KH+v/YK+QBdr17WfE2pZvgPnvfj+etthhAkAKcTVvmxLKZjScUq+9keGyfSX46N9
Ay7B/uCCTMh0SmO/H+NPcUhvsXbZu6/11DihWoC8yf0dDCk5NrJkQjQBV7DVakUWeIt8S5xvU0k+
KzeR9gZflV97fIFGYIasg7ljHIt3CmCbcY06d7oyRs3nIUWUjF33qV+lxa5FRM+7rxZGnDdXAXvB
in/s6e19KH5lSz2ad3yHJG9l1ahuFQT8ckmKJnjC7ePixsdBQj/ugLrWmj8bDCOtLL1KqgGuhCRx
jcwv4BMl7EQwc6i1qrgGFKqlrqd+nlpt4/bhVeiocxP/09fAcDh+wcT5XngT4mbBoblUs7eYc+nr
wq9hlKm1G4BkUC5t4rCd9qJKEXEdcM3iwY3LGuwY8RMj9hu8eguniA3RPPyI4dcmKNODq3hv4KcF
iV+HiLHImLwCR/3uIMWkcOQvWyUMRetbIGRbgl4LUsO476rgaDEgDWYaWZNExdh8CWTUoWSAiNwi
g8ZJ4gWxOhjszJc68X3JNmCe2suHWk5/76QW+U9cs81/sgITFvnb5v1NJC1AnNutKGwhGRtwF5Mu
6nCSgjIbj3rz49nNszjRWYM71VKjpOrug4Gj+1/uMvAIcfnELNJOFrJZusfjggM4+elWN+8sbxXa
py9kQewqd4EuNe11DpXX9s49yzSuWabgmEVF2iqTyn6HvuEHc5ziFWbz4cODeK5G/VVFW/e2J9N2
DuK4+J1WcqaE4PIk5DINgMlKTQuJ8vrnRai1XpZVrSTXY5132hSoTYbTvkNRYFYY1SQhapgFWuJq
BnST3nvI8XZ3n4oJiTDp3+5szU7vKppasIXhkgAGcF/LJJ4BGXoykjWtBXtgm0T7/hAJJn+XxW6b
we4S2O0wQZJ9Bt+Ln0pE/QmB1WYbxksBaOy9I0NaV0CbS+1DyRY8qyn2VYgUxnSGHV0cU9JjCqwK
J9uq/kziK5g4ljMTUkb7x0zdA9QMrvqlEyyxU7HsiQ0ok8myy964KesA+DLJAFlBTupPH1nw91Kw
Z5UYAZcRaX8vvsRZ1BToJMO2ZUeOFMXHqjl0zXzJpze4JHs151531ksOF/oA6PcyTbaPeLusjL+6
l7Z5pEG0Jvp98beoNVV8Yve0aNb7/hXxK5ulNxAJeey+mj7J3T6xATsa9a9EqCkR/8r70JmmWCHs
BTsTWzgKTpi5h5kqdHoewu2MccRgRen30nA3cNX4W0ygA2EoN7kthX9FzCeyF9f9gjXFQdobd+4d
Wv2hXw6BFxSRf/HjZ9cjT0QX3KVRY7KvzvYjc4RFwC7Zz5f66PPgzEWq64gJ8xt5wmbIxWEXUF+G
7sIXKmTqK6G3IQYS3XU9YSLb8rwQBIklKZz241PzRpbfVBQYTz5hJc05d1AMN8dlKjB0dBSWki7N
C4vBhRhXgiWp0wjxer7zccPqnjrtcfeCv0XXBqxIHNRPHnz43EcYLtjWMiQJE3w8xEyUDP3bg3NF
1ErDaWiztUgfYniNGLPK2VSjVDpznScNMoAxLuLs3QZ1IuF541QpN8FX4LSVxDRfR8jSd7dYP8fj
G1KbQZAT+XEKznkPBfqAMGnUg6C50Oc/aHURam0rqwB6rAILTiGK7358Bpy/sW7cESGWQ075NHF6
ysZj1VpFHKiUKJVQp2Btj/uHXAMjL28BRuDWUFH+eDOqDaA5b07/bJmaCZrSBw/qByQjfm1N2p1p
bdC4k/LV3hPGx0vbN3xDSTZVihUISINFfkty1uRB7Gaytiuvs0lOKleoyetfdqeYP2nV8Es7zehF
XjYdRQ7HKKE8NZJ3og9COJiSyLWqvV4jQLRhH6B/FSVw3Te8DVPv4x6E+A6wEYklpuGVU/3YElLg
zKTe7SRMRZcf1yrVZQVXqJHuk4TEA4dj6L4s63h78KwgGax+g8+SdGZNRLAJdDxChfkK9JcXN/wn
0dRBM7C76Re2RU3ma9TVeL0eJX/ExG5CFNA5KGxjkHQMXE+fr0aRgWNUXDZuwa2uH4Z4vBUwPjcw
oNNVpIGgmQjUrGhC3diDiu82tk7wKHStyJ3e3ubuseJyiI/ElR5JdEModvPo7qaL+Cg9UnlfjUH6
rR/FZF1Jr1rKU9siutNW36rIrMTulYi1B6N4W/9bK5lX10HNt/tw7DaujnniTQlPArOGkBf3KxU0
WmKwzRTPk7Rn5PXgJsb+uiTM48MHPvMDkXXt8ZtzKr6k+jvHmfwODioRsds9eR807CEp6ILaLSbL
FjxcP5NnNIvS6S29F2V4Q8NOum03YwwAFb7dK+gclVT3wwWp4crcZWSMrLJvqwZnsrGd7XmkvAja
x0SJrpBJ95CXx2lI870B4nKjmFOY6bggWQpJRvJSRkQqsDLykbDqJh4bKLvAeCyzlU3V8vfeA1RB
kmKulfiYpGU4636EldJmxdl0Tyn7ksQ7dZftuxhXfkxRXFK7H6MMQIqSxqFwZY7DS+T6tTY01UOV
b6husb+tW12SqlLJIWb7TNOg6lg/ztC+AmCBIiBbdiVapoMjDL4m7F43tsEHDhJEnemlvf1IYIPW
N0OK0uLpc8IOJVUnbwvDUXxxQpz9lcfLw+VUbpQHoAI5AecWmA+beli3VuX+Vwuym5eqHAsXYGr6
cF08+CtcJ0dboJAxUWqAGvjKqFhnHh30THRGO6ZLB1qZa892T5Jg4MSjdCMIi0modOMLfli6rOpz
V+TWqVx0WLDBS6SFSN2rOagOVWHfDaOkogU0u11PEY1oXB7e3ugyYANa8+SQwUu2pjS20km3IkZq
ghBEVAdgJnsm++FswJ9vSNblE0NtcXDGYeuNIzTTR6I//ob4LTp5ouxIV3+BjxGxcVbIq2ol+t00
/r8zy+Az6TzidTwnZAVhkyMuaCcqxVKHNb07pqNmqGL4OcIlQPBDb6WahOKp9paeBgE4vjijgYwy
up+8XiqKe7eSn+o0B0ccZW9Zh4rtwsngfolJBaQKl19dtWa43yg90mjd5sI2DWSCTGJNYA8wakkq
oqVOli1dv4UjrUoAIqdA1e+VlTPWKJyLE/N5Hws65KBDh8benPd9o3cOJt8IK16ytL/BP63J/2GS
f6qzfcb6TKICYDgeon8S1y7/1/nrYGwCyEKd366AMLObhRHfTKWPaFgqGJmF7vZe9X4Zc1Qa5eiM
XNE2M8d2VLxOo+myBUBHC3zN4Q371CmYUYQ7OoUNwweFneHH1mNXHzoO4uWKC1ayBgqjRBabu9Ys
pmPoTsq2moP0+nKV79Gl0GiFtIbw4zF6wrx+xpJnL3udloSJKJWSg4U9Iz+5MiHXfNmFXT3UexGF
dyWiqhEQAHvJyZ8mV4wgq7oVgpRoayTkeAplwvvKFc6kI01KqYdTcpE/PWY1NRyy8tfqI9pZq3W1
bBXfakkrRVEK6hGZSt60N03Oh9d0gtfVlYcGeDZKYhuTPss4pFfT5nWl/6JSH4evJ2+Zpmy+a+1k
xO7o3luzYH3K6oxGO6wRJpMCrJOfWiB8hcIuGBt906DtrqMEr7IZ9aFTUKxV4e58sJDpvzMp0/lf
thfmR6VLp+e55AMAq5eOOAkx5uXO/apXhSNwQGsWe6G/fmhJWyvhM153H6lMchnAjyHd6tTQplfL
PejqdqITXeHSGQ+EEAyLTkAbsVhRSGjXVNTX4HsulyLuUp9893CxZaE6OCS1aL7jTD847HUbG/Ph
tmR9DjP5A0UA/DYlsLDt76cAbFyZnWbjXpV4iQjrH8JraABGHbA8Holul4cEMOPnE5ePhyTO6nvT
SO/qZvtHrmOzzuzZPphGKjWFU62rcZCvqaojvWCKumccj4RRX1BFH3UVMaF7y06TxfpHn5tKoBC/
gpo5fGd54uu5l//r/NKyHSacUN+7TcYOSKZB8jnpe8QGqR9bC//u2y1cpFBLaFck0q7Fd/TWEo5X
NhMg12l7lNUO0NsOQHcV/T9ibq0qvn0omaTfCKf0Py97ZvZOcv4kfsuprceoEmIm8Xojq4wCPUqp
r1hMu1SM3uhdP8BOBL4sdit/L5UXeSCu3F56MgA7u9KFN8FCucVrr4kUuZ2xvjE01GuKwYiUQgbE
VX/Ag1UVW4kC8lEkCRwjGmkovNUJlDAfchjLGJTyeQFuX5GwKYaKH2r996/qcxYmgRyQJBKH7Xqg
dzKn0zkwM1Vx6U5CrEw5N+MjsQcWENYqVHk+DNzS+0hMgey2j0pns0+3SUR6uhAeaTIlKg9kYWio
QYAEe5F+520UUifiis9Mjyw/b/cFhG5t15Yf+HwX/3vHd2lTs5usu37iSKdEzK4VQ5pNoNHM5y2n
57b/jKuslOUFBx/6iokdcnKHSgoxbfHk/xGHJchRqvtBh2j88K6tZzEVRdDwkZ7Ew1Q86HbRkCVO
UmAAvwNg+VtnNwOSJo23kF1fXohEpzFsuY5bVZYqkOT5ReumUtf2O4Sd1nW2mLNMTVIqeUjWeNZw
yNEhWQ7i9owH43TeD5e4zOh1TqHZT7kdlgwgP4LPbkpIcs4jZyyKJABbdSl0ZJbOvQYnryakjLe2
c0HYUiV/K7GjLWwhnPVoN9OUuAAoC4aFulwFgqSqIuYlUOdHfgFOsxwsPs3ZOblhaEFgexHgcUYB
qhLUmgts9EjVFNMlz0H6ysj1amUnckrLV+cycjpRCMbowoHbv1PrpAwHMNB71dyr2hh3pkYfTLmT
PZGY75Gri9wHiKR2bgjIEX60U2IKmziRnWdt5XsU6+ZhZTYRXGIBpbQ9OKvE0BCGiMEhG7sYhRqN
/v8AYf0fxK5iWg9lOZNY+qOd1Pm97Ucv/5syMRyJzvw7YNYvolX8bBqUQY8uVQXgkR0npdrc1rnp
3zIqC1cqi+Ybrec4Zp0twx9yrE19+var39jt6j+vT0P0M+MvxOHUuc76SFD2wx7HZ6sRPJLbJqJ/
Tx/9SdZpOvGXXY54QvS51FL4REEw6ut05Z0EzNFx7zfZjpBU2fPgFCoTF2D1SCSd009/FhTOXNOh
bR4ja9BKqR4iI83ZCkHQHvTEi1K3BHTBDwPf75Qgzovzj6xXz0mlt6PNtBjn8KGZPcBpPyK7lfvq
SyHF1o1I3aLWsTiQGgnXUw8bm0UTSD5vJdyyQ5MBTYaGUMwu+sdqirmD9ghHCkmDptlbCt9cq/pc
YCKJ+4Gl1+5czFpjBxK2h39BG+z7SFXJQF5w24snpXlocAJeMoQd2yYTq3Qp9WL1x86n+T77mv+9
SPmOUhtjm+1WI4Gg9h4Sqv4w65fLgAqQiJjLXa6OlKy/6MJppu3UyfcvSWroKr1b3R8uGylWeGaM
Jb3dxXZtcby+fXoSZzuiMuRwmZDfRsRd965tPWb2k8JDVIDUbekmEWC7D2UFXsMTZ3O4WZJXc3AL
npSwaym3mu6xKaxPDQjDemrFpjLEzw7QSITTaSBm/qILiRbfN9CgNSTloKL6bAA7AA9WG0cYip2r
0wXsB+yYScbVOkeKRFlpJm5JcWpGvpASQkdmTSVh8fyYR957oRooY6tWXOtBeuGYtBAdlRW3EZ61
FE9CEyVV7ANU4PZDSt88kt7DM0yAwSngZex81xRYpxAj3iJeCLwAiFB6yLjaf1SVP3tQFssrDplj
Q8rdlyv/oX1xHMw7mh8bVsK7CzC1ChzObBzyAUZ579rwb/8GVgckra4SxVTe2pT4r08j52OuYUzN
uKPxcoEhz1giEcGzuZePrzYFo5K9R1zZshx3LlaU9kv4ybTZ0Vz7AGSttVQ0JfMxyfAxmzFZY/AW
SKiEOUWjbrKMEkFSq+6dyzEWmlNcsOVoHnJXOZcsCn69b89CNSq6mBFSQucbKiB9DbTqcM3QTn3j
mABo+rdRAPades09RE4VvhW6I1vXjL6nr/ATpq362m2U0N7xwjIwAQwqgVLRqS8LY1hLl0tfBo5+
p49u8Jxn2QYiCcTp4XSTpHWbKUXPafxHnyNgYzSIKCByLCN/cobe3VNgVlMv1wcaeubgEWSB7RIr
8n1ar5A3M5IUKHDBSUYJpggLUeVoUS5F1X5BkpqyLzDDlGUIuaCW5Xcd4R6wO14shagI/mbMUfGD
6CYqazBUbOfvm426oIN6zHCw5nTYwNyIiElYpbtCH9gdueD/0ifEjDPBdnw5d+4HDewOM92lUe4i
ZuemrDH0UkloR3yusZm5zXLKWo1T4DKEgCYAZAjK58IJ5ATF/vjJkbgRt/AXT3wELZglJYcjtjM6
sX/2zbEOayOs/MrYZDe9Sls5ZmFyZdgmg6MrW8W7ek6YnOMS7F5WR9XQFaoY6bspZkkOBF5/slti
eim7GZ/YV4BKbube6upKYvIPqL3cjxu6YCCAp19FW5THLKgGahJqzB995fCPTg7M2FbPs4uFBE4G
7Llj8lCWdFx0jItd90wwbgpQjhhukGCeAnSR8qC5aTxrK6QrP8kVvQJJNLsxxcm+b6I1FIoT1bRF
n3kOb5//pDL3eUyMvwhvbjlclEjE1C6OSGY4xyDjevsX5fQorwpRlvngZ12edYeuyQtI0rXtnJwn
hzoJQEwMeupBsBULISmE42N5rgR8+5arThF2y56iVg2NLk+UsQjbdYj6u4MBRaFRVbiTlgfCeAGX
RGb8bdgMTlMpFSBk/DFTgQtnHlVtGzcxn2M0ChlJwLS+I+mtf+iDKsAebk97g2Ay79MErVBjzzdP
7dAQlidCrHWZMRA8ub7VA3p5EvF7860ZGLXrhsOh6a7eHfIbzWySJRkAlE8KNmQakw1NISOewmnB
S8wvHq0VyOitNsMd9WsiO2tn8gxCuvVZsxapJxr4Z+/flS4O7XYmsVouIjjrp0BNniqYPh33nSLr
oKKg6uo/9xTa3w0cBl3lYgJb7sdixzkc2JbDjAaIAKsKzrtL9komWX3/Ey5lHv3YUxDCEdglCnZB
fpkyXr4CoF5KtKe+5Cjm/9jzLMV3rPNtzUjp/5mQdHDt6DPkqwANbl8VpkiBmjKecQhDN0qfzRtk
P+yxy9FE9ZJSbqVuZMplrnfFbAQfyXijhfr3fNqwJiXfbhMU26bQZb24XFGKOA88fOVqexC7rcf4
cY+ykbPo4ocp/OUw34uZ+T0L4rC3jGqBd1ZRKhHHbhqNGnOtq33Zg5hZRbRLKWvdDAL8P5K/GGh3
MTU4DY5It5JvSMeuqvj9In0jNn8YEiD8CfCBx+9cbzHIfge4fbnQe223UBNT6LcAc6fqpH8H6D6x
ERcunVakAap7iiopuvALuqparWZGbsTnPtyL9zzd1cYo5u6eyjTZvziFs1pt/QyEm5MwDm4nvmQz
GSAJz9FCM/MhyUa46pvy1d8RlEr2GCgPKTHca6FyowmWk8W/iNBO9QTOtBD9Pr+b56thEUu+gTwT
u3NA4bYxhvkt72K9MYuiy8wriwi4KZdsvcnycVAftQ0St2mmCpM+K0IJ2KgVhUPCkKFVFPnaTyrC
XxhN5mbzsDtUwHUm2YVJDsdpwAWKN2r6u79C0iTFDY0fcI43ygdfmLeDLssRNOu0HVF7JUvL1m5e
z665bo5sko4nUFLCfK72Z0wsNqxL2LkT4Q0P74xmH/a+fseWUgmjm6p2zvhR2T/8IIdumYdK7TCL
Kbuh3mXSr9RlC9OOKvUum0+IbBG8b4qLGxJ0GWHmUHTtRL5UeXzJYEQpQK0sxrmn2AtL6WBfhOa+
C8AuEeurOwu0K3Vmk2Jm7tgySA9JeiXlivu8DjSbsMHauMNiyhuVdHGBzhbgvfYE0Kew6Fji+vH8
YN20GhzgOGVgUdZ52GxRAsmDptgo+zd8DPYD7UcnizQ9vbcUPistpEqIfr2ch2uAzwPLUtLnP/IL
e7oPoqVNzjNg4kOPgUPs2gwcdKe6B4m0POgWpQEf5sF2EKKpB+9rj2GK4MYjmPBsu5zl7zl1Tn97
Ssm2aN0yR5eF4Ahk/elQQ9beMya5nWbqgfcEdHkhy7EEhhz3bFQ9igYzmWfkNXl9w6NeAsBZyqWl
gZqel4rXRzZoyjombTvcj3DTJKxaShuTmudDtfjY+KpZGmjY7UwVDSAIUDrj+irRUYwrIsfFNw6d
Y5LzEOAaUFhBt1DpE2sDusKGFWnLsTxJZNFy1stgkVdw+skIvrk6w/3MTyvHxYkUYtLIarOM+igP
yHXzsodzPWJsWnx89pSFSX7+rKHc6rx6uYjR6rmptwPPa22wlNPqQfICWbGv8CkFN5axvQOJokdn
kT9fYNcMcGjVziY/ByslF9bi/C+9HoptNwKltXyU18EjXTwcRvgnIf5lO2v+zyMPebeE5C7gKiZc
Jnh6AoFsnBMl+QkOeV3pIJ1bfV8kBr26CbjAzO7o5L3kRl2Lo7Yy0QOifMidmSEDwWtq4aQ2kgXe
06VWI9aVCIMe4KBt31re/5AGaTG0vn+euIlb4GkdNpnvYLeSxF5V7qxyIpT/YXX+ZFDeNy0J5gDA
adLGIMain8fQk4hWEtUMvAqqVRUWeKCPsNiq8SGXQXUGEBPqvRpV0po5oNMrptFJuNuM25oYEzdO
ZGQpCeISPx+jzNNwajmqBmLqiszUO/rJZZlYZIVbgtSRwtVZl+7W9Oq8p65GS1IVpSWC85hgBbx0
jIlSkK9orF8dm1KCD0sPkYNXMCOTsYkTrBW2BAeF0Ik17UofFeK0UGyJMgo1MGQNg3qYy5bNHlt/
oZLLT7Ya+nnQ7Uxw63EdBFPkBG0ptocdxeJSzbBWJbpgrKyp685XwFr84wOoV29E3vbj0dRB1vCS
2FtMN0Vr3mHiQHO6lhRUxv9XfSKA2EJcsq69HB9aLJlfQw8PVOJlYLexzVltKJaw8YL1VxXl9c36
Kwsqjat3pCYOjcbuiWGRYmRLS0v95xp9hPXn8exLtq82WHYSCYKAlsnA0AZnk98ukYPKAfTToAAS
Mf1ILAbV4CeWz7bGKTmj/iteeSIWfR5Jm26d5igvV9dfYQkXw1sxLZ6oN6pelCbW5Jfg5SahNzbx
dRZVix/HmJMBgAhQ56vrC032NvwygZAMa1qcf3/QNF8AH7G73+pRfAyO89NjiRUBjBdC/7wqqkKy
7QKOPM37dY2gXVi8i2JRVN5RZIUb9/X1c8U7tHU5DPVabqVn5mqTdJplXIombQaPBHpSYonRMyHh
XroZdIENvayuILdhQIW0BBu1dbFtzVJ1PnN84yl/ffNNudQkowJ6K1uzyb0SNrCgXftAV3p88wdU
2XY8PL5vpizHsCfLzWryQT2yzzt8W93VGOdBo6/buePyMBnmdAkZCkbuI3lfHUDtSREL00qsoc1i
5nqcA7LIkRDBY+0T2tJvVWzxN9Eccbr/RiDqo+tr6RxCTfEwY1+WwsH13wGqEwl442H9xxlmv4KA
dFkKM7Tqbeg80XZ9544h3haVvaId0wWK1282O0LW0n+9CVV7WhbRPYCOPY+GXqI2zswMt7plz/te
/VcVkVN7OSo2Lu6Ml+XiQnEDqYpaRDZFeLd0hHKpGSOUyamcM5i9aJDnZu79oBoyKtM4iDE3aCnM
2e6YFN5exCl2bIIl0s8l2HSZ58I81bmfubj1BsipQdDUdbQnqplP5Li4mVKnuF+T4Nwejjag+xZ7
uGmu8Grkou0V0B3GOQAFnbJttK3At7Be3PkwpBsuvXDcTwN5+XXxwvOxbwLCSDMnNT6ixF3i/0bI
SmeJ4q6fhb/awdg72vwkS8y3BZgUHmQjY/AHU7fDb1gSN0vwIv5FDBoQ0xnvC+gVBTR7tDrv8ZvL
i8JcWpYWnCmzwR+XZeWjK6JK/Nt1F/uMiihkDgv+y9VNP9dZSrXglgwt7344QIFb4YMMMmhKI5Yh
/rS+ICX7iCWbDgc9TsltsdmuPJa8FNCTSjIHkB1vDdYlhVraIdUfMnRGGuVTHfe4bG9Fxz7SFFzH
20VJidE8wCXMKwvItANpjg44Jbh5K0aUA5i/SA9ixcTAco0ac4OcIDzWcS/jr93uDxiSqKv6OWtn
RvNtYxaz/Re4xnwCg7FyZqFymQOTzthsBcOrFOaqbjCU0Hjamy37TmayD7Sp+0Te0ZRxLqAGG1Y6
gInLuz4uKWb0x1HYDjTR48Up7PzQ1rkn0NvPj6xfQHT/z0k5cz5UJ4EA6WQoH2J34GhPKTT8Y4EQ
6qEQ11H0Wo6iOC6rSP/SVrnoYoOAA1Js48ld7WaaOt2tnJ1kui2zQam6z0U4W89c4ET7LyLuvdLr
8S6UiTCkVY+1rvlMFLX0vGNDPofR0PCOhWRGkiU1qWQrr6yK8e6KuDAyz/s+QyiWLRuDXYfhHlNn
EGtUGHgVqKfZDVO+5nZ2qKEALAUf3+fRpV4SZPKQxpMI8T9zsz8QNZnu1Q3gmt+SCLmZnbxhc+cf
El9BZ3UHIz/IjPTUsQ5DXQmEsoQaLRVQ7pPO1VhsK7dE7iMfr2twU71xbRUW4/9Tq45vNh5Ebt5D
mFmyopkedPazo5EN4TteITT3Jp93ZbsFdNmC1/8h208447Ak9p5XYxxYqlwAFjn2Cxu7Ehm/E9EL
T29nz0LUOnPGQsAqUvmHbHDXBuMo1TllQ5gnublsT9LBlC0d4ylsKpHt+/rRZpXzLKLlgIyxYIzQ
v6uEnA6q409MXfpufbmOzmgE/br+KmtHhyAosVlZtj9p2PBF9MOEShCRfpqW3KcNYBEQYXobZ10r
iBrcYlpl9LiTsCp2x9SI/bh1HF2IjQGvznhrmJ64tmwYaBpC2eO2oOq3x2rgLZqzryV8M1w/vE+0
3OPCMblR9VItCo6W25Mut4AYEbBfWPiKGnPGbZGAHCVCVXoQXh4knvqU7mXNSAkouuP1MfjzxnOr
c7jPqO8N3EOjZfXfLu3KvJbI+wICsVqnrlDp5aHzbSXMWT/76gyS+kE0lBXm83cPCU8fPHzpjznd
UGUZnSkq7KxchFsVqjVi265IQrCBGl/tVdBUajeUr/hf9Ntm6MoAxRMCt5HLom4SW9D83xl2GcCX
UK4B85LcmQPDZB2kN4MeV3za6Kh5E9HzlA/u26xpNBrrKGeqnEL7tKzjIfvDC4iWagBffe9rZdK8
LXGZEUaFiN20eC4fRunwq8f1cJ2S2YKUuuOVC46siX6t/m0JiWtRZnr/WLYJi4xR/Ja6A87nn7W2
5/cseFntK1iYdRmVL654yg7YzunNDWvcG3p2UHLgK4Cl4e89EFQJEonqYjiBFarUDvcq4jj58uKH
MzoXQhPcf7XSM7AzCUzk8l69jNOfnLfzymIy2uZGIAh8P9TtyAyW0o0lfMclmEoXv71u9dJGrUbn
2qH1a3hciHo0kdqkWygjV57LidbKxNOeJfbB2ZbqvbCwB2IQEVA+OdJzcxmjnlY43nh6VWi8w0dj
+2yqkakXEYqv7YtqD/HuYEIyN8ceU47hY+aKuxX4EVT9X7p1FaN3JgQTZbtp3JTD9JgzmMU0+W9W
dVQQiK92iCiRKdQbjqE69MhjJob/cOqlivykW//8qlFFdY+blp2STd05ybP4Om90mvYxSKeqKAKQ
16sHZ0WBeLf3fC3HBExToPi18qJhezxepVjEhuXVoaCt6318K9tA+zcF7aClGuX+kHOFhIUdDN8L
NOtnxsUCMXGnLMqGDvZHkFjLhwatmR55+Ux0VI7wxhadmdQst8muqQ7XIx2KTBSQI4s2ojSdM7GY
PL5WdGjqFiqH/NpYWYiC5Xb7L6iLEPwCshOU4B1eroYri0iY7I8OwUTJBTrMAszldO+c3lj7a9oh
OswsPnjdqN23bBqlHHPArwdbr4Lsy8TeT0y36zFH2wmilburl0ATciX6Tko4I3BHva4kbGLSkLzE
1rAVYFxnIuJAB3QJAsrcbc2vpYJaV3ATzGXQQas+TXbBa02XKoc41lNtINsElVV2/HaE+KLxPMJd
mOY1S4CuSsUnat3aN5c5NK0IYhyQzBaOH2D7LPZGtGcMGoO1URJz4+iP02NAiUbcIr35ltiMU/5s
FHVoYOrGQz6NXYQazrrwp39AqrjKzNia8sLXiUDJqeujPIfav0KpsbiODgpZArnrCwswE0kCs7jV
EFmTcPKFAbG/6/qaK3hK1nKav4XQfztUs2kbLazEE8yVyrAF77ofOKCHGH/lm53xo4raPwMXH3dM
36AvWgpmB8duMgSSEPYvKbKmmk2qBh9ccoCjkR+W268W1KydgGshvw5ajmguZDwas2w2xdBhmwvb
Yr3GSEUxFwhFk8NsA2wVGGJpOYDVEtZFqUXngP+4CxznmsMJyuSugQ0M645nulUJCjT4312Dx35c
W/9LFshAW9HMiuUbaT/GGOY9UaRKHOXqBXzp8Zeh/PemFEPmk0QRf9r7Z/m7qjIlpl22Jywv3nAs
wmj45zClWYr+2zardy7yb74e0yjKM9Y+s+sP4A5u/OvuRLgnWUJv+wf4wNhwWtmPPrRbbDVk+iXg
bF3H86OvE8bYLENVbdVqaepBA2FBT3/SZ5eLmu21tzsQkxiqTjmWW7O9f/OuJV2xlJmDKglrjjOL
RO/gYP/jl6fPDVRBjvEi6IWcLbZDSwCsUYVfjzydqjk6sDYEPyBcSfSJlV7ugbC/ixe6ua8Kf0ur
XVnolRIoPBIgQ7c1UnoXU0lP1w95Pe28B3TWueqUxqsGJkuBhAWhsn59b5pmUh/HWYY1oY1jCB9s
G8IKd3eQQ29LjAGVPLc9CCL9HZpZQvag6z/ZzSpJ23uvSUZCqGskH9RoWPVN9+UOGNKT2DZjg0Yn
Tu8cjaHYXLNGJ69v6FfekaP02kfaopTQiJmGsr1iIG1jRTThgJeAxDze+JgwfpFLsK4AjuKAJEWj
qf/vvTx16uUge+3JoNjVNvooiy0RPhMLSM0qIhaYWQi4oY9BItG+LAK/Xu80280fXdvIYVSw6jkO
xjEOU8OzX7Pp5DB+ACPrY/dHSJxHeTUxB1ahOzSX4qzlyRmSpRPOdBdtqJ3O2P7V1nJ414S5TcNt
9ofpWhIP/7LzBnhBB7Bqa7ZrBQq/dhhVLHlKeTc5aI9PgCN/NLwQ//y0AVfCgMQTGLYLCkQNloHg
IxeUM3OpFmL9Rw1We5+gXSw/sndpKPp55vrrwoeF0iUihSUcg4p5ylzRBQ0Z9RfZIbPPUD9yRjTZ
nHr8P1SJg79lWzzihthMsty4/ydscxe3RWFleXS7khQ8ZXfeIzhzdZOcwSs4j/e3QG7nV6DxZ565
VZOdY65i5LuJlZETvleWQ+axUbx8ipCRVPEE0yLm6IRg6/kQUCkjneMjl2l2AXI886PhwgMowxeS
OpTloa0AJPoKvsG2c7rl3wzlB9Ge1uvy1ob5zWVvu3q7dsn0RhGXRAyjdhzNj8wrjM9YUxR3OJ30
F5f52nXKTk0mpxBZXCX8uTOZgqlOunxX4qoMUZMmZlvagopvLVPdfy/h8POpwPXzuNQ/CCgeMcbM
m30xuDL4KXsL/iTdrk7Sq2VNPgYsUKiBTUg8AkCGuOzpJO4QCkg9L9K18W+srOt3zpyTHeigTxs9
qL/UIpPYCTvKqva9p82lbNJP7Ko/mCFuNrc11h9dxThH29D0O2q4lOwEoOrRoQ3+GUcHXdMW15ID
ijUE1V6N31I2NgNWw8WI6/lqNDyz4J4SGCDJpMd9QhQzPBp3rUTeXsSJ7Jz+xryoiTHY/aHRU5/Q
oAiEh2Qukj2I0/0l0Pd1jpxDXMvNfKORbp3nFuGpTd+gG805sAlBpWipSP4acYhOUCLkB2Xrm0du
mtIlGRNzsbDG28PCi/p9W6lMbZMmZvkE6biRYicxlr9UuMAp00TUJIBgj2x1y0af1ckWUqqoyuNg
fkKKplxYXM07DEj6h255o3Hh1X1meSEZL+SqqK8KtohD0dCDZ3iQkk5MCv+5n02AP4KH4b4Ktl+p
tTuFD47fYkeu8x5WrFuPuGfe2xmR/vKoYUQeR5asSx+b/pErbb5cCUlIlQjgoSe9QtFgxrT6JooZ
XGHrhsl91i1TZcXc5AqUU+HsLaJ1P1DK/gEz7su3pXBXJ4zr1sp8L+/nSzNPlcC9BCv+uRRcFmF/
hAwd9rZNoq5g8on1QIORFKcnhOC+ofrrOgdHWY6yE1FK5ly0NYy777rYKbQgZbksa3AfSWxKINJz
WF8KYGUHfZb8XXhDuUEAETyZnH1LL9nU56mS4rnFBv70RXiFZDP5UPFQAvcmOyxD6vMm+oILuCLi
NmclQlqk0g16raUfJ+4puJgjc+uPlp4kxC7cGgSLzP1135DIPo3HgOwnbMn0Q6Zke38zPi7aLnIk
tEhRRSRTcs4NuqYrodEyrFhAK67FRS51YD48Knk8lsDOtkddg7HDKdJ/SZPTmW6bu2N9QSSLQKIV
vxt5X7lBeo186xw1OERtN85nhBSS5BRuuWNtq5D6WIAvxOmZih6VIypEbCB5qTK005p73aTEbsG4
Pi8zY7uznvchAd9UiNLBqbbXaYcmwyi86YSUf0ox4yfekLjXh8AEPzTtDu1vR4vlY87xoc9RdKeK
XeIr2nQorj6NvKcTC1fdUaXZEoAZBJdAkE2p5zktXkHH6amGBmx96+onCcm1Gq8JrGi45dYJY/En
GFOrCTbWI0S2NdclGX70p7l7ed/0HmE621qPmVxIB5eUBpM6NhNiBTXTQPo/X4BfdAzyo7jXMsPn
p+kWtZYCFoeDY4KJpHrF+BCgkUkgfaXgmPAsYa1B60B2Y0I6/1UrK/P6edt9hCK9UZm9p/O5VJkf
jUKKchd6zehKbS05qL/nMRRMzgRivp1aLpUJEwcxl65PpR/aEqbQybbnkfNvVEvLIsce9eiRh0Ex
RNka0fudHU3tyOcaoV6cXXEtF+fE/B9qo9rQ5g+OrlUxCtyIk8T8guiT6cNJsuVu1RxgvU7SroED
7U3lsWUvsF4UW4jbofQwFbLLusGuniFcrjQPaBSgN1/RifbkVRUOAZc+LmmUMk1F8XOUJIwZYjd2
r2cfFdogjyqBTCMG87Nf57DDKf1SSm2JTvJc9yZoG4aU40j+yW8+GV+S29SqgFFwMkZadVk/3pfi
1Nn6UYyzGDUMnCIHbOmddUAhy2ISxA6QBQMw7/FtV1lGO//JXbXqwJ/vzP9WYnnbjJQndKeEKyZZ
xX0Bmkb0o3yXGBDOmrpAOHZdXrSequJqWiwzdVZTWRbEeWaqlU3S5ajeIPYB1aHW0ZRzucTfiVAK
EEAMnzRKkdtiJSXsjPDJqnOg/jfVDqMEghyoLO6i92U6Oq2gnakSdaTASRRGes36lwATXSS/Xwkw
up+G5xEaN6GUJDnTjX8goSCwF8yoWWc6Y/P1v2Dx1XmyO+EsCOTAIkkIwXrUxk89qfe+wnwrBdlW
gU4rBb2OPC6ttNaaChh9D0n8yT7CKyVYQN2fHG+TVygYWu8ERFTWvJLT/3NVr5Pi1seus+QJPff2
tz+a8KMK2cP/6GWvijd9NYZLEpjnMrEH5bknfVBSTTIGyPW1RbX5vcqC2fCQJFKYO+VrfVjtYPgy
k1ShCAnKwRNTC4t7SJjnvb8BNF3Vyke/SvE5JM1Bb+4WmNSMTuKR/AW3GonCXG1weSeeh1QzuqwX
jAj5JuDdGkpX/7w5uOFjg0a8yAtJwrsEiy5FUqjtgJFlZM9SMDMaPlafKFpaYRa1CG8U3J5u454j
T9YbinSjQdsP+QmbW5fl/QOepm2Muoaj7hV/0PZaV6SKUst3X7KIGgNwuRhRbvldjGmjnuKkfsIU
zPlFZdPLwZIDpTcDR2yRsVRx0o1JE4FpT79faK0X0qgBFFuNFb5oU84ZcDttHAteV6N0Evul3FNR
B3Gm/p02AxZu5euy+iiF8yggXMqqjwDaIsQb1ysZayihXNSwQXlqUVazPWTXIVEOcB+VyPxU0bmt
uP110+DewSFNN/UqPk+1NNov+IfH7MG7U1FKmaPDuvkiafronpIM6LveoZ2VCPCPqK90/HtJoLUF
+jnlbD5a5eDXQfcPZSdGFfCFXMQJOSOl9Yt0htWNFffvJkiBJnEs22AWuhkwKAHMBDmKL4qVZm7y
5tj6AlSyGRVHGUq7s9yx2VSVBV6pfehz4LDUejTueJas7Wwt4oZ+nQyHinHyh4SIKaD6N+LHlbIX
jycj4V6rZNPbuE1JpdJYYXHRbxzMM5iKFGi5Nbm46KL21/2QJy2dL6z/jIu6TUcdfRj4NysUEv5o
Pz83C6DvHOTDTcIygBO7wNIyY9oTYgvTBjhi2nycs6/5JtVJ4SkqQceTvd0VoNUcWDDFWRAt5Jk/
DeGnj9eJC3cQeEXieseNR/5EzT3IL6R+8icrFZJPnC0kTyrURljht0xmCE9HCkVRBk1kLZ3lbhB1
eGRXRnZAuroUvVihvlZ+KAB7+UAX1y3TJ5xprtlumPwS65dLTbmBkxGNRkF6hXDCUtvJjqznb6CS
ykHTU9K6h4NBQnxrUiH06MbMo0XuRdmsipYXiApF2UcqmvDvEILKxy0U5G5ZSNq9zNidNvAZQYqE
63U8skCyT4nCj6beGeYfTvedgDwUkde+G75dGSiyvDohuRomFSrfTCM2bY1P27IzmMhi92v/dHf2
LoHBFKW9npaXubfDG0K8BXE40820vkEUlC9iVGf9phENVg/2iAuzZfKWSEd3XcHX6IG2oSXze177
35FKqDT50vLBY0xLx3SvcMN5fGN5Zjg9XyV+yq+0v+pMISrKHmB0NoBKzO/rHLwIC7k4ZXkOqh8o
E/mdD828RtJW+FQgV5nhvqUofGs8B9CUWT2ovLaEhBZhS60JKhKp5niFqaWHIlEFE5EZXGt/OtNL
gyFpPzQkjizrOzE+V6K07v67VdKI39oyMb2XvecbqPbZc0TkN4EJN44oYTfENb46KjngrImf92Rv
Wpjsh9h4Nmmtmkfuorg68sIShQ05weFTAFVdmka7A8hRB5ouEWxEOXemjxB6D/XifGkhAXqXf+dD
AeX0sVHRcBmIhnCUY/4lxKfCRHqnZ3TcB5krCKIIEpTs8ZKnXV0OxYzIEAaWiEBzv9Fi3PG/U6dP
sb56jEBvNmngNbzBipHLabNZStWHLQZiP8dhNX0JTCVPlyHm8E63uPb0sFu5fzLwhgD3LwN1c3hr
1YYwlmwjYY5Nz/rt5ux7QWn0NJPIC1P66lttEhIx7m9mqa9EXBfmkEk2yKrHVVERtothes5uYnav
uNRrhYf+352LS6k8yqOmw/o0xSPSPxvfwUkHcTOYz++NbuSQC6hr3Kn+6trQyytCLwvF74gTLdck
H3lwtCoeJQgmgs59+JxQjHDlyfmkKW7A9pu0H04XbyzOE0hcxWV6L099PeKt3+3Fdt2Vu4A+etDs
J8MDOQk7Gxhnl/4oGAG3l59UYA8lWqY5k5GYHI2JSk7SzpKVLKEc3QH6dk92EwPU23BijyHis+zR
q7YngxqwBdyt7OUpQaK6FMOf/Zjk21bRYPSq33QxMvxuzINPmXPhHY52543X3PdjNM0VoBFxb9iT
it1U2fiTRxqd2Zg96Lu3CExeKxOC+xTcW8dK5jChKYbUftM4fBfhGXyAbl9UVAaxNNtFuyhiH9VW
W2xc3mAdKWovBAZL6InaDkWHyEV8V35yb96fngxTnydsVOyAi9XeJ0LKfXcsP+8cWYsPg4907uvj
PMcSmT5K37MXL3gOw24BHXPlkjOSTpbzU22PBhyWexCvIHlpWQUkRaMy2J+YfkBXKniZX/XczaQS
FXJmRGk4fMjifuFsSsAGKB99/vbmwQVRV0iQSDDHOWwtOIaQB9GoV/xCZ587Q+rcfW/QTnhOKsAa
swFrwNrIdhNJDU0Sw4IyXbhoZWyNf9zrzdSsGfMgu0a/ylDvc0LHOdWHdOvT7eWMB5/ITxL8qqLF
5JC+j/r6V+V9fLvs+9oF2Tj8lMCKT9RHZ0aHQAQuV+PSM2N2LgiQDVcSMFJxXqR0mQg0hsHD8bep
Yx5dnWwkSlyTwWz6FRs7FKZEQa3DIWrFfZFxeb1QamXS0bjms7mSKX20D9rtiIQ/WDzd1lqVRnIt
lgiW2Wk5CNPYz4R7AvhY5GMAfl5lPBnmPbAOCOrq3hAgxRkwR4AUTF97L+intTcSnT8DIRAR0Y9K
2V30P9X3e3oL3y7U75GSzQSrpGhQPjfG8nDL8njIiDEp65MrMwjU+LOPPMx17fsSyg01cZwt3cmR
c9+uk+Sc/s3uGI7Gb/AStY4D6tPMqtE/f8hAVjCVYPIi0HiA8U5Rzlqney62BY2XwPzT81Lg8njJ
u6AA2mydXW19nGMUwwt1eKKl1stUkXnuZ3O+dCl2QsMQ+CPlTtZUrxDvO22A3fpcznHiMzsooH4o
iM7OcAQrBfC2SzBYfNw46LF1UCmLONlNkSrYO/W83g62j4agp9iroEgc9iBl+xyvS/vNfXw4zbcX
Wfdy5e7abGxqRE04UM4BeAmyR9GV3v66ImOvHhCpgJO8KarwQOlX2q7iaCo8TowZwmb/9uu/A6rc
WvuNxGetR7XTgGpCuhLDDAFxviSAcn2yVyzGxhBg4yvOk/jDSyl73QkNRQeB3xeG+q9goVDbixhr
QP6huI8r0045AqwzET4LH4ScpErfoU0wgx65J2+VpQgHn9rd6Ulru1aQ5oh4Hbz1miwV2ql6kdSi
agjK6qIXDgPo1uLcfBVIVPaVuwBZd0cBKHWQysiVE7MQpNP1Km53Q/KejDP4tay1K/D8BOCT0tBe
PY+KsAAWB36ky1fgL91U5Ll8eE7ooTJIDhshRjwd6XqqLOmeSrFmbIqOMYgZw5pcvdULC0DHjmi2
mz3qThAU8H0RlKUyVhjjshZaQZh3TXCknr5uOthpq4FsXmpxumKTtgWKdMHG241RmloW/aTHvHg/
aORb+7FuvkJhuAvxuuwXP7PW6ti/Wyg9xJVLMsBkJPmGzI6XBEurL1ST/44IMOHIuzqSFZhlt8i/
RdO9T3frbt3Ru6HG6FcQ/gqOMFyMUELWXSnpnbbGMARj7NHOhe+XYP0FsizznOBMeBGddIaPySLJ
GXtyQ1e/BITVMFisABEDI5k0UbnEao/Ty21+t2SPX+m3E9uKEIdr72G7Pe7gAtos3hPiaYoa8Evt
ZCNKX5V4oEqqL7qYE2437UGkzcFm5JHlHJCYcV8SfyxYdEJxdFk6MDpuqqvqmrxRHr706KPbuA+4
TULAASKg56ouIjg54CIEU6XFICFqNI4Gry+QJaLggQj3atkMZi/PvzLvsOoXnVltP4d+6KmuLfqO
VANSKoyTwfWgTHW15XSNJ3oXF6UrexSXMEcCPWBya3QxlRk0tKpDsNco72mXwqjpWFo0OKc+pXnP
0OTmi7g6dsaOxGfLHOb3dyQ8o2sLmsrONnQeh19RUyOfgYm88WqYWbZodf+qn8+MoRTYYGr1PSxN
BS1at49d1pfyM79Ij94xcR/A4sJMw94itJAr2ccLkKW+RFlsIc6vsuGTj/a1XvjR2hGHFHF1hOu9
y5ZzT3/jhm+DqS6Le40o0mKCewWXTZuhowHsH84pshBspEkE/92yd+YFmbULvW8Zki60ycst9tiZ
WkUX2GXn1emIOesM3Ty9gVuqNEGn1tv1WV9cv4aJ0NlWKI0xaEmhPxq5PEx9pYuwK5e9mQiV5Bmo
0i2JSsw8SCxJeOg2o4zYrwDG6sm1w8qqEok9aHnaCWesHI4InJKeu//WdoZtoD14LPRWbgINA4DX
Ek/uxfbsHQ5ZD+VjJU1e+yH5vcVbTEWi9qGK1vM54JUBIugEnPOZpb4CspqXT8MWPlB006+izZCb
5R5uG3BikfSjbDbIzUjH6c+0GXxopg4KVjxBHKycoo4KN3wOK2zKVcJKhWPt5X3SSqfXAcntyauX
uv4fQxArihbNTRhF0bRhMLMPt9cq5+NFBZYJN41nn0d4qN/ZHd5/WV+7f4ZljTE6lkk6eEKKKL88
E42c9MhaH5jMu8RY87xGKqTJrV1GyNJzUSkMuN3RXze4mXCCSWa7S/ijm+wMgjaZh9hHCuNMOBqk
BruJrfAWbMJOEnoGa82bUt4PcqhvWWL3RZ+dAVTMw0Hw5ksTOxVOfvgNTaiV+Mwm9rz+odB8P0Tw
QXOTpbLyg2e+enek+LbUZHMwflmo4qz/ff8aIUxN10pWGRuMB9bjw8Nd4GvLeXoA4W1bJgYv7gkp
Uf4TdrtqizX4TwR7Uj/m1/ygJgVhIA3cGu0dPNKvV+NT7IMD/5ecvwrw55T/8fRXAcwfNHSAq9p2
/+1+vq8L4b0L8LSb2aE4KnifbkvjbSUSQGs5UiHfFzoF8bNpDtPX3mjPHrZN3ml/zQjf2us/91Iu
FNOzb79085YdX8vBA+MvW6daln9JiCiEZ2hOjbKCkgVpvVYNsgw1jnG8ysO9fGPX/+EAD0qv0h7a
dh7s/sPQFxkhCzdv3IsXA/Hv1fw53WrDCL1c9EW4CVslEyb4bhoHTmqt5UMglOCKDFT+GJ6mCFkD
AHe2NoBsN8yVeJKV2KHg4RacNKPCn+ozqus2tnj5UM4eM4hOcx9TuGUPChBz1m2tJFhTedno+cpU
ltRvD7tSOyl3AXQcXPM1Enon0e1UdwEU5GAKMKViQTPVpFBJAJCeo1zrfMCTcssL7pb9DAOogzir
FI/hEbzZ6NCVeOi9RNolg5ST+wF+W5eP5YorMgIdO3DZWZF2eOknd9CQD5vYkpTxxerD28De6o0Z
sZKs1vWNHj/wG6puqEcCdq9zJ0GlRBdm1p+8umLQtMSVgKHLOTO7BRIpRCiPOwGzzoTxelRepO0H
kOMIiau66SdsCgeL99dnQiChFM2joMGFwOD0B3eFKQ8Iyd/2cht6kDq+TOrAXsH9+t7TH/URh1yg
ARkTRAGam+ZsjC1D7E6By503wzYH5TE+EcuwGXBvFvPjeSz7eKusKYjpUfKRulCRnVi+LmjtPP6J
ChdIF7FUL+6Diq+wwASe4RVVeXoa45zoaBb9OWbJFjkogg1i7UypfQCeqdsHly752CWpkvatI8RB
aGl0VekVconX/2Pck5eo3VNbgh2JJICpsCWrSz1HCtcXrHotR55/J3A5qKBRqNU3IVamkPFbYeeV
CEAw05W+/mTmwDIJtu9h7FoSYZx76G04LThDPrqAWN7ETREx5pPypUVh1AM051svxA3LCArv5HFk
5x7tcm2yDCBwcTmcYDEFluzaMIoeDFqMCEgbyX5pOWskc/Fp/p3A4TpvcZ1nHKPwegaRkUFa0JSP
7V/aIwqj7Zpek82Os+ivvZDdY5wWLT4KCh7RbFhUMqUpOlFuiakWxaYKVl3AcSbyMHSHk+BG6L++
ijFVLHhIbgaYSeM3xDapO/uX6ZQg8Nzhdd9oVIU+SjoVvMrRKItdi4hKP5Kk5cVg99A+yqszFSrl
1Z5vdOuSUvv98WGiVELoZw079IptnhgzMhY0vx5DYifG4C55plExp+sBQzUYt+57lXPvR2duQ4v5
JWzxQoK0UBLaNOYtDMguhFhG6X43kfCUupL/QI09ce+F/FYCFzU0cpggeegwCvcOwINOGeibVFhU
bCfYBirJhqlnTvof4v0qxsnKQ0FpWLLtvxDXjRy6HyMU6O+G1jY+fHmE0xjOlctgpApWl1UkeM+0
Q7z3YXDG9/7RhVTRmBAJ97iKWTB+F5YrKyyiKgVkUuFj0ZGtz2n1GWf7I0X+AGkbD5Ut3Z1qqSZo
zjYemXCjfyrL36JxJ5SyMS+p9oIfejKxPs8aUkXtYHwcLRhWbpaC4J4LW9OUemxvT8Evjkuy5MuL
OOodrXzpau9NTAawTG++oY3E3SgKkbXebpMxIeGWrUEsI2MpPHebP4amacw0l7UEcL+Q6d683icL
lSKXDJelaBX+FMjaW/bsdVNUd08CqLmuW5u0JkSis03KDPDg18k63G2BCz9z16naQj4Jvtrz0ycu
xWjvxlasRDty9LhmbGwPGguHajTbcgKhJJ7wb2LwU6cbzTu6UvN0qbylxVDCuJ3OsTEbc+IUMvhK
/F19c0j8cykVefhO6g0ayO6S/dC8nE6mmlnPnI3UVKsG0B+b/LDgV4SiAJ6/ZmguSeHCBBchItlP
Vu0GcbS/z2LjbiSAFXkAC6dLrAnBonVkfUSMWWa8pz/ynTmH+ffuR4TurCJ6qP/udRP+UL1ArbHh
tLhkpEo+rd+XpweojEezmueK5o/QMG74TPZdcxcWhDHzSqDKxUtWs5gA/dlKnX28vBY6JlY9GJVm
kJiuHOZopuY+41ViStYUMaGg1MKC0xM9xojhU0fQ0BzZWZKSA1ae+COTb6plI7fIriNlQLlIQSJo
9oxTQdz4IdF9MwJ4eLPA+FDfOuPD+6M8SbCm67sJoHQrCg0HX8XaiW3ofGT5h6CeZLSYue54Zrky
Ls1aH/bFcG53E68HFuFZwvLKfmu64kehbyn+hItCKF7b1VcosRKc8C2IFDGgJ9FtbzPzErw8Pe+r
6JpJpSrJAAIasCMQi2QTIipGLwT8cI/LoPT/eIHQb4lZw3daLLOHiDfp+Ftd68nhiYgCXitD3Lcr
ZS4ua7OIg0YxzAVh0Ns9lAJd9U2xL8xL8lBq5AbHY/gesC4Y2IJh6dJD8yo992ojxAopFCqC9vSK
ZtuU97nXk0jabLHbTmVLDEgEYiwoajD1JzOrdPkoRE8QvD5TJtkb9zBHj25uVEwnjSphSFk7Fops
PhumGjKeyii6LHZFfAgyWPq7lPNRAmFnFGE2pHYfJK6GDixiAqxF478nZjCEJNXphfhhZomVkbJE
OVaWF50xsAm4rLbYCci7jKbpeunRyqoKo7rLEqq6M3suuD96t/jUCs3fH7mV/ZsEtmFtWX+qdNc/
7qOY1aPoWjDeNSulJt25gnqS4kiE9UhmxhyNyZhF0TfnL0ig3owQaxtCjg1ICVohnnZUuPiKZvKp
7tr6i/CZt36NKNs/vwiNnNuDTn6LfEtAMcigq9Ef6AK9Cu2zPfV102duhBWGGrlnKD+oxZN/F5Vo
WC5prZ0WxYnOCZ5som51hTGHB5SFBUSFa/cZvSRzuVXhUOBOwj+Lm1lxryHQxKXpA24iARyf4pef
Lq4N7GtvLBZ69E2MHURHn7MRGI0m62IaKZZ+MXntutaKnmOQDjMyZf4gTb3M35wHqZKC8Hb+zLGV
ss08WaeX3xQGNS0c7EXHvkM8D8SbRNJjugIyWMMp7MbActOJRo/VKzcWEMwEgpoN5bo3sDTHT7ON
CI4H28fZ2j8GGoPVFalcEng+lbEjtfheDE494VEiDHAZKn6EsG0HLtHv2G1wah/mKY2s4+aTjndt
e5n4DLZMCZ3wQNXtz9D9dNBoAKLjeRzBXc6valfNK+Wq4qV5XujAkh9EJ9c9fq3jc1srxaDKhxMS
N0EOYB7wrgPYJK4Kddv2KywqP+AQhBnithF9+iCg2yEZsM12YLhzTgSy1lDV+2EfejJQkpzsYj0e
c7QG3XBZ3dhWCjLHiQL/J73HNIh9tgqLJEw+ZTxSWCozl/XpITZKrseqJ2SGZfMX1Q3HArI/3AgI
LJCXB1TGxfll5f4dZCIhWiHY6V7iq9lk8pBuFRMWW+EdeHXkKienUKeMMm0hZb29M90bdYRuVjHd
LFfe/R//x3VD655l+O9XObcqV4NiHja8RmP9ceYXTGT6zn363JwyGrgxnm3zt8gV61wHkP0Z2jfy
KVZlX3kffKWPQKZnrk80jbY2wkK2pG12d+Tc9fFRPJVFY91zjwA9Ks4YN3zvA8KzSHEDGH2kAlIT
rcbD7yNdRfwHnRDfYBgkQHwYWA/88p4cfBPzxx2+tRalMOEUlvFzlEULOP+ukMYLnmDhZIQ6+ZID
4d4pjydm9ndxWBITYm0tuJLdU5lLV/7ZdQpeZMZTeEM/lKSCvqza2R+KwNZB72Rgf/iF+ix+3xs8
Ch+vhg+YdGjuxx0LTbE2Q0cy2ZFev38iNjEwA+L3yZZm2lHYvJbYwl7HNm+g0NggewIvBmnqRt1f
8ayLy0EQWU2mjp4W5V/CoeikuK4I7mC0mtUEYAeRgP6J706IbEaTxA27EvdlFCR84sRB8a76C+D3
52hruAxp4BlfWNA1wOVheuj2vpHy6Uf4stHTICHW6yG41IrWG4Jy18Lwqvg2MPq0aL1BLGYEuuMa
HCCTRiqK8X0lV7DIsU4BgM7+RZyJ9peIKUhWi/LESUp6ihaoUBvce3CJ1M6nhgcrq7sNhEm8AqO3
0lEfyc/0Ra3fPvbhmlKAYx4BdKf3BsTHSt5Lx5LjJtKIMuCEHZE01i/5wBsG9NkxxUkzheRlZfei
jgEw9jJWA/SfyqpXbcNjnCwJS2gUjLnMg//iWlK/NJhGF+twFo54wLzwZm52oBhpXCbhVLBp3o/3
cqiVn8HkdT5jEg0Aga6vFkHkO7m2qk6Rfk7T3BOco0FWBU/RoBJdv3Qk5gjWInwt7qYF4XDZGfd7
Ck6/6Bxzwb5Z3LB4cNIWwCPP4maaoz+nICK5If9UmnLl6cvmHk5/5w9vKSgGGwyYUmKqPgngLmyo
rDOvQkCVf/bUN70rrAEXsBmQr3jmNj2i3k8xJxm/9wQkrOtTR+zU6TNFNrAzKrZ4ZHUHrKUGi79q
3eW/zx4sbfr4vEDKNRAIzMwEgrKmJgrbA0MFp8wfaOinmr46UQ23tJTrzEfKrTfboyD1WK8AXPqk
v5/SdlV/Mfy2UGqVyCUtoNcKFfC35DL1nd3eg6e+zgJ3ebpFsv8627SUjSDigv7OyY6hjmZUrJv4
vlLW3X1STTBQet7xWFmm+5jZVhjeTuFuE7n6PD0EOksuILIkEqWDJmHQW582KfTy3e0jMgsBBXqC
itoy+BmAEVORgAKXpNy0L97CDsoAXyS+tpeoPk6FaVGoF2EdwCgl45PLaSzXIOOrjMpiTLV/2xNv
VNlMWVn0WdzWuhSXTday0zGeng5uh5CR5T8wPqyy9gRT/RFWQSDRXIOET5KafAPizNOvCqQGEyBd
K1SJ0fGQin+vewNFVAjxXxgSKtPNncdPmuoSyj0XRjFhQhACdGxcbdyE10whWDO9vIC4+is//8mM
2MDoUC4VLaf9huY3RQR5lEYjxAS1flz5XdUmawHkFoXYHiAar2G8/oXL4XVIaOJtR/BLaFcXBKrF
J9CE9m3qhTkkpdm3QbjjZIKnWlstzlsDp+MdYFJcmL/IbV5SdhM4d8c9M2yc12G6UCeX2KEIjSl/
6QuLXRTP/FxvbD+FArNvWH8lkbQRZmFU3Qo7PA4H4iZK5N755mH5Ztggjk7e4sz2OGuuI3y2RMc4
J/5FI+gHCmFU8/ivoliCwT547y/w9pUZozyUc+fuiG4Yp2B5XvMxGF/VQSwZ1XNOp8mlGzzpMS9S
6L9mYgaEZIWWNgALZd/NFbibbpNEENcW6dWEPABYsWnIBOOl7ejHMX29N4fA3TDSNSuxnir4Zmyp
pkKXBMhGM17zoNgJPEYDFpS5qUFuFrKjX5xm3agi0KsZh4Bu1/+pBw5oWAv0DdY/kt7cJCq40gqT
irMC7+u6t9AwieWc0jQ/8PnAn3iw1oIeLtB8OMxLAy81hr05T43bd+3XZy8YoRTuqFIZD8dUJa5E
SXFA6BjBt6omnXArhIDd29tMLNsibIud5btMX7+joWlWFs05YuB2DPV2JDrEom4uk4gg0EhJCgH4
STiphHdC4KUybYt/2mdpg4AcfLZxQoH+hcLGtHzoQhhfzE/cUzl8bjkOteqRX0IDaIf2K+poUGx5
SzGKNcGFWa0vVDCFMzd84fOAj0aslyoiI7OumNe+HDCkQVwDYf3LxZzBZu6Oi9hGl7fkeBS6vMr9
bxejk8g237DG0p76wWeoT1BL1/gWzwaROPb8pYVAbxRG795yIH8RmMRAjNVkIuKwAJT4S7heeq02
gU/uWmt/zMwVGkgfTwLOdVgib2Ubd7VLgtJvvl9aOijrBrAD1ApS07zSn3IQhdOmAoNdivCYmjRM
8QiynEK9EIe+fOZzjCGjinZ01cOpzASKCnGtfGCixbVGsf/gWyG2v4qmrYxCXrvW/b1RZ9Yok1wy
QXqfLyu7YzuLCI9oT0bMi/y4vN5xSRRV0ZwV+aW9xSE80cdII2rzp1kElG6OqNNrPf1unhy9BbPI
tXrHQpGzk4+zqMNXbjhaRaYCpgeKy95gMDehDVrqZE6UIzQYQabg/6Y1yl9K2+Q6J5/N1Vm+EefN
2V/Op/VR2JTTZc4FrHIR48IF7Z/pBxOkvYwcYywTM24lyQcWnw+uwsxj4xmS+Fa5ERL6mX0vKFO0
tQesXz1+97KMSiIzogNADoQ6KGhISqxTF51LT0HDr741EOo1vym4dK7jJfGCzqCX6Gkju7oLVQcz
UvPSXBa7DOErg7BSZofkb9/KXx9LX4uLI5DYY3V6jnBCF+IMvFt00R9T8M71/o3TgaWao/GCTXyv
VDePxTB8CG1N6jTuZ6HQ9uUEbi1C/aBQM7z0c17Fe739CgQjANkSUBMKa1kGD1XJ6QpIW9UysUDk
rRb/BdNPBS/bqfjfDs60Wnnhl8KivjROsa4Df+2gjoPtQ6GKsjfta1N5VaLDkIwh6rH1tGukVYps
vOeyQ4CmvKuvDYZYCx2pHxm2WF5CZyu1231XB6IS4RoGkFIJJ/ySt/TZ0N1vDUyBtY8h5llCOiso
sMPKm0BqeiIGgf6NA8gcmkLhmkuFysP5YHlEOoyT5GU7bka0ULJ0TnyA+I0jZW6V+31pmsbhVacL
SYyBm1geNW6o1ur8gXgUhRtsiXrbEPR54tVwaGLyVAndE2azVTdtZ+HA21qvC+C9bi17RMfg7wr7
LIJdewl5iSnJwHle1XNkQSKdIukhEFCurm18imI3gXXo+Bpr1FIu/o1qVewb282ljV3KssHqXZb7
YmCGC9Obh0WTz790dgX6GrO+sW78i8cOKyEyX//2vtTHOnMwZ8JfsoPqibBLBT9CuoypXn/q/EOk
ybw1GdBtmPVwW3MbX/rEW3RiUXa/R5GEhAmd5qQPCOSHgVDuTr2f4oPxce5KCP2ecU5A1Lf1zm4z
8mDa1KfTaD2qHn1TMPV74oIgyLadu1M7VCRsxOGPUubFFLZDQREULYzjkJ2Ni3sbt0mCo4kzEJ9V
vUjCFU1YISyYRcxfMaehGl/MY6QAMbbO7DUmaoflMuovXBPmAAn2HrBaEJvpyPegsT7lultQ4Mz2
BFew6UgeQklGZEoRRngttTEQQc5YCAykIRkyxKx6IgbxI9W9WK2fhaBMC+f5+uaeXo1HG7MPXxAU
HKN4pBqXaCqUOVR1vdLHmswW8liU/3lU4xWXqHloeZLHrryoZkxq3iIugrgrJ/JJrCvGYf5BbpiL
UVoEgwdsqP0+PGO3ti6nS9mHrgoxRKUDb8tKS3SOjsqBJWi5UodJRodsILw24LKn20OabTzKQPwN
bSU+PcyX8oikM66tmEGxyiR6StqdRC+uyd1lUtFMd0sCjAZrBxFaXsrlcQjGrbS2XdOZiC21Jh5K
1tT7+Q3S8Kov2iZsSquymKntUbjVJVHT2fjYy2kNGelUpB+UZzdHQVyYPIsI3R8U7/ZYheKGixCz
h32sjIVp2nOS6D/Zc2GZHZwFgvCRDjuBFqRm7YgGBSv31KNlc984HxV+iKEs2IWL8j/V7W1ra7YP
vYBLMzSg3GMHq9+WP2ySwgNczCcR/TUQA/LUCyLyyoF/0oa7qCIkf7BPT6BJ0GxzkSxv9BTUgFmj
jhy/TWe/VoEXtdMZtmvkXEHcwQ56aLVtU6mAbXOKuHnn+SXFtUmBnSPgMxJekNw/qwPTUiII6PCq
Bkcxm+Oah1ukfkvzPR8uLYu0XdlRbQmi6WxDOfW5KgIYJEImffufs1v9SZx4pqXG+kdJLwtziCdf
xe8SvgQhUdAYIyfs9Iulh64rd8C7rt8j9Icb39fzSlPo070VEG4ctjveWEmf0mjGr95ssNbejf8I
euhDGEz4Yc/Cq47ha7mNLMeCfI4Yk4TPkpuRc49OXecVXJb3/ue2KsdoDMplSQvrygay6cpRUU7h
FlaJR6nFNZL2LycA2NAbGGStqLqVvvOnro774QXe3h7kY3eELzbGbDCK4hQu1IJQKQJ4mkm29vrH
39sLqUAnJQUEAH1imzsXKZITLKdTRYoezqGy4QcEkKNTVGqOcnXvzCfY2p3RPhcoqUhBK81LcGm6
c0yiPCmY0BTGWgxeDOF9CgjmpGnqys0d00AsyJuDSfelrPfQL5s6YDXRLerru5++etQthmc7MxuZ
3y3Ti/0+tlwkGwSkUfB/QmBea4d0IceXbMxYrsuxOdK31VD+eYTQG1Dpqm/6QFRPZwxif49S4vyV
tVcLA0MnRxthhMpjqoKp7iPVczWZvxxAp0JCQxX48kH88ZhY1V7Q1IXT9jWt5HNVjqm3NjmHDk8F
AcIsKMFo+BieZJ8P1EIws6JUrW5hJZHFGGKBKOLEEShHE6I5WKFjeM8bheclsuaTAR1nLLhYP39C
asRKGGVe9uWCmvMMj30GjowqHGgywCL5YSQAx29nKoYh6JehQJSwxe6YPoCzDDRGcyqW3GRPY+kY
dpdLPeU36yu0jd1hzK20T/ROM5XgjceZadKfz3JffJaf1aO3zyUrFvHZsJTLfBs97fOoMSjYnudV
9ocjLR1POanKTTXA1UrNdnHUf7Sq2bdJ3hby1QUbA4SD1SkW5gMXz8udxolMzMCMzovGCGIrP0dw
Ce7PYBvdbstmsJBJedW64Vu7zNA04HFkorRki6jBY41ZmVfc9+9XVFP9nVBsMKtoi+vX+eY39kGW
P1j0fj0dGeQODY/Gnwe+0VynbQGJJRC4hePQu8559Pv/CmgcvXVFZepVRRrT4AZzUWxLPvQchJAQ
Yk5wLj5J3+82jXpaYfm5UfygIotr0BpWAWGBmuWPDSj6xrYSwtkHhJl7QJvDbtxvAo9Y8O9nS9rF
eCUBjSiCaou5m2THMT/f6GaL0MAHJTNOPvLw9olxhzRpkfymIGe9mYGSasbBWGdH0V/7ar5C1Jp7
+Fln6WXiQw0xWSGoPu4aT6r34DwRcg5YNdsCox0fZi6tBZUw8kt9Oxb5iGaj8UAwCSY7CoqO/Ace
WXMzwULcs7yP5L6pMM3pRY/LhQtG9bs3BcQg1wXkD0KeLB5CULxmWNZRdnWsibxKhKun7wN6rM0E
1/grBm6rcYIbExpdmM9Eb8myzEbv8sBelM43e41zFaFjXuAaUSW9Q7qI/NdzcGOIT4BWql2e9UhC
6J6BXeWUvdjKGUGHUy37E11pqsf8xLTbX1f5DVxsrsvWFtRsIJwPbSHTzEMG1UjUw3XW/hzD3I1Y
NmISZ0f3oPdhLFsFsT+TjNISTK4An79T7vMcGxxEvX8g2ZyytFs3MeGda5K6FzEWLGjHxVyBME39
APV0POBEYcWni5mOdZqtbJtRVS6NSOolFMSNsJheRJnvwHWhTErLEayXfd47lhgXRUmNhYvS5MwZ
Rch5Oy7n8vTJr1RpLsZx/IUuaJD2x0www/3FYR5XoOkWRptbXl5P5aR6msTlGIvHM2/5nvB2xCvt
PIvBvWnHfYrYyR0tXfHfs3ZWuJZjwedWHiz1OK68OfhM/G+houLg90TLcfRp4C3+JANfi2866E0B
tIIXruGVrDypS2LT44cP2PcQDNzyDLzdf16UMyYK1DEMpavPnpUHibJj43/cR4mbcSA0uyQOv75I
gBSm55sC9gGypxOmr3FYhEsrBtVJA4B/r8Y525MBhZUvWtYi0rsUVwEfdAcmoKk4mfKiORWFUTr0
roljlRGOqcGtcNDUJyVyifUPEBB8Fxeig4tu5n9K3xsdwKcvS6F8l57lwoRGqoS7daoMqqiELmUD
DrtXjjoGNegManVyosbHVViHyx905Bl0qRzI2xcY0v2kjFJdYfNmlo7rrJW2spxBQEtsYFdJcZcr
5BkBLUYwFR5KurBOWhJ2cAehPm6hNldgA+Xp2mknuV0hcqT7dCt6Dkv07RhGePfSE4Go19WnMSFE
h1tURqRZ4SFCzJVjIVsYMijft4NA66o3OZSXEdFAozdk+T37T+OiZWd80p/l0ksROirhVfYp89nf
7dgEd0XjsHhHdwnkXd1XQsgcFB91Lo1SYNtX5NYpfzwii3/yCpvDkBWLKuzX8uFpeJjK+c6rm1mN
946+Rgi/2mYwhijCxE2EVBRuryXVplclg7xHW+jAkAdREOO9pKdouo1a+obVrE7G1ufgjvJZQQAZ
Xs2C3VvWAKDDZbTiR5LlanNoN4LdsLkELnNuKEFOw8KE7B9DBGJuZbQtiOCEjI6A9xQYXto1TbVO
3WOSrF8C+Ym3A1wKTbj/ITTO65ed8yuHHeyXudrFXkTKv0pimPLN8R2WbJjMvldNFFZwnLAMn7g7
+voqPB37/LK1Cl+FCXSRMXd824VlrcmElVL1RupfLsD7Wly3nJzvjYY1SGXWVYV3D+Kxaoeozznx
jZsstUeZmZiSLAjQnVttNjE92fVhskT30uOO5uBs+cwP/o7zCftlScqRNBC9JUIibYMu4uB6NB63
INu9LDyaQOvuf1gLz/2UUSr/ekIuhRiEfpaox79S0ULHZx7TLejwH7Bps4sb56nPYB0CJhAvVQuW
VHLjMFgMSRe8bxBUTKWQebecocrSMmHPpHLkpvm97IhL/pgBiUtYIwKN04U1XGu9UYlyjf4OV/xw
+TyVoX+35NDbP4dmZhUvQd8evO3yt8xAjs/c1NRMOAbwoKy3fv/3qwGFrLk2xfy3Fdk/X98Y9ObI
w63XD6kWdIAGT181WTZ3qKcspYsONZcMxLGtqSFEIZV2aqN5g75/oMiWuZIMVSUeZvDwcmpEFJGE
xm9tyEtWF7z4Yb4rxUIWkaII23M7jSKQqim+3INGGazloWjYbI1yM2YMWs5EzzrxC1gboHH9Avn+
nBfAFwzIrBdthkiEIMl78N9EzbubmcJt6bRdQ2/Htv9NXieb6g8WOymSPOJwBo42jxTInEy1e5UM
itEf5Sjf0fSPUZQ8v1AOBvOopqUCunj3zr8YLcF/HxzSvUs5PHpeapnSPAvGvytvHGbYKuwmXOsn
Mr9S73H/tVJPVeCkCY9llkx1cee2yYzzKAqXUATG3SefMZt4S+zL2dvyXYC1YFpjzRNlOLiKnKWP
zRmfyQlH/TeSTd93SfEWrC8fEaHR0um0isrz/gT/4wOLUqoXvFvbIjlF8cG9OXc6rcDulrkFnQh2
C1xeVAkQkSZWAQ+9MhB5n7NDZKWYwW1jLBP33NVwkZrUQj12PgNB7hZmnDcBzKta8n0vagJSnlWR
/LRgNZK7UdQ99N9aSxWtrWsQRvZhrmwoGUvZyXOr9d6h9pD7Pc5M1n4bw/A28lPsKAV8RTjBvpwy
5PJbLu0GjVQrOKfgabZhn059JUeAQcX62REj10YsUcFbkpNNwdN5ZJbwaZmaL+HSsXijKK2KHs33
3xRfEb9100RBGuJHiiCl/jHcodm/eKjgf7niOkS0NWwX7NxRJa+GM6zl8C+pKa0j3erpvufwXI6h
Crg4M4ItgBV2a/ktkQZVr+UWxBYIsGiM396v7uKQH/T5g2+r9WF7nMSchjrjLAFVaVFbapGi8K5K
vF14NQB9vEVvsdglG6vzHKgaJX9Ag61HQfj2oBv+FEdOZtr60ucZtr/u52f12bp02fwcUxC3u+t3
qPgiN0+vBLmMGkO1KLRQ2YeQyDdT+6A5mY2mV7SaOGFkFYSWC0PArEImpKG9HW+iM95dOfZt7dNk
E3PIDxJIvka+/qrUF+ncvmsUCthW2AxZ+SOJERTn/e4l0F+bG4CmXPEt7DbXiIGpg+8uMUW10POD
p7TTD6NNL0wYVe6Yz3eNqBo9NjmwwJPme3w+rqDrLLevMqCIZJUmsv3qfKAFiTT+mR4cjQDFGDa7
mK1dgYSvu2rOryq2eAiMUwscEfgf/dMYmzkyfiNZH5yOOxNjLqE39m+B3tTkHJZMvybFZq9V4mcg
zGe9fJjdqzH9PFSVqiTp0q+Q+ff4jSH7azef6cZSgEZ4syMFjMUmZIv9wLEiqaCiw4sLJvltqsVI
hveY49qhjBhANk3OeAk+f3+0wNc9mecODMWx1W7h7ujIhVb3ytVJprHa4J/vV+uq+dxkEAL5PL3N
kSfmYNl1UoEA6mpLo7Tt6+hHjdK5sAtoEw8NrWiQWpfmDtgDOEi9n5PNCZ++UZKu5bA4qdJbkRqP
J1CHbWkYLb5tQ6XJyW2jVPShd6tVlgxb7VcQSZXE1RP+QX53mo54epAFGzrNK1+WNlt/xwd5Gcme
1c2gBfQwc9KgUqTiozfg5sA5HB4JqjafrzN7NQN1iB4XdgSso7vVh81qTJuasrTWOBvN7QbC32A8
c5t+PCBgGAsPycoPHqsgfDhq6v7g8HTDvMURT1dL9SilrIzIHApb6xtikzaeJL6bnxLHxRPakY5l
M6H/0o7OEaQf2i5vO0MnOIc1dxxu7Bf8ZgSpyJkLMPxHTx6k+AZIx8c7VurNK6IoeG/4KcE+yy93
yWRrc08rzWMWu3SeTXjVItlSHPEsWyM2SzPs9DaqLt0uUSHlwsGwkSDNPnRKMaBjaPRHijdfkQci
xGl5tWwQA9QdCMQbO2t7wPJqOtx2+K+XnR6XYErcKWTNzEJ8RBV9z5YscPEDIJg6V7Cb6WHcfpS4
9aYP5vsMen/TTjoY34KUKLVpl/JkB2nO2qWjLqpYC1xSkr2VKtsibQXue4+MyYI1Fk0krWHuyeYE
yVyRFdyKP5iNaqCLsarfbkB98CDHJLfxmwCl07O9FJwL42MpdOIsY+dML51mJyozn0Jeorsx+fez
Ua/0RYYmgcck6myHHQwiMMTSNBzdeUU2cjgbWopFKRMjNwcw8ZQKHj70Sv9UVLdauBTkJMx6V4Sy
mRCGXNMnTTg+Vg8pBM9PSk/x0kufTN1PWVxUYySn//d//9+nSqGDwRCyzcaq6qYrmi/ZusktaJ2I
I7wiV0dNxAg7hJteRer1ZtamxENSqdIs/oFAi4V/Ryc0Vt9PLCqxCWBKCDS4f0EIF+oOWRLMVJ2J
OiFZk6o9xB0AOQMz1r2QXcawQ4nhOHDsCiEiKIc04ZijOQf9a2y2cOJgYUx/kxsfpu2Y95bh/oI2
exxF3XT/EzPp2/tJULjB7uC2Lc2ESIbO2v0IcrJq9J74nymAut05rMHdigC3RVxlSiiVc3Wk2T7i
dhYIdsRfATJvnLG10LEQMn/DmSh1g2QECW3DusG1Mf4lJKmMRNAezpXhq4xVu/JDLMEvC52Z80Vb
XK+gVvr5+rkLXco05niLVhYzjX4gnqaDDWZVTNBSieM+xTAVhCtSoX2zqzTM6G9E4Wolj89E4eSz
xLIGHn5safn44z+olkdHx3YcQOGTBcns3yBSGzHKXG/Im7mDtN+FNrKVfKcPpaVczZQLUMOZ5C6N
2IlnjskmraC1xwZ0UdvGGMJPwlgFJ+p9vb5XBf0WIvgENh4R33lCWTKiotL0gT49C8LOdVxl4z7I
JdXZHXxFz32nez9G0gtBvXfqUjXqkwDijdBmsPAlmslqFwFcKtubBIm/y9pCS8hi+PdYygg+KofA
5RQHPnYJHE/sGvPpzfQsGPH5S8bUW5NSJT0D2gPOCDE5QtQaf7BvGGCM2u67Oq2ewBj5U5aRchbD
cbizuYpT/QDE9AgieMSqcEmK8IZNVIBicaXpdEG5N7zEV4LDecv46xTK4n+hkPKc0AOFab+Roqs9
qei6mKja3EMK6TJkWkZxmlAcOMIORddsG/PYyIetMO962Q4WOqxPhM+yvgFrxrQPiv5f3p9IoP9g
bBScJpuqyWbJ94wf09uk/tguoAOV0w24Q4iaetdxE7/Ppqvln5UtHCaJ0j5zpqCmOYR5G3w2Mgfc
tnV0qlWfp/OCjuVorptLFB6sYLvVNHMzT2PQU/Z7FYqdMAiEtN8bURPQNuEP2N/y1qAhmc+p0cB+
/oRX2pNDEol4/Lalc6A7Z/hr50qhkymIJxyx4ou1M8YS8K5ET8OZgrHe0gorun90it33PxkS+Mbq
56ngRjY5rWPzM+DP7u/jY3JIn3kBhgnFa/QAfvDDTKAPtcr8qbS0vbG8RDXSWTKzKKs7ensNeHbi
SS6WDxcBlrraapnKkQf+3ZSOJSpRTuiRstkdYH5liriPeLUH0kMd90BUB1xb5dGNdMTAkh8Vk24s
jxqdbF7dEmvi8nekKZ+RORfEoXtAp1DUWY27p5rBM+u+ayP6oLS7LNSso/3sGXSleRgFm8yF+X04
yG57OMyA3QuzBJuPv7f5hBfCRjMVRz5MM5QCfaruyhUUZSmsMgQ5+rGTW35uRhhcw++Pk0Wid/9l
AiDo9p9PpFWDl0ahJqBHxWZC9a1sgwMBACOCd0SIZ+zI5deVgv+FYqPCopxAKYe5EHPq25lSSnVg
Bxd+c/LPsX/m94C1oZY9zkH4GY5Xh0EJ5HJl85P6vXxRXbyR6k7jy4GTmSzPce9DILLxsrloFtOz
9zY0wNZkpEx3Mf1dcORIVwPsyJgFZtaRU6CnO7dOcLfOCKL1gl52bKCoEYcR2SCN10XOkPdeKyqN
0kzffFGgHcxA2fl8HE9t0xaY6u2IqlNqgXNZ+oKziE9t6TdbgFvoxriaEZRYgSgfBz/QMUDOWzhe
B+jhv4iObBxhfX23PLCj4qQSVQx0b7mz3bpoocMCeSl6J4+5kvyCWIUb/Ko13j+onv6YyM4PSHtm
mlPg1e3lXxCJSo0XsEKu07lAVnam61yVJiidNvhwGvA6S8KHlbYIk/lrZzY6sZjOqm3+OYFers0l
udPBkqCDN05nOhXvaZJB9r31kOLd+w/L3AlYyo310a0E6Z1tqx+octK5rg6zsJzS+/HE4s5uJlVu
GI1naIbJlSuloGtFGG2Gq0RdYkaOtnRljyAiqfKNSl1jvpvspCI0qNHq0CA0ip3UXgjmT4UJaVhE
mjoUhrBOibV96eLwA5eP8T8DGbam3vpojBa0BlgVPsDyNetgvBh/KtQ43k7CeMmsvOzZoGJbVUiw
Y/bhDBpb0waWaIHQWbYWnbXoQ32cyDJmn3nwuG65VMEVT05hQRPOAxQdof9M0pqifFDKm082VMvY
TRbNDnTGKqEQ7N51G0HriC2AK1Kx6sFAL+qleVwFlzi+c0Lgg38dMKgdIF9O6IuTQ67v+TIFMkKb
nO8TFCErXcvD3EerGNnF2G6rLZMqJ7sJnfBLXSmiO7gyob/AhcpI/adhNWmFzIm0U4k9axfk/xDX
WrcXumQHbC4a0+0Up60wHSllXp6GWpXf2fXUna0WC9FoYBJS4iM5D2UR8g5tu0GyQoTIR4nT/bwN
3X2FDRDNkZaj7otaBHp+splExi+wXgNPZbP8lqCSM1Q/DHbFxsvuaQko5J64fGKVurlTrsSXrVME
NrbTxz2oFMbjNphtmSRo55XoMM/9/uPrpE3xo3zF/Gh7q3Gx6hKDILtldvjJBtts792bk3PFwGHl
YSdWRcjUtRMk5VpMIQmNyTFZg0zshrxyVcCp8PA9xveQ0ezMnu48AbBpGRYQJekpx6g6e8g/YZV2
R2I3a5T+ZB6d59zym6IPN41IwcJcnYaFceSCvYjavZsm74duDiSHI6kMSFJ3igLxUgyw+BbHuT+f
hXEj5aCYBBb3fJQKLyhylEDEuS6a+6LIaPhgr5uP7XdaKzlHEMq7nLgjvzoOthRjPkjjIjoSFmxn
kUC4721J3W0ButY+5fQTJ/Wa9hrR1pNOERLvdeHBKdYqTZ8IU06CPqBFUfMpisnCZ9qXL+SYiEo+
96iUe5vBTdoWPhl5nIDUuUpvMpk31NJ3Sg4xWdlpV2ZG4xtDLb2kHvbfFotEFpEMB3GLzyvnuEB8
qTgurWzQSVGu3zxKAhVBuyFcAxdHyhCsxwae+4Jb3gIIMrL+3GjHtU2caL8AjeZjqoj4fVoSFgAE
FA1DvBsBt1j9fk5lPPNT0QSYM2FozypfhLuXWbKe8dGjB0JsnQM+w2Z6h3ZfJ1wYqLNkUanJQCk1
GYOCZI60s7lgPAZboazOBZ2aqawJK4luyzMjLfEWlA2lcqCir+QxBQeeLPkyOuuGFovI8V4Ffi27
KR7JVvn+7Igh9xcMFV0bbwJzCv4H+24SqWXfT0AGuyxKaGPO1PLFtPFNGai09AZMGwTavopmBgC9
Hc3xeKgkFGr+tIy/CUndX8Iu4TpbgG94pEcrJOTo6LOlCE9uMB2sanR7Kn4/8cnqcnfQrhP9UCRs
m9WhrQjWQriCqPLAiR/1Tn7e19fU383W01qF3EVpyNv1yEY6BWnpZz723Sb+wIHtXlrEOQxLz5O2
ea8Ar+BEKzy1lQCpvEm/NNEqsp4YsX7pxyyb9ehqI0jmVDOFIIe9FHbDKUYlEmjAWN+Y1USKmGkR
U7ccBpHt4hCIRvZZXH5MWclHwFW28pTgvegPGXCMwvXzt3I5EqMP3gWVLQ/vnrB4qi2wX0qalrwn
xKsYWkvX8Z/bZgceVD6QJAGuZeidZe8ozU/IGsdN0hkdyj6svAuYphnzSE/8ciYnHXZf79aZh16T
xyWwfJncVB0O7C1kw0CTu7fiRbgQEp4BXuNtkDAWlNOHQG2CB91RQ9rhpKkNB4Ba9XMqVvN/jevH
dvUO5nHw+XNAac5slY3GJqQoGfGNW5xWxeR+HKHNLX+dcZkTPBWGBCRiltfmAsI4AHToNJw2XAMG
pMmFWGAKnZkkRmW/w1ZnVaTkAtjMw5Ws39rrdj1d0bWQ0en3XUpm6KTGx7YZaaE4KrkeFGFIFBI2
j/j0PZNeporaEfCD8yyrWIxXvI/zqX4sSZfij8KxP01s3vkszCrrSVUberZVdAzkjxwvVwtqPN9C
wW6loIVuoGo7eYnNIMKfRTGBbbgLCH34IfSPd6GvPW8R5LCdQONa74EyKqpN4YRZiXZyV9yk2jmv
MXQ1VPQcF6JKdZ3hrrH9v1582x1V+EKARUDL6UbDCWe1YT3BnIz0fQ7cR5DF6vjvIgCAdZdHBrJ+
QmQw+WzVJ/QX4QFDH7u2eKVnsfNpndImLitZ3MQHMF3EKWiOAKJwr2XBgUA6WYF5wxanZatYg0e+
FUbmtZOV88l69j+itdjIKcxQNEfG5n8KJuoCitgufWInY/OIEHSNn2ZyCIm0yyI4cm1936W/dyMy
Da6Je0i8KblSoKvl7QiF5E/g8K2BGfRsg4s7grQpD23xMvyHMVJYSHLMhkStgf8roEtNmCaN7xHZ
Ou8wIfeHKEJbhTHj1DiBBI9zmY5zLSJsnDQ5HAD3/DiGkpF37/2IkDlSrOu/M5BFMXvR7jYIQi9o
zoAj6lAIlfVsbsRFDbnAJMNDV67X5Y5Gz5zrcMSVgQCrsAcKzNdrTRMaXBuXGuq4njfCo6bctkhJ
pzVoW7NWWe+zSXHqkRvbopKlGox7KqRuUVimR7LPjQhNPDIyeDR8gHetX/KAgL09W2ki3/TgcjMo
1TI+v8Md4Yi0fCx6JeaUC2Jw1pPxNcdNA8PBJGSNy5QpkxIaDxLOfepx3vRkO5NQiYu22i9t2EqL
X8w3gPYjiiGX9zhEr007K0CCWadiQTheWrkePOpchQ0cG63YFuJ1f2epBLFgT7vT6XfZT9Jf6erY
VVQhGltPxMoBHSyT5+kkpvBl1msAxCvDonQMrdSN1NsbEryB3LFK4H4hwkeTNNC1cdnrxl2aR9Vv
7GzahShtWHSS7LTSrTbZtMT+FF2TXF7z+sa86khYaOiZlrMAcan0arLO5rnxerlL9rk3LixdTIwV
34WP9ed2fxjsA23xBpl2Ms1qRETcRKKgCZXgtors3lMPzvC69q72i6wb2n7i1hzSqaMoHypn44Ng
H06dBkzrqDUcMHfa3Cjv8US3n9VPHwUgzArssXG+tbkDujUYknotYVmo7KP9dB/D5rEvwVjzDQBj
lLIznKMIdsxF8TboYZjFhef/96YKOZCAe5E6CVPI2t3KzHcP1lO7b2uZVyNHLmFyw3vRy4Bm8s8q
fbT/ZqOTQpbsy4s8meBB8AA6IoTJehjnwsLu+FYYx/iNrX/FRz9lIHC3YHqnAmp6nzciuLR/3XpY
O61oQhP01ZlD1UGYsSE2QEHLPlRJVf9mUEPIagvi5svMrifGaw4/h23FXScC6rh21KYkLHz1mnhR
oVnxuuvi4/kEaf9k6o8kFJo6apGHLDhwxSfC02OVziAi2MSadlqpqqhyD2NsAcRP4gboI+v6cv24
D9dHbomdMnVjyFwnOt0CAixZT1vx9vjVvfE7fozwEfghVgKXTjQUcn+YlSa3XsSKMuhlLqGH10UF
ouf7TpKw0o11ryz32pW4EQ0FGYwHNTHCgMNyBHOPJMBW2WcnKy3U10+ZEva1angTib33U3Jv0Er5
NKOpX625/yQy6jl+nS7KEoy8SVNFeaJ5RyfKVobTSuP84/ViNYvJtjMffYGST2N8erf8MnOMsgSI
eemVaYDt7TM0bHT2gqi5lnfwXftAJZd/UeNmZE0b9afVzC30V1/8HsB4XSL1X4PbPjr2HkTSXzVl
IAxDg89LedEpHGZaok4Twr+SzsXAZSml0izrvY91QpdNcx864g1Fvn5yzwfQvYs4JeXqMQarB/D9
Lfid7y76SZ3uAX2jYP1Z2ZHHNdnsQoz44LzfrSFjV2yfixFaSa+rBtLf5IR9rDWfdlei4A5DlH0l
CC976Gz6XP+UJT5NhzI/Wrht0jt+cmzc9LAWbS7WBZ3a56QzW6JtupXVkZvhGttTV3ghcWhiX68T
fwF5u9UwtjyP8TElFn2IsTzq9RcygAKEZ/MDBeiVRxH3womYJ9Hp9s3Z6RPVBtS6SW6e6iYAoG8M
B6tpmfqEBctbmjfA3RkHPe42mMjUuhSmGoB04E2XAK8G/DA7+zZZB8X+bcSKe9Iw3OlF8V05WHIn
krS7vTJq+g1p509KowJEROT3m/o3jEsNwNK3tCHl3IUJt6PQQDkdFsEs/4mOdMsmRrUFqBI/CzRP
2AEuXmFG2dX6kRG5C69rsIAxrM0kkzQJvfSrF1P29mAgGri/7VSwanVh4Qt93Y+UHWZA1RDLi0Cm
o8WZikNcAFtaOUZcmkQOhm37vG7rGV3Oyel7OP/qj/3F90eEOaWUKFtXKZRvUbIqY3ikwrTZzK2r
4vJKSQe5sNMAtUsCEx9bgRS77IQuKsCMPpUfH23V4/EqySImUie5KC8MeV/Afh1tcxxLKEVOH9ni
Ff7i4iZaSxJn8i7pvyaoCo5oeay1FbrQkYNvqchd+1xK2EGuSkIB1ovfx3t6Kn3s3qee5BFe/EB9
EQONYJlwBbAyZmjVz01SgTn7vd+87oj7KvdQ06un/fAM5S8+HGCQR/QEEvznwh7059z9yohtTnxV
pLwFIZZtbwWlxj61HmpFF4Ot7oiOJOhG+kFdK2ER/iFWpWbEWfyoxpMh8RbcECR1AdzEQBqGzkYF
C1v9ydC0IBUHuPWDcbN8D0CFEnLzwaVy8Imo6abGqq7AUOwRnWQrgx5tO37/5aTpE+FZCjBvYu+F
AJFQxWH8HOA2w9Nx/FsCeCwpDv+67ri56xjfAUuMjQSXMtwn23Z0FeLqfeKktnNoTSQHwmj/sgRj
DANBN9AKhYF3nQH6p9mcXDF8rZXy/eauqrE9MLqFUUPNG5NTwXtfgYqv+Irp0IiwS64SIi0TgHcP
IVLT0a6YmjUepvqZAQSQWaUhUUesronrlU7h9pr3XNrSWyLQGaM7HzGyrfbAwFQ0+Bwmg0T/+tcM
k3H9i2GM8Gs0zyp9NmCLbijhnaYuQP2JZQbUq/fQgRbb9HnfnJiQOeuZNMJGPFgTsVdVuapsVK1z
y63e3vtX1xyi9ZrpYKvQrmvbuCXfKFJQTjDoTPlHqNbHUgqxGZVWvs0TtgDtLpIEuSPKpiEv1DQo
1yKvZIoOQ8Rg5Yu4Z5doPPp/xTf0tGepbuz1qvC8EYvjlMcREiTIPPb7JU1LL7rnrL4hENAwKz4V
l9mTIBLwKuuejmj+7f0TQFz2ekKPRewIzo/s3I79+N+iNDFYRd6rr6w6/LdsLgaEF72R8BVI9KVD
msqfskIILnIXOzAtR+DGezqSROtUVzUKlZceoKZp2lqQO7zV22VWM66Cj2eVu4ppWcap3+NTvOUL
dP/Oley0kuHq0AAwKuhuFPeP5H/YwxqPA58noILr+NNGVubDikQuWPRIY0BUw2I6n4v4sXaIgX36
oSN1uEJZSm9/5TOX/hFUkTa0qhK4DY6wHr1vW+avY6m0UTq2+x1FLf1FWL1AwQVy7tHS4mToBUVm
Wk/f7k5EOr5WsvWktCkOlBe/vg+VczqBLgEDGKTOcYQIQriDLWNCGzxlzVkYnWWv8zMr2DAMKR9t
NCyyZfrzOvdk0ZjbShNfbgty4BNuOtzH4UYkqJ9sth8q90eprsxR5t6P/RWYOy8QMpOpftjRk7+w
aSbVmirNNaSbgER2208kgVmLTbxS82+YPvUDPK+ANTP4ufyZwLZJAj2QqumuTKxz5hLh2+NofVJu
hyabcuz0YeZj9hpM1NI7mGKuOefojYZz8BHpbAbM1Vwrqu5FernERhC11QDZfJ7rTMMHyyrbsnZh
AFqeQ+XoRRC2UnrJHIZ02nkBd5tGEEJBBBhdudLO+HI4b+XOewU7A3RuTQsIk8Uoez5IApkUKBto
Th1u38QIgqb8k6ORqinrOOOAjR67wQ53a3deuWhdXfY7rjv7BizDFobWQ5dtNLL5ewCVZJyAl1Ax
6bp5vJ60soPXhzYJda784e9WEPYWN2wqHTbO2xTiP52gyGW6jbYHZx2Q2xnAps4EdEo1kGXta/wW
XUWYASOZ+fIeDwybb6uC9zbhvhq2MvXKI4ZjfEmuDeRYVXkNneURbnMCqCOe3PM1AnGwlf9YafGG
wSvwQ+JfWR+ISGgX5rrfkxaN3oSCy67jY3oqJXtcnP37mbW5+1Gl6IqpOulwiv020wCylLOh/38B
3MQRKSG7u7MkdjIM5Gy3zilBqLkS6+E/Csm8poBwYX5rf9tGk5TBhVINXjUEm+Um8pFSaAAX7ClI
ZnijkEc3IF0w3IUqpZJHZurzrzC7D41Biwaos89qHpBSYvTIFqd8IfyWzc2C/AtoRzh2nvWjCnFV
VWfjg+mWr1ty2RsB2tTmP7PS8bqdPdUbULa1FVVIvh0hSTs5hyEpm/W4WJvMznCeNoCXax0aoR60
NqiGmzMrsNt/CYtPmllHOKdoUmfq0ARtc2qNS/4UD5bZgDRGdF4TmErDSEJu27OCNByp8Rb8JDPt
RT+NMacC9vUmTROKRnmcZhte+lQajjtSsL/KYksQNCDiOwSYQF6H3/h1Mh8vrWxLO9LIjNLoofN4
dljrhh8i3s735cSyIWFUKIvaU9s4wY6l7wu/NV52Bp121/0QIiK6iWofbSFGl2VjIsAJwI71F5pq
9CrDz+PDr7qWci8W8pmzQ3ee2VgadOCQApHo54gTX++yT3hIFX566BG+X3vQ09eO669IjpIt05XJ
owhHlr8a7IypI36NsbiO7A/buu0Cwe1gtQoCxTCSt/io9A1otgwPKzOzPsc4telpqJB3DWulfMId
UZ7XOjAGM5NXnp8pZMj8NyFofZAWRwc6Y6oDSfTFz561fIVGT3fa4N9F7Kgol+ssvkpGJdUUec2g
2KGRpgJPTOO9hKzK2Xp1xxMXwAPjAy8pDx4TV/UU46Kxuxtk6nLuY8R6/pYn5CFz/BDfNI/sCp1O
76ZjN7/3KloIfNhJ3u5TldyrBPkrv0MQE7J2E+PyACuklNI71vfu2ppKfQ6im0BTIWq0G5ewWQQL
anxXVpkRwnOw9BIlspjMY3ymSCHZsWBNrFfqYlUNCvddFbMirf8LJs3S4FAoFWVSOZ54AIO+UdwU
XKqSiXbgwpge9gx8909eoykIllsR/Tmy+d36nBP3nRiFVdk0L8d6x/nWw31Wuy5EESUu0CKCu0qu
B9KOb2Sb+6x48pcCw9T8p18TkCRE8o8D5YQuxLYmGIKMfJQ/JiCORV/QPGQJ/7ZgvqhUVZqvYg51
iOHzbotZP+XbzTZy9bi7lv5pK6BC5pfwd1TQRJCfSXv0P6lBvPnBcNmmN8y8MG3erGhJIAqcKFud
gHHGdTtVXrHPRN7S+e4hLHdM8KvTKjwHUzBhHOUEFWwyxkKp5aXsn2MhRpN41u2V2OBsqrooSmi0
ycSlqb/7rKrlpGWi/kKX/P8vo4T4cs/qx9dMeg5KzI6GbHepv+qd/G9iRLU0ZFtqhiifKVzfXpQ/
J7+yaq7yxHRasExCjVqI+N3izspLroGSIrp1aMt/M00/Bb4tPKZrV3moY21KohDndFQzvqFX41WR
+Jc6M7OkloNWKlN+3qF3GNXWSTwCjWh5RD4jIIcOLQtPFbeYfYPp18F/gGFbJjqJQ7PkPvjPI6Mx
87L4upAVNLc2Ko0FOZEqe/X1A69phxdfbPvzXqTYZwPbCzeWaFVtR0pwcSY2qISBH3+CtAaR1bEi
eeT0QTdmVbFG4E2tWnVgIxKd03k90StlJ5JUWyO/dOQ2J/laQkAz/1L/9VO0vVLHyPcPMDqB+t5q
iN2XgYadAHDZy/rb8sPxSaLzq8w9Gmkq7Kp35NT1OqoTFZ2C0QfIITCAgte1ePt6hSlqlruLgHJU
PV2pRTtcHwPNMdDiA5v2kKyEKkrGYNSel87Jbl+c5kRzVV/HE+2AuywMCdC4TIaxrfhYR41Yzm89
7zVzcfxgIS4ZqzNBnQP/QKGS+Yk9rD0ry8/5XMHHCp1KrAjQQjIr6PyC2VlOxntWg/0TwksghVmw
pjqci5CW5RgWXVF2W5rk0cAKt/GGyzm5cZM5TxUhKtlGoXVeTlOx8zHtL4IQKhSClUmYdp/4G2Ns
0oThY2PLkJZ/jy5yjTyarrrV2OFV4HzveE04lHbu9pWA842RWWqaS6bndAc0M0ohj4WKL4jPXYuH
w69AJn8QneDWiMGD2hf4xZE5l/wQmTI0vwuF5hM3WRoj7L2NCm0k8Wu3MUIRJwWn5ESEVSO7U5sL
l471yLIT7ANj972SLz9oxnNaVYNWE1sTT+zCmP9BhGTr5slzJUk2cOQLhh80dCGAzmAnJIazU2uk
cR2FQdXRlq45teYkLKiKUBlP0B+DqFEFXtchXv+2IpDX7lBVL1+4Hv6evBlGUeEExTcSYIBx9HlE
P8Wa79Pdsu1A3+A0QYqtHl5xhsSo/twyowrEEQy/G0K+FI6JXd9ItVKGzuZekrkhwQ6OBym0MXEh
iMnIjBRfgUHhC9J1ybMkWw19r7Hh1u1E87k+L68JbqCMNwbGqnmKm4TInObBfAvVW75Gp3kEvBhE
K3FUg2A/SDz+E8TttdO5ypVDwIPhsv45L6MBFyg3Df20ElsmynnPju5OIUrUILLcDeTnOtwdXYnu
NW3NZGrGN3LmzpK568aMO9zvKV7TbaKPjBj8vKY2zlQyHNCLGGk56U9QsoMjUWKyLho2y8Y3lLNL
+xJW5Gus8WBO3cwuapU19WhEfRf3PmX2V4b8l6G8H4lZe32r+2zm2AaYeNqGWuZy3h5P16sp2pXg
7ebJSGsztqDNzBdet2UcnJUaqoqO92aPxFBfV+br2b+2jpdcGGqXU9YaTSu+aDTNkFRWbh54zqup
+xb1SMzWE8GMQ4iw85RaJjZ6Ra3E4jdZ0AkwoPRhjZ3VPCeyL3uEGskLvtpABKQ//7hLJJiRGRui
QtXMV2zC1anNwsAsydblkIJOtFJglBXOdjcsyS+h/wHWnjs5ZE2Ukwk6UinbYy+YkG7ryq3HQY79
u6bEJbX4BGGsoLBOOujddwODeoO7AbzrlPsbJgUZWLb6FsAq7zWva7uwDa1TwhU65vw04DDFcQA3
G8RSHc7GYnSnBJ2MSVQOWLrOga96C8BoiSjqWFzPqIsb3cyynohnazPLIPf7FjIek16iSnLBh7RW
1BTlE+lj0xfBRiVCkbinUCPezDj4+Fx+WweKGqNAf9+CYKdFwkxPBBkqYW1/KlnmpGCSAn2OfVEK
RNBrwDUGGqzZhdKZ85Au/GN1x5TFXEm+cpxYg3OY5pB0R3yv+dDq8ViNVRPm7Vtlcxm7gLA8zXw1
fJfdXwOX7o+4YXzsMJ+B8fiwdIYmI9BjPy4aL/CXSSyTt28+YU2wpDn2GTMBs8J1I1pTv7dmV9/s
RVQPJQuQHt97zmUPoi82veOQz50KHhIwHwWsrcE9LPFEdBcgdJPazKLNdnI8RYCKwCXodDTTDz/2
g9x3/kL9B0KYyt7em6JONqVJxIf62uytVxKs1pIKhuKPmf3daNsc629Reuiv4uMwCJYPyRpw5g0h
TvmEojK+q5ryfQrLDju8G7JqAPCwmHNdDhjIfJcs7Mk23SfsCc0VEuiGgzuJ1S47z9SJPgHlj+i8
Uq1h67/c6Oyuu0VS/TUcBol+8RDwDTQ2faxYGJZ9NrNqrA9DXbf3blo/L4+lUqz174XB48/6g60s
1qfflbkBMAn4XE0Fbhpv7OA2MxbLPmQD6i0zHOBRoQ7aT9b58WtZgJneAUvF0bhfzTTv2t650Vy6
2tIMrhskUmZquike9k5jINQes9ZtEtzadZ/p9UG73d/XO8BaHQL5KYQDVuD7c12J7M6nHZVVvu9i
v84KXPymGmgD5PFxo8QN3BybICY4Q2RCNx/kimgwacJtdPYGhldAqYt7BCSFSpyCSpSGdNUeDkrn
wimImZhmL6QXaRqu8oEB/g0ZCgBcCVsaJOR6lvAkDyuY8oBoIo0z/ujxpvouVcuTBqaHZFIlyjsT
6i5/bjX4+YR20ihIJ2NycEidJMGSZU3gGqcSoLeWRPQCM/OkoIZpXTEQARKSA8IsQh+Y81FBZAKV
vO8HGfwOlPzh7JUOsDgKjjiXVlU52HiJXzVigkJH5+351/DArP3TCb7HsAqRKgtgh75Px6s0pEVF
C/cOFq3dI9CV62wmVT3+St6EV9YVOGdH7Wkcz4IFigyLsJ81CXFWEEUH3w7yumzd8E2jH35E2mDS
F5k0XQog80WI2y9VskhCQTMLetUE4MOMMWTWguYxb173Ev2e55AGlK1tNOQP/knyUr7nhOcrhrCy
WttIoSUTUnZj3+CshEjziBKfczeAgrgC2p4pI/gdm2wzYfQ6etiKK4pLsEbYBJKhIlR9pab5GAoo
gO+qdqnoH1t/FnkBdD1c7ifYMbdz8xLFBzhzDQLC3/xk6dgXV3bY7Qra9IqS59dIoVboD7GiCMG/
91RPNMPLzqls8w4HXcfoP2J3rglovEw1Tin8HHAMmiY7rHuu3pCYIIbd+ICHcnX9QOHUWKtuGN86
C0B66aAVl8IDVePaW0Fs7KUfNJb/RADeBnHsBy0Ja0vAS3+0+bg2Z0TuYRwngnLecfBz/Q06WDTV
LdClgP/OP72NM6w/UYErb/w4AZJBXLK02r9Wzr3Hl81nLEQn5LLtXM6Rvb4V+1Zzi+DeTKwjWaMT
IQ666XlUEe/8vWNp2lVIgKvQ1mwxxYSJuRoxioUAKodBs4wjsPzOafM/kysK2A9UJ5DVcBWx5DA9
GsP/BJcxB0M3XBbBQ9EAvH8yNSGkHYyRRu3HR2V0lm8igiSVT1hItEDrZt0d/BaeL13vdXnKstMy
APYuGRqfymM7RNNfNvP1QClPgnMfLRTHzzfMxqEMlyj+/jStq9ZiEPP1l4WDvkGciHzzZkzmoSCb
yIgnDhWTj1Zuwsl7grhWtOT9MnCFwE7jx9CJJFF0JJs9bdtuAqZXJofgCaPj93Qwu8lP+k0J2Gk5
Bhyyh2N6TxcDwAuL+CWonVgS4zxXuGzn85zRmGrRe/MF3CidFvddWlmcNfgZ4dI6w81pHqu7iBKL
WkF3Mzb4wfHa+znING7DFQO4r6uJSCypiSkNG4CHUKKv9oRvxUn3PXNJPC+LLrnvQCpRKM/tXUlw
qY1ln/SIrKv0exwqLk0C9Z8G3mOAIe58M/YtWZyzSADQr+fHYO/SvrA/Y+3BDRxK8vYjXeNjsdk2
OqjpkjsgK6SGRLPN0Wze9hibMj3o6m9Hgx+vKVMF8rtayN2C2PGw5QkQf5RAY49Q7U9aNGqPDuYd
W0OttdKEN6UlXib+tvxpE4uMI9N1h124l8h5OeFEQPicL7AfEJ/w0aWQjsZlfBECLYYiU6kaGZQY
s+d2/kJeHokDZnmZwUwyC7jxCD0fb/LO0bsqmu2MxlgPTq5KyPAaWNuVn8whiBQs+lFDbn8GSM7w
zbkaNeB5pcCMmtamPwBBfWBb6s5a8UipD9U/bWXo37kiEAE8Lj22ccgr8L51HnZf770V/KIikayR
58JjhAYl5Yer5u6kADLsFF90XY7kVAGPRDXQx6S14kuS18sOYW0ke0lIPfr9/CRzgGRrM0uKO6+A
HvXVmN1IyyEAdyD5ITfqbXk3n2qS5ZYjLZy2sTALyvli4vIGXJCael32AJDjy+O9h6cxqGzUWQEU
ZZOyQJP1WYnT8jgAjlfkwAYU7+7tPGvASQ+gdiv2eG2gXE2nb6He4A6veesQztUFTnwHi7F2WcYG
sPD7HsR5/CB5gTb12/+moPlMwOxHhoA8R3YdbN6f+b4nee3mKEK1NoN8R8Yd0cblj8+Q1/64zKg3
IcyjrfY3y8ZxGBqxOmyqdIhMTAgubWxS53Ej3/mR5IC/NHUO5AFdVPzacrLXwVPMSAuXd/2DMwxQ
f3pWEQI8h95R4TPL2ZlzvgNUWOdD7B+QkMX1G8ZMbPaSSy1x4rWKG4r5vsWWIVn6nJhxSOtyETrS
XN8HtB45sooCFJJ1vYPe8O0DJpAKxORmjovyekrc6AWcY4uXt8QgTZ0N8NZWp4y49b3D2Imujvaq
aC7HkQkV0kYoztjmm+RE3IlIYfIdzRE/7JK0wfuSZdIak6CGpPRrWy3Eq6j18ALXJn+z8ntCexz3
bRBSwWVC+AZOlEczJCVtOvJcvL26dN5TTCjywczecUyzHf59cqVxrw27Sev8Hqol/TTZdwn4FpkH
woIO4zEHt/2BIxXNG1ElfIyHSQywyz0kGbEQXZXbcpqOEE9eKiAvbsOnEohzN8pKlhRe7oNaOrB6
7tYDpA/LguCNTg4c6diBQt+vcJiPKs9KaISBzLZsAR1qIjoGuRrfYw+rPWjVQ/K4jSjGkC4xve7j
FWnZ4WKVKDaiDphyJijSMg7b+49Q5yTnjde0qQgAk706p+7lVHbnkD6N+0d5r3UgklT3BPmEhfKB
R3mUynPUcVEL0441JSbKD/S405powE87GJ3uVY5tx3BMByPVHP+qW48eq5Hk0tBydWla1H2N0FIQ
s4+XvtfW9qIytSbT7GdvD6l/NrmyvjNS5uecSUaYKQbxIGIETCcZXXEQFkdXpG/yHQO99QI/kO0n
iUnU3mJa936aYTwrO0etUS//M0q3QbM8zQdin6ghvsnOtM8yZ9Uocggl99vdI8ZB8lRd7q+HYm3r
onXJq2LLCJh+OFqEakIoCjkf6qqYIB/PML6NEF7CJBMcx9YbjGalR+AyXMFHWNIIxAaaTWpabETi
Z0q+MShFwwT+DB4wQWHHWEsF4IX5ihQZUxEnFFzg++3deKPgKpJE1B+TED5zOdoR8s2wdFkCxlwU
XLQ+dfYOKwJp5oLkiJmxPuZSZdiT4zBUcxjqIADINzI694MKOSrcs55f+ie56MvSXbCcDTWwCWqD
840CgpnOP9dCv7GNrHmatI0m3bLdoc9a9V3alNT+0ra28zP/AqyolVOLqV3kQr55KLCoZqd1g4Rd
N5XYMWpajqNiW9nQ8s9c1d+FXitC/9a6+7Ty0tzZA+npRQhFLhHAM+LE8wEKpLMMgjZPGhSxFCSc
L5RtAbaYL0a+5o0E1MCUYGIvgM2oxYGn8H1gq31kiWy2UOP1xlvdbeseFfS5W3DGgDAKnaPPpWtx
0HNDsysgcQnRWIvIJIAjsHj7LfAdvbK8dLW02CSd1nNfuJdBzZsUlCQF+ii5+cVhCwIimlJvqpiV
ZrIvWQGjd+YhPEU5xyzEONjkxFkh3AQtM2YhXvDmopk9Fm2b4fIxauMalmtLqYqTyWK9qLTQ7VcM
ngywlf3Wmp4m8KgCpT7nhTzo4Cud1cDIC9TJfkst6JyeL1WOmnPYST8rMt53blPPn+QWEgffpHPl
cpCsOZm5HeepK6JJoqSlJ1YOINLKCbbdHMqs1rwpYm1bGNLl43wx3Pk9wNGw3RFtpm2nIWuqpKWj
0ZMUwm5CAGyqP8rCv09mLzIaf4u10qEfrbyjvFlQ+VETGXsPVTO24fa0ezqmYm8ZHwfoW/I+sZDA
fcmS46M5599K/LPEL7VAmppRZYUkBCvtbk6G/lcjtEp81wQ7BXcHzbvn+Hvg2iskoMTIpMmn+ZHa
qB8hxdmkE4LVsOZuG2gQTCDSrrYcTQ2UyPjuq2u/YCJwG0k8txLcE92FAjI8ctveT+gm7LrBuZ8G
7D0VVm6N2WOOVxBBGps64nE1e91ix6jambhU9cgb7LTOvFLBiRy9QPBi4EDYLtUnwjc+QRvUA/pI
nECyPddOqsq4CsYGvYS/+mJ0R3YDGwv8oYt0lB0kCGiANuoI3AdWExmj1uHGquBp3PC65ZpjCqjA
f3QXCMBKGebMNxKwBGEilRIoBCQ/o/w99VfkImk1B0AOpFXi2WGL1knjQ54Vb7J9MNJ6nUwOYn24
HAt9+4XpF+Nmie2YQGe9j0Q/Uhwan2ZGIRA6x9f4XIGaVyy4+r4QzHKRwzPS7t9K3bS8is7oWs2Z
p5Z9g5oh8Hieh+nV5I5Xxb8vbSWqjqX1Wr18L2N5+29Vt5O+odN3YP0n3Z3RsqhipJBUhaRlFgGo
iRYGa1/v/46O125ixiEf8r5kHNJPtPRiugg0iMuZByWfqsoM2lV/b2pcdd2GiXcCjOA50bCx4AFZ
zybSw2ymTlx2dJo5SbtXG22HxIWOEiTHvAdcRIecsnIZY8k6/qyCg1kQxeW6igJZbPC6tOkf7Iia
HWI9XiLpIxCVR8Z+T3L5zOK0M0ILXmAxRMD8V+pM6VxbHHMOFQp+o0ppmuKL/SlD5lYjf0vVuDZZ
KYrzAdu5XXZpimh7WX1Y2DaN1kdg7/iPgB/dEQEc4OlAfN1Bmn7KU5r/UjrXhzkExz6W6k1vgy92
xG/rGjcmk7AZ681w3Z/3CKWsxVpBIuFP6dLocQNmjKbw0K/UJ0dZwExuUF+qFFXV6qSmGMuRoFru
gO8yvioyRn2qiyIU6HVSE+1xc8Wd6Vb4S0Upg1mfcc8EYdwxrJUYquQCQeVmYl3kc9WhzsoTTBxq
13Ee/K1W7W9KoqNCyoqTq0977HWARWYRDFw7v8IMeFXmS072CR3/1OYZNlHUeWfSzl/HT+YWM/et
JnfV7RVnc25W7FweWdpeMsoEuNP+PGCOrrESlGpEQXDyhcKA4tuXUux8DzOhZb0lJ9hfSqLIwSI2
rFKtBxcBAZbZYg7AjXWhhI1Qc+RVChyxK4aU7fn3Np3xu1F3FI/02WztCj0L8SjTd6PVkQWll76H
QSCjZ0iaXIwkZvOGLqdmQLgLY74V8P07XYAnviUQi5qXIqjvor2P/OObTsoWEk3+FiNuB4jSfht8
hkjN6oNLpWrtU33j8ylzOI2DYnOlgbJ+k33V4lkdg39L7zOKbsnt5q47ryo4pHCUvrKsSG0R/U2j
DTqbhToeSnPzjkG3xXc9zCVndTvM2fNNMrs3aK6AixouFXHz/dhYt75c5iLQPCUPtEu6uWQwmPiH
syb2MD16iFzQHDXmx6BuPsIvZeqxqLG2VjoCbe/+NQUqaLkD5jDhO3//rETf42zizyHXMk1jpoc2
D+nvFbNWtxZ8/uDUtOtChhGDKryuW6YJSYqqN/Lk8VZdEDF8RLVPBMeAHOL6d4+vXrCl9KENzcma
Z1rxE2wvkyLH6EEmxfkCvWDePOfMIfrRRgHGFcwNegIDn/HHXy/Xb3ful2/dVCvm2wzC0o/WWRY6
ecyK9YKsVaidMqFPSS4XmSrPkV60ZZTA3JFDmVezmqe6tjnmIMtNe8RRvMMcDOjNMaCbP45KeMqm
Kv5HMh2X0svdZWFWEm71GW0gsam95+AFsL+eLeb5ybMrROq4lszUoGNoOiXSTCL6did7BUiP17aT
6wvTplK6YsQrkwKNTIR2/NaTRzBYBI+q3SYZJbLVnv0yQoSWBEArR+CqoalZX0xzvKlb78N6GQmk
wGkLUlpfmHedGOQWHBpMPeVgqV2RptxDjfaKkEdBz0LwBSKOfbzBMFZexhrBDVtMRFly3Lz1Rn85
BEByamke/caP6dz9awS7qGfdXAXbzXC4k4Hy/Zt7OsLfrrLL/HseGNcJ4cNw+SLvRJRMtpcvqpGQ
TGIo4X6QcPGG9j9mjbBiotJ92PUHd7tM1mBJtdIn3cjyn0Iw4+Amq3mEjSaPRse2WaBNmMBhY8ZU
SFpKEcccOBf4RvcnSSfYJRhll3mKtr/erxlHekP2wrNQQChrux9PP34VZHI7654H5BkvGPNlbBpw
t/ZWNAWCDEg7JREHagmRzZfXeLKhpNMoagCg5jcppm8EAM1ehJmdubkfKVmxHbJskct0M5N8x+bA
m0YzR5l76jrg8ysabkRC43DnopwdLAlcihpaPrwPF9fh2XvyKZjeMOdH1MXh/0nMbrPpsYeou7a1
/LpXnzgx2qhpNKjikpn7bMbmPYx30oEOIJ2CJmh5vStHm3RChaJ50YSY7ryNXvNwxlU6IZNdHeLo
eH/60zRVNcYUXNiz3dFGuQ0gWChvCXMcQbYeWTI9yAbxG2iV/gjpx7a8ZqZba55OE80o3OW5bYzG
kHo8XkAxcnFoIAVMYvYTsp81ESL1TGT7qH9duSN2BEeScb4YgRNxXv+5FD6e1PSg8zqUBwS7yNHa
VOce+TKv12c6klxfxZzNOfnLH385FS7Y9YYEI36CoSP+kg2lXjEo2dDf6+GpvncBUFf7Fb+6syiK
t/Zg3BOTGJNb6IFLFRJ3jG1/tYE3a+dzgvrL/eeaYhO1odgj+rZj1XhXb4u7e3cY9Ws4MZF3RhfS
xcNfwMD4PcdBYpIvTxrcqc+mCH0s/4xbLuLv91u8V0jZ2CY9GjiS9zNd4boI1Vx2wCHfJMKAxBad
VjVDUGgDX20HlHkHwBjUsC9CZQNG4p6HBadKw1fno8fuui1uSqA4Dq3Pa2nNJS++OeKilGy/NDcK
7lHdfdMTyTKvS87hhO6xgsCtTeznBYzd1Kav91oqtnCFAKp7yP80oHXFwfesusk5iYGPHPhIXAPR
wxgycZ/J0mGcR9g6bIEHhFuy2ChqbCxEWJGXWEBg0od9msBCbhDEmncCsQ7CQktMQ7R8YO6iaX2D
M97AUDU+fzvj2AyoLcY7lHZ2O2y3cdQrEP7eu6fDdn1vwgIrBp7DbYzkT8DYeB59Nn0ueczXL7YI
3SNfC1UPY5iRLB77TWyS7dZuFynsuwcLUCbqSZ3zLd+c1cgE2OGFRI0prXDxDC+OYeqa+ZbbiEG+
MGibG68x5A9Tl+2d2fZ0NiJtvAoSgYPqr208Tbr0NUzxZTrJEvdHjaPaKfW4mwOSHaMGGxFlzXy9
Ptg+jB0Fp+0DiyKfLd2KXGSbEigngzRxVvhRrsq6DJ7HClhYjKr6329Ac+uYhWDcltpDfpgTGZan
/0MQGtvfDtPW5HZVGNLTZArpYSjCtiWNnboRAjFpc0/u8NBKbNJZyumw3CNO9nwUy4WZzK88NmMD
j9fzMxfOAb7E74nE7GwmLDMvR6JtAzr9EsIbBjCuT9J7y2soRe0SGCzvXNHBVrzG/lWmyfK1bRXI
MiocZRFh4kfwKAOqzHFK2QU9MLo32V7blPV2vzOj8H01FJTFEweIOtjcVbed3d1T510LCrvmT5o5
vXBVx+ILaAbs9r1B/KesH6q6FrePL9RSbzerZU5QHdJtIY1sctQYN3AIJmuRqVGW0VObQJa4mRDa
gzZtx1xIoa9n8YEZSU1b0kRbAxSEVLdCcuxmpYIQoyyVV6Ljq32ddr3IxX75X+8R0YgipzQRAl2s
TGcRpS9UyHGqdFebHf3Pbld7bFn/M/mV/DNwVeC9qj7RsatBOnGN5dhgfmwfrIqmwKT4u9jKWczk
EAVodPm3GFUhA4ylXXQwWN8n2DBXWAhPFg52HNrGymVmV6gF1WjEJQAsr3dcCylWEclMp3WvFLmW
z0rcUM/BW0QwGQy1JU2MLXEF3Yl7Z+N8a1qGEPBGixVAnAKayl6Ac/mwCXYw/Pk5Q7IJZMwDTpFF
6pTwFQVN/+2xz4v58SFPYgaqb6q6OnFX2QFKHTf2j62XltQ7Z+FIvd9aU+Bx2BN9zo6m7FxIXlvN
R2XqhBzN3pTMG3FWs1x8V4EbcJYtaOtphxXAL1IGvGyn3CHgBJrDjMhoNt7+VJr9yZ7Lada5FJvi
l9ZTQjhMYDsmodFW7sy7b4Go4jacrnZj9ZTwvT4M4jRDs63yCAOug4EYGMXLhObh7HxxIpYKmCXZ
1rsjYDQnGSRpp4Iok2VcuPxWCQFaUCR55wa71K3qaaUVEhmk/rNCKgpu40tdJa0L2JZsIZYnH6DV
v3bAo9yen0gNCEiWTNtesjKFM1SC10Dg9nvQZ/zC3kH4Mx/gae2RzPIYbJ8fV/PZTzuCRmf8MINb
9fAYPFfZgHPoSsE8XeShpS4ujkWSaBj5ELK0uXAKqqoUh9aLA6tcg2LaHDr03HcA8EvuDZM5aciL
xGBjKqaYA6RhoFJqsXmF3l2DaRdZKa0XL4TDDcfQOyOWNTbNY5RsGEqzTpwCjCBEAZG17yIup29C
PIx/pKl63jFZUuZsplt16mUjvHtJM143WBDOrEXjtfu2wHGO1lVFqeRcoz3TMxJP84vBermG3cPF
ZXG6o/oKNH0/IBBAQ0eVQkpygeLLGitFv3I40c9E2vFQhn6tw98t33VM2ZU/9F/dRPFHt73p49Yn
kYWr/unxxtQPocxta13akMVM9gPzo0MgCuc4m3DTwfu4gXMjNNBBIiMGYuTecNGr+ak9ScOtWjPa
GgIBkiLeSY46JmlOzk7+y7zHCpgydzeeo13dFYmkbCxlkzsprGhu/jsCBfvz+uOfag1s6sXx6oO7
ue95R1q3AxuliX8Y6DgNBy9QuGPnj8ZhNPOS/PYcMf9KyAY2jshMNT6Wd2/Q7WNjBbqXsJXIWaZ6
szM9ZLPN1BdgYnF51/Kcn2HiT8x+Qen/ok76u2V1e6LH+hv74nLv13MKfFKvoR6vVrKjUc71JhsT
J7cTUQzCih1ukHMLjUOrbHXOk3HPGXcZycmhVPPBf1lNRDOhyw0hbt9NwmtBXfim7A4tjABXDd43
qvFhO+YS1H+i6aeWMP1ONuSk+H/OhQnm4uSN7IEWEw7WiatBmaDSZFE8bX77yR/OgoIGm49E8a7L
FbtkCE7hTyAExv5U+3PJzK6D4KkhWmQsY+ArWzyOaOI+WKDLr8X2nGtxtYbNJ7ykib6INctAvbyd
FtxCHLROBvWNH5xmRSo12fgEQ1QCxycO2kYt1IavGG2+burEkjrMF8hTVBb/Hn+WZTToRpKFany5
bQkDvvntsK0jPlvkR+nydhxy8dJ+HG56zhfKxWVZboi/TI2dyshpsk56d0kX5a++w900clPevULR
p4lhXASft2TDryXjy6+t+3vsd5Z5gcOhGMtWwCoJIMV7r8/42liGSyiAyeRGs8gAMU8SBtVcYhxt
NGNo+NnCffBuAG043/CMb8xGWJxlv7E+oOBGWc7HX1OezjvOHsMOrRd28KBZ5MFV7eCjoz1L+5gZ
NS/YBaozcLNvfrTwu+FX6PXuRY10egR6Y6Cjaq5maIkcle8k3PCwUjz0nzAnh2c9hwWeedz8WUja
idpwj5LwV/BdCfV0Lngpxr8rrAypNM0Nk8mvdQ1m7W1w0N5m7qQrKXDruWTXjD26BUgcupvEfAJ0
OnRe9MVQXaV0GSi89D3BNv17lP8PfB3KmDZ7EybQEBVa+MWKX828B5Ra2QASoPuGLfD7pfq+URAE
bPcZGr8wqQx5ABnuYmDkYzFAzAbiR73ISkCNOLvSjx+4+4SY+5Gl4jYaNTCaloOLvMQ5wQ6Mq7E5
kefnR46Gwwn6t7Dc/ld9G/pA7lk02hP9Kf4mcIDF7dBbKtjEnEsaCnuoHsfEHzG47O+MSLuZ0pfR
mnRHVHmRE9R3q/xvc7ximcg2GBaGFNhLqzE0gOgU1aFQJX7Ewh7rjj6Bp7K8ww9udnADFxghJy1u
FCWoAgliE1Z4Wfq/XJ/tNkqkpzdGf1l3LLOpRKPQyi0q4RGO1BNQz9wrebiStHHli/cxeJWGsyxD
r9DCifEQa7IXdyBHGiy2Kc5+8rU20gfXPMC+rYFFa3PHWdOcQoejOH0SktrdcVuwKSibWK2GOYmL
6BMba1OT4bY5F4NzacfpwsiHnevauqsmpWHM5WNJ7hurx3b9cTF/ExfAy0VSZxpnsqv+3aGwr92J
VsXe1GvJv9eGa/dxiVbN4qmUeMrGWNi013NpvVQYIfQZ4YH1WxetmtwbWFtMaqBH7hjE7KOR2QsJ
WDpgCCCtucPEAIs0rHvjsGEgSKcWNYygF4F4vYkh/gSHl9ur4PgcZRPBYSw9t0TI3CXn7u468crL
+eXcw+S9XWi+9qIVkBhDuVVHBziGaNUzPrND9Oc4gVKzg2MZX/yLgfg7AIXgKXrbyi2swC9bgAIj
Lo4OgHDrib/6h6wRMrJC5QJo+8/3cNv/aIKd3YHOlf8eZzvYundx0b8cltbod3mZClU1R2Ufrv0b
MdXOjTuD3o1Kjab+tj4DTbsWj2P/SooHpsrEXhWrveyc1xpsmGLTSZsNvtQ0y23YDgSTlmoC7gp4
AgZCyy7GW+7bqO0LYRsSSDFMShmWOmYh1lE0VDU2EYF6eMuMdqRQ2NEHCd6Y4mjURMP7aCJiH+7c
/CmO+ZjDpjNnDZ2P+DszMhHZ8VuwUq1w2WSum//gO4LcciEMRZfWgBWpA00P4z2FZTKil8UvrE29
mRw6lYaEvVwgaHQMrkBQqi1u0V8YQ5ra9Oc0xQEONiWWThCjJNHnqJ2iJlJmnZM0ofHwiShT2N7Y
Wscg3ybnDRrawfxDciKZsnBEEweuSMfcvqz7oxT2Mt/doUhWcAxh+YWpATLKqLfV2OAEcR+Ma1sC
tZo1L5CTmuoSP013ydXb8EM4DNPqlbDDWqAd7naI4oKNDI/UsKQJTlytCHPClG5/sXbxl5+ub8sL
QulAd9ziWuhDLxfBDSL36Cs7cdQiC6nJsD0xZSAP/0C8+bYMUSpiaWWvt7CgdCk1Bkv+F/wYpIY1
3SEq2B9jBmfgqU5JzFEHti58gASX0/FH3bJDu9QUtwbIixKI4Qnuubq1ts62ugueoTNCMh9z2fzB
WxmurcDAXV9leRYbafBs5DU8tn6Nb4u9P5D7YL50et7mcXf/9f4/MGFqiwDOhJG/bV+cGtxgVTl7
EznQXwJhnkbOKmuvTCM3BrXPXigeSvbpM2sq4sXVbVuJP+XbzZBkJ31Hh0s0UGpIx0kcEYXxX/lU
1AptT0BCDQH/T5ajnqmkAN4QQuLoTjHzDS4NYq/6pzXTvqCwFMwGn0SdNTD3WP6eTCo62UgtCS2Z
GumsR/TjcujP7CB+5Cj/G2hc2s4oLwSHjjl+lPjiam8M/VEBO/DVVyN/cr8GGQykg7nOKiWyohX8
8mhZtszEU5riupHAgCZLiKmo3bpfWN//8g8PA6QuSYOk5cJzW+3CWov6Su07zX/EbN4QQBxBruX7
llbBUzYPl5FDshpBAsUV4Fa5iqmfd8skDg+sagQSvWZuESKUIYmqxkgikXJKvyw7wJWdggxyuo7N
z21hEroD6Cq1OA1lh9qHxExErh3qut5ONTJKF93Nrpu7s6mmP0qe21/sFc1GgTcfk15ByFh3ucqe
62NCuQ+vJknJp9qUk127IbTiXO3i7JqC8AiPEJslkQETO3qqRuKa3ORtKwz/iO2tYsT7itJhM1D3
rq8Jg5/qSFMRljs7puE4hLtUf++BPE2crjvV6flezVC115/RJ6GUkYrfq775iVGioTXv0Ri+QIl4
SoLEfSxoX84smTw7jzhdUOHCeq9Z8ekVKZeUFudirAh7eeJC7DWQ0ethDuMCYiqT34LJRHaIwx4P
hNcTJ2drtA4y4QKhH7huXBEjAekHfLJ1SYzCx/4PAm0mnVJ8rDHjY0s2xxu49/JWbTS/wAPtR4vj
tjme7wXkZyJ0o8aG74s/btHlSOcCV6cNyaizzF0bmpeDu9BlhTPnJ/xUWZMP2RXdAK50XCWIHgiP
WvxVokSlq2jjepHRShK+DprI4lsg0e/g3F76w6G9l2KXPiOnYTwTCI1z21WSxupYeQ9+W4kVLjhR
I3mKdMMW1v5eiR68szb5oZoocOOulZKrMpsOWhKG0mnuaplJtMfv2wkk7EYpNz/GAG4uHP3DeWk4
hxg5JExoEkVlHBTfTKrJsty1N46lsI5kGXzXu/jkUjfz5eV5v3dNSGitP/rP2eyEEZNFb+85mUyR
BwZ0+AKN5QlnYoY6Ch49wNyRFKCKV4Ytn4+ht4l5GC5ib3ZR4UMJuc0djgkNXfLBLcTma8bXleqO
t1l8zEOtXOWkSBI23QH3jXQ2RPkH/udggUFvTUHes1G1Z1+TkhTU7aM8b0xKOw1vYMfzVPBlnQJH
Of6jnzdahVvA95pnbn4nMZaDqxcjyseu/sBA0uV+xvNBfoNRxtDa7nBJutWiWFlndczpI8sLWRhV
fqpFRbWtDVlWsj/GW6jwaS96ZjWKMB0k8zlcxgA0l6Xii9g/BpzVAZn8QiSjIm0vPwkqJ+NB9FMj
HIymynRtUKFV42foEKG/BQ+0xN50tj4KfmuJGrHpvP4/NiiCHLcxdZsG1HESbgYu6BKPG8hdHfvf
JmdAhpXhpegtTbVC1YAY9lRL337HZbE2cqZivqpdIxK88yHqz4esTtUxvnoWaopJuazZQeLeGLI7
Uc36yxWr1qd/Pwg27ZS/s9Ei8ElMcqhBaQfODJZA32qVl4Pe934cSLBmVCK+haDErxSifoWApBTJ
cEVYnq/3Ei7a+LSys5AVL+a6+muJi0tYljrRauVBcYeol81ftzLhBJuX7BJXEDipcUks1Gp9h8pF
vtagxDwd+70tCVdureRsSfYQHjK3IoarymX5/ovxkA2AcYQt+3gKajxWM3gGXKe71HKXfR+CVQLF
aZRlOPyiqYjNTXyW5v9DW8t/tEOuA+gKoLOpb1xc91s0u1D44pMphA3FpQPTSsNW3+bh8KZfUe+4
86uuU4fE+YXTyf6FNKY+kE6SxzK4Bu2fH5CAYjD2kwH48kbvvWap1VaO0ZXtijWnX1XbxYflKoEm
KvLdCsucEcQEtVU+BNtaO9AeQgUHQxcBe8uen2EzlArGKaDbo5khVFnmu7AFkxDw6BzeLs1h6sHb
75RyPnbzPPPNAyC0BTiMw+3793BL1ek3Ei68TcRsNT46NDogMmN0A9Ri70wIB6fLTk3CwXhKbgYz
ckMr2oJ29RQGIQDW1uz+7l0ayICKEUf4cQcikHXvKzvj53AyQURLBdAkWxCEH3e9mMChgON+em3a
yzRLaLlshHvwn+R+yLVFw2JtdIBuS9HdeibwRL79S6n4s1Qlqiw9wkQ0ezCsiLxrmCjElrUe4D3Y
/dBIFwNlTwE0oyP5bcRegvZ0emhShNzbpoCld+kg9WyKO0v5/SJrKMaYiAeuYzX+gfvCraBHcQBi
xkEKdzayR1rZKn7ov2BkSZMLlRahx/BkMIP3FJLmZ7VAhG6gf51tKLUIZSGyrKZU7DwLfXBo7WcO
7CudT/YD84XQzAFoWKMc9MaM/F6NrTOXINjY7zeyVxhPovrHEzfN25RCKgQ+q3t3jEaGeZ3eNZz+
NBfe2MdJPGHHikNirS8PqRrj5qqCa6VgJVB/eAf+JzYcXnuoei6ClNxs1D6I5HYe+KP9YYDAx619
3jjWhkgZ66NC4fntjzw+tgPp5dUGIXLobnnuI6IuRGGU8QPe37B3/lI01PQA4Zb71bKGxo6cgZTT
m8bWWgMNpGcWwASZHlQXIXoL4OJwHVITyu0bgJ7lWCH/urjYsVspNpTCz/ykag4qoZp2ErvObzTf
fR3cOKd7VabJMqhAwmidotf+pMY7SEH5o/Pt42rnJuUr6AItySU+Xrg2V5orfMom91ApeKzjL56n
N8xpkOX1JQEDMe40hHCMAF11a/id8rvmSs3QaJp+tSFiZOvONeyfJ7QNNXrI+QYQ1Leq7QjKe+MD
ObD+QvZm7HVIxjfTLkPjbrNBwn0tP0l+35IJ6i6iIXaW0/ARBlSWWhhT4gkAE5Y59qn/NI3WzdKG
F/2T65NQDcKLfmzeHnE80lcxAchfViMFWwr7GMQyJOWGgGdFbjY4zZUVrnx1DPAG7d/LlHieOiHo
gggodw+0xj6ukntElcGnJiH1qa7hrAFcPqoyOtwkygvMMfNCwTj7IzCby1sFIlYmNZdkTiuoBKsH
5KY5N6fhgvC9heoJCq6Pi5h1MTU3QaMiCWKG8751NEbTH+FfDsdnDFzSjnCu+krI0/LJg329Q1Jn
WYdpxFjxPpP6gXKyuT6S8TiKevCokOWb4FH/7PaMthgoJZkwXmSGN8UjitlU00XbDhGEe+oaTZIy
jwXNVAftCbcdpfGSWjfiAel2/A3kXlJUaVeKixqvXemHCGhAXqBkjJdVw1X2hIwEmFTPV1npd4pz
3yhE4/N4o1wp6M65d0Xee72BP9N/SgBT3sBFAKHoCV6nBbc/a68oXhRQCeQJlsp5kFbHtzOmrSd3
XNHZqVE/beBGgSu3QNq9TFqyggwhdReH5XqIKxT8i4P6MFzIEoeZ3jtJ1aGuOxt7ee974i4YyiKp
8iI5a4RbehYcGxJBrUBtRkHzAybJlS1q3Ab6T2gE7lNiCNgDcVLAcUGXDv1V8oIaFwr2vFDXIefx
Dco/iNy4fwaUirL/IbMjOFkoufmT59NAFvBQsOqrziPPY93G+HnJVdNbyGIYuWzPzYiAbhRpRrCG
Z9YlyVckL4v5x/KtPx+W3lXPZ3Cy3vU19r+1CBNnw95lLKnuCUSXP7IU3Xz7M53fWbwtXgKqmeYU
owPvJXUYvI/K+dZVQEVnrtErapBP20X9/DSEBiHi68JSjZYnQrpnnQ2LheaYFcyN3q3f5oNCD67Y
1jLEFgusqthi3euFmo1E+D+wSqP3WP+/SVYPPL/k+/IDLMft3bivK8ItHPe7Ja1MZHrkkryLo70a
jd5LRynYrYai5nSukXsioEYQ27aN5yrk/3vbjK4E4+xgO4vv6KnpoA2M7xtTz3gzSX/eyw1WwWys
q92cCdQI/j2ymVasqk27opf4+5Pnb67EDyOpehPcnFIQXSijzByJh3ToMwBsNT0dvVrUBsymx3it
1vWyyCicGZx7kGn/2MpwcT89oLk6fKXp4bi5NewloJxBFWnsEryrOt9RVTgC0dJJgXZPCMrZqcuO
JUpnlDd93BXYGrnd3bR6EiW9nzKcmZBJdN76rd3hqRBtWNLWMEHQRaCi5O0/MEop4JOhSOPpR04o
z+Mn1/hCQl+UCWcvTRO5JjcWIZ+umr38Jy+BHD+bm/P9iemUQBepsGQHdiaQv21SLFjlf4GO+l8r
iIpOdFQt4LZLymEQAUl7v0IZjvrDgY+iLod6J+jhXxsV4yDKySIZDIVwHxCYg0XIIZ+J1ciQnVD5
RIJCWiEbi9gmJjo9mdwymVmtzJNNXa3Ddt61CQQj8s9W7yIyAs8dTOGP5XK6j4bkFozHHv5vQZOm
oM/JSz/aOcsdzmiBoK2yZ7kft/hA6RMeh6LFHbwvHAdzYG1+aoozksdXumuZdzWHZHtfK4vZqi9H
v04E2P9RbKLRlzj9m0utG8BkV3TxxHKTuXE5PsRFD954sR06goHnOXDbtscMCT3ygIrtK5wXKSof
faqs0BlNwkFqbefH4sWS7llGzdwUBlFhi92Pyd4YzHJcHIWPBDcg3836N/pHiWehDJiSavwpbkST
U/gsdH5rFnU4UgesbncdPf5d6NMG9d9VyMMHH8LylSo0ksYecytT3pTeF1aL4Iby18bho/DE9ibq
q6+LgYt0wfO57C9BXD4W19/lH/tI0XMmh2U4ZI5KCRqjbyhaSY0fCZtJgFKtkEvtjn5ut7zch3TE
Ti77B9JV/y87fIxG6/ov889KzhKkEzWpIPWixKqjjxeSKT23vOf0GjGstkjZVFck9bvsr1zfdEJ3
GgnWTQB/Q74xhMxkn/aFjzwweIMVENyKY7/RnJkD5Qi/pHa9xIsFg9wfJwwTur2qnhE1W6nYqYS8
5PQ/4U2WXz22lPEdVUmuRodvN0bD1KMSM4/036AaLhjM/d+sHjgGKyYMtSrOyqHRjCVkZ4yMEGL+
cTgPaRrJVS2nH067NDcWnIXAPZJ+7zsHDz672VLyzzR+vPtzkJJAVGWZg/vjhedgQfd8q1Lj5IBQ
x4fTrdYMeNTzubWBn9587NjgCbb/d63nJ1sf1R9VJBBPkepgaUUJkAtq/0Lkz4lHWk3mw5gai0pS
IgyXvCCpA6ax1gmjBcZl/OOs3+PHVPHJ1nA4bT0hwLZ0Ec2swfch9QcRi+wBTw6ZJMBtxRzFzhxt
tpdicHJaNRAR97U+apvmxIjvLfOoqd0d5ivzBeZKCWISX5IX4GFQXk/OaWl+UPUN4V/BZOX+Fon6
wp/smtWf84LGeYTnCHeZpNXbBPChWKDwAk2Re5DB3yaEoSBkkb6BVOo/fs6yuqWK/M7b1U8v3Rwo
WBSPoNZ2/YyvN8Jwe047Cgh/Dryz2yBoJ071EKcZwsyi0ZqnJ7PTa38nbjK8F4lN4hpnrayR9jpm
RXP6XBlufw0PSdsxtMTNJeHFmeiooY/eNpi7pUud2FStGLRKnRwCXmwTHOkH5lsHeK9rbm8WN7D1
2Q+Ejk+XtU8eCiyDKxY3uIg8d4nzbXaypF5S/Lwb1fnqL3K7QmzpGZuwN0704yD++FhuGSsqg5kf
Qx8q4nQrrr8lhhfyBnQD7OXHZPjFEprPVq6eY8AUbbRWDSodazkYVQ/4oiYPr6cUqSxPKexta/GG
3QgcVWTFxtTpyNQgwwkmwhryb09LBZ9zDOtQ4TT7PdxL7yE3Dd/EYWBj2QZYdak1ATMXJZ9fS+sQ
JibsKvxBqaMYZNbfm7ZHjOujNtbaFFUjG/jdiS4IYz/pngdsuSyRumtoZOxyuZNoK9lEVrY/tR5X
dHzRWew3ugEhY3yNtYsXVGDSdXyf7CrqHrGMYrYiFRT5Zm/P0BDzsac80KupQstXtmt+pOUq1COK
epZvU/s8GwMJX+uhIbIuI+K/pK2QR6T3wB1A+Zaazuc/v356IRkynVER6M+QhPTDJ+aScJx1oXHr
7ygwifXFFimGhRHfe9C1Karhb59MRt45es9t6ArdeTnU4I4PaJWbmz71apK+jS3ayGfJBvF+gJwr
bo0dRlEvV4+BaXDIOv9lkytrUJ9LJdI4khX8TNkE9EuO7HWrGDcMKIB32DLvThEuaOv8ZM7XMXVv
+EqKwewkRL34Ed50/8QNIkVDljQGlW4+Fj6JpNQFe6V53/QrVmmvTebDmNEBgm4iRKrNtC8vuwQd
MqcGXjd0Pa02A/uVtzOeb+ClKgK5CEHBo+iBng4iijdEfqupt07wWQeznclbFhQcvrZdZVbLOiKT
ThLa3RKmhj/o8PUjkEgSm8O3h2H+i4GE0gau8VLg4XEoIb1n78zNJ+CWEQUPcBKRMntwTHQEHp2O
4xjzXDIx+pup1TqzzzLefcAd3YqB3lZgVvOCyf5Bx5n8g2N8xDC+KqylV7dgP9Uii7xUHIedVsrb
uDjVlmXq9f+TADFSSwR68L4VSQN/Ma8OomAFxhowmKVF4f3Cz/Sn3/yepgLrgKyMYPtebOarprZZ
0Vnrx6UQsrIP2Reg3mMe+uEoLVwJkGUKQ//m4idQzl1itzc3WCqjO1jLszOd6td3ZCXQHMUsu0QE
wbh+CNv0L1y2vl8MPzslPQNz57YixEI8hfeybunJZWvuF15+7J8DOenivOMXMCPWMARX/JAweHBh
CrG4LFPHxhP8t0X4yU8fZSesiCmHnk8UHDynYy+mkVLoVNifXqeQ/sOf7rWXNHwV7IrSIMN6mVzg
PmAJo0p9JV4PzTrVSREQ/+ZMJFH+AbxCVmr3xYYe4U9OpNviUKiUKxdqaXQE/rp2AcY2kJfv8b8E
a3AwN/ybJkKvx+9ZS7pPX26r5bOSG7u+yY1RP2ARQJIlKElegM5vRwJgaYDefyMCjSsvrF/rhvPQ
dVBuYzcYH8t5YHGGdbI2aDaCrFu/SbxqkLpfZnulydarE1EQUmiW601FpD+dAXJERD3c6Jnc/cSB
l0hpBbR7s7LaMnIYx69aaKxwmmC4VEhVnswRqvPV8w7oR+qNz161mtohj0tkYdod/QoQL0sjzfZt
JOcLlA+cev2+zPR9qt3CIu0DENjDAfOOAI+IKjr6GzgzHwFZ0zXjJyrLsJ9uI9Dz5t29thXZoADM
9Qw8+TxWLFmZf+3YRSa9P3dg5zZyPcUOIFREiq0NIMR7o6nKo96AV07sFms8kLhXL5IsZMq+z7k4
peHl1mWV1NNdbI70aBX3RNE7vPucXkMTUqFKQ86dEOPDATG/v64I1kczs1C6uig+w4f0eDZRxijj
C6dXQV4WoKMJzNIgG0izZ/gxcho96eetS1ZrSQGpUHtcjOuYHmj1RqZzR/OiOfPsttbZoupjIyVb
aTcPHAHh3wiHnxmHwOGoFy+tPka0HvKiKrglEBIYC1vA7znxruNJr96GwYLSxy1mPL/9pgNEIvAy
bHzxebg05FOjI9JJOUYKj6Xv0Pcqtrq5/8FZa9znZUWfgPCPue5qScZktngTigz4FtU6vgjaHpQk
qKaPGhHNfdGjA6dU0kSlDCO1/HrqPfn4RPro4l2H8JoLaNTwDXD69sgpx++OvkM7+l9VouSSVnhD
/maYlb1s+W3n8DUquTc6PiYkqW3sn5PeBbUdpECM4UvRuHjkf5ViyTMMALwliAA3m20mKZqN2P/x
2y37zw1eJvdPh4W1PHpEs5Cimfoh7x18OIogbv/t9LHIohCrOlRT0AX3h4584bPwt/9e8m3A10sQ
6Jbdu+ZXk3yrtRfqJWGiIpj/5CfMEpWnNM2DGvZBkuk1xjjZ9yyfmmUzLITkHacSakXaie4ULTDT
Out10kzJ4mu7hz4mb2BBlv3l5nT26KeGrvqfMlG37yJnjvgevPn2ndYzOJqg6lbk4saz7/8guIyW
gCHV/FlF1GqTjXAzECpqivYHFw3w7ZjAPNcVeLKkUl6vYzRY4qutMAnQTS+TvPAvLa8lys58VLSf
5JrfooFpMrhSFrxABYPkjOeS+ijpC3fzvWByrTJTVtbOenl6BfC8/Jagn3cNG8PFQPHELjsa0CeA
UtAThE9ul3dT9J0ykNidmFniSjBhHC9WEKKGTj5s1lEokJlP82xm7aADIVVD6b+VG+80CBmVdWbC
fResTuPLR80fbMhIZbZxzHE2OBJ/HQwantuoDZLY1vcT0lNs3quGsXqGaiE2ovKDrpmhrM2lxV2/
9qSuEQQd1CFjtVyZI5v7UM9u+xDSt1r0TcMuBHPHEVlYdgVUK/D7YO3RRs8fzjh8DFc5mkNV+QlZ
wCrGe19VlYBqXYVFQdgG6vtn3TcSKYLgcaKbo2OCOBPv7gTmqP5rMByx4S32YzzBC/9tHkl2JgKg
GVwtmavt4z//Z4/V4hWUJbPNzrTsPu4EiGa9CSanWM0ak6fD5WsGZJraq5G/gxA/dy9C05i0viFD
I628L/fn0WmYJnesR9fAmp57fqvk1Oes3+cFXUn6NchSBpUyVUY/KrFIVNUdnLtsgvpHUmkzui6O
tkXP2NBsrM6g6d3FEm+JfWPgXfgZFX5uTbhbljCALJsMqTmVi0jKwhWWJoPrI/afhVP1VKMnwau8
VKIht9h3u8n+oc4xNIeUXV4jo2Tjud0Q8l7Aj2KEXx+CyQSHFGjhVJD/014eOOCGdUMDZsTj66ju
DhZ0ZXrYp5wPHWaU1jcOn3holv/BHvnmptJ0DpJ8XakDCA7HRSkxHA/GEXh7QBlF80xjd4Y+S+wa
bBJ1tS5qfedEkHpWYI/2zAZxZiulWFo2J+ug+UHCtHmYwjeR+dEyYQP0iDpzFHrIRWggqnMXCrtc
HKG7S3vqM2ePHC1+PXgU6lb5y/Q6nOPcT3HQ2FH7z940p91AxFMF91l50iWue2cMF0ocUfGoX4zW
nWIqOUoEPQ4sPemOntNpwdvz/+1lDIQ23tYnsDzHjjfHOQkmR4PQodj81LGA569kJh32+o2dLWXO
VtlLbPvQvDPajlwZNQ4pXAnQc7po6SHPQ2iD7YLhfvtKDXotXWmMTb6RH0IF4bRYxkOY2EOK/EiG
8XR6vlE3arvyPqQN+mUQ88iJmuQUagA7NXUQIzEog7z8IL+qI9qZPNa8Lkqk5DlJDozh08pPjfRA
7wENzHvRbcjVZKhYvQaSuBqALOhMMwHpkOVcVepg1ziQyva9xm4i2ksrwGRc34otfCRjvrohLwMZ
lQST2bZVwDagMEZbtwTF82IDFyU5kzuRV8yiKvTCys4ufPgw7ePkUjO36KND8eDZ8qzMrGytRvxK
YSxfmCcq27rLKP8/jYVUDpFxtFbH9XkiZPUqdy4uZiktYrl/cT+88AYblMkrv+BQEWkt7wiuBHKp
c6xR1sVfEz68lMWUYPz7EMnXaHt+40tD0fSBjdewl+IespZfSFPqkvdMcQ/WXt+4683KtzSVqcmW
JhkeSGGOHrjfKkBubSFbOa6woiMuLmndmWd3gFvILparsTtcKEKaR7qeIjPRCQSpNWXTS/mpUFYH
Z1tlnRE8i6q0AAlRfjS7SieGgZ++HINDERyNXVwdMy8LMjxcAuoDApll6yHKY63uIa5nOR52RH0I
TS+b/xwRCd8AsXB+X3hOUn+XBx6ys/PTIzr8pGhyBzp/c8DuxQC/qLoNZb0yRNzj1gWYEYakrHsx
mvlilgGGZfnpUo4seKPXqdox8/PFRu4n+pv/5lojNn53QrcJcrPO06RCH2nhbl9BL36zAEMM243t
a4k718gj/jrVhzLkye/qyDgi285vRzXQ2fBOnEZ+pYQnd5xm0XKXOlMI+kDvt+fIansIHP7E3M6k
BgsgdDLUF+jd/pcS4TShxWfWCydz0cz9HyE8olNBc833iHPWeDGKZMLKh8VukvpG3on5mCV48Jks
q0JBSl/fnM1ITIlaF0isIq216cQC3WGPO8bOAvDCL/1abD8jO+MVpl9jNBwkbLELAxRnKUhiRg16
ansIOIM+BbBdWjWkzuMZJNjISDibS8v/UJRtBsTdHB4GrcNVbJ+j5oMHSOkuGQhrgaUICjHL9rpv
xrqWpU7X10ItiN+ORjFiXZy9smYESF6lY1ojnFfP51fbF2OJv+MHKm3lBxAsIwx4ftgGAzYil961
wy3hOBsCTY3Rj8sgGde8m9d6cjwtNBM0e/CPVfDHEpEpl6c3DN4mhAGSacEaQNIPE38BQ48tkdx5
OFIf5H4J5PwtCHI+zi9PhP+M71sTf8Ck793ReXtCCP2JHsbNGQvfzCiez0tqv/B9hoNgzLkxmynb
Aps8EVP+Tq1lnXotAh0q5lGzXAerAffYYmH0TLTyNNNFz9TKVehMLt8+uCTlifRoMHLXmI0GeUpz
VG07QDEOH5ehmL+0FfISfN1Zxs5e2C0ZPr0pPf0AGaGNa17wifi8ADoj7PcWOgDPGSORoK61xZsy
9zSd0nW5Btjxbs/HBZtfunl05mvPenVdj7wP02sdDS7zMhQp0IOa7IdoIIwKnLWDy7ocdSHVk81A
4SqbJYzQiWY37PD1OFRsoDUs6LqEzF5WvEn1Y3KUueLsgbg0+3928aMVi54c5T1VHJ5NlTrueOX8
OG1yQqGd1S3JrjA8OP9Nvoe6qdqkrUaJWl1wUKYF4DcGRTePPWSzk8VmdxjYb82aerFM2buQRDQD
lqZU5N/uJaOKtt+cXLGlPmfvAJDtZPPQlt7QoCc3b2e9qSuuLJ0gjafzHV0zWsl98HzPMKYtqBm2
qrxvL1Jparf9PloMrHy1WG362mpcDQXdhZFs7Ir3jzbfDE1Q45B4PCkezqa12uB7rqcgx1c1uGcn
l2dnsovRipWPwIp5Qy5qkbN7nTfGoZjJfBg/632jmaNxEQauK6Wsrung/COyibsX81RHio0y2qgG
Zg2sx+umowS+Ct2eubRcEICGSFtkwEpzcQpVAKCDsz9B9VhPDj4HGa92YE/LeJdo4yP42MQaTrr9
04dBS4VTMdB5/J/L5UwK2J5B4rsNupHIu8aua17xTxLW8Byor/TjaNnxLGfEP95wUDEAQ4pb8FIX
auArLy8nRS+zukH36ogKcinOK6Nay1ZcVCumQoeDfyQZOE/mVIDDj8JejgfktzrGBdYX6qx/uy3X
M+bKsbu35gC4DxbXD8jKyFxwxvdN0A6BBDssTx7+16FnClDwcWEDM5w79A08vp8kBRLe+miD1m01
LsFWFS5co/9V/ChRE5nnQ4SovVVH0HYWkynqWEG1ylYpslrh8zw6EYXyraRFTIf+UPIcLOjUW/5Z
ME/BF/dL0v/R2XbonYnG0MxQlz8HpmdU4v7V47qvRC0jr+8RjN9HzTIOmEbcwdq9j5GfW3/D8Ucy
G6JkdfJAnZWsIkNb7kEEpaB10rmUIvzLmu37g3TOeE5xOh3J5uWaA/NyFROc6DdBitXpn/c2072n
JXt3hdu9RISiYpLxIhCdasXIu/peUzzYJBtC3GQD/SDerX6dwJSJB2ByiURtFx12N4XeUeZjpOeT
caoK3ArMs/+sHWhLtEANIHsH7rc4gMWWbSK6FTex1IIjaFiY7f/263N/Xy3p+VsQSBpgyhX9+Jy6
nnJUAbhWDlRryWG8UhsN2IB2xpGw0Z2Kk8nRDcfxeZUAE1YhWVw7poDe813fHt3d6jOq4E84WeOZ
iZ4f/D6rFDInPJwcFpteXKIZNSycMJ7bFk+wMTcriHpZN8NHJp52yY2UQakaf/grHXMPU1LeF/c9
OtR09WpKg8wUlIfTyCWqCvdJGmM17OAxpfdUmzbkBzzqyLhjOFEFPcWJ12tneGTcO0y1xvg0PrlY
T2QlYNvb6kJ/6Lp29M466gXMRsuveW6vPM0a34PkqOV6BF/IqJ+cjOwR2Ll5jmYXcXvGVi9AkYWj
wd5yAI3TDVtr7JDZmVsqNPNq8LfkE9WYuPO9+cQ/r5wD3QM289cPCsxxiOa+kvpnoibhIamPUhYr
yE9tdxRc8V+ohVRF1EA4aV2I4Sm1ymJKrOffSlu+0fj5BPrW+84iGmNEwuCdCOO865wqt7351vwh
cBr1EOgwXug5klRzGOb9x1vPqxm4UjIhGCBSxde5SIwjBHbM1CS7V0bgxLYZmPthG/73MCcbJePl
34bGXO1ueHT1w9sIDNxpArxE0dwBNhgPs/kPtIWBMjhdDHOHOmgdQSnDYTq27bmfZVmRb1TQQsd1
D68TQmjQ3vQVhxR7Lya6f1L33zWE0hL2U4YTxU1TZesUc3v7RJ9y4BBSCtdgA74tZsb7ZdEHJnIV
+QWnICSvJTfCFgJCg+neOx0ZZRtbKiTERgYRDWAfZ+v7yCvgEybivZKsDxKjlH3pSPdCxf+K6YeK
b/rIpo9DPBCOW2A6zyT6qaKB692w/t/YdPqyAkWS0NJE/EOoNjlqgx6IOU+bo8ZVQlAGnl07o5r5
EztMg6qbvsNOPa/EJ/WuNSx9ho+w8tJBN9j/rhCvz0hFmLQ9PCKe6cEg9HuWNSNwJ1cQP72DZaI9
5ihAIRS/YroG/YSvNA18yOb5aLt20XIObcM4GL0xI2EME5HrHUBDt7aZevy7UG6xaIbRkOW/u/Ws
7ISw4owvkRK7aUznuT5NybQgCeGFh5zGZVcKt68zyijD1/6MVW/HJ7ZHxVcZtePA7ePINwN33K5R
6d0x7plJT4lAmjrgGTphLMsii+iSyU95YVnIU7HcKCq1rKWmdDfya7tBuk4d1SwfA4aCu95Ov9d/
Vpj0pcxtU+GofbwmmKC1fBODzGi/SCKom0L36wlee9cwOLMv1BMNVa8B5Ja4YCIUUeBMDgjprqEc
E15z1ayZ8QX3noPIiThOJoi/KeAVdXw1laQXL0mPPM0AOjb7zuYZVEa5P6ggG88IjbWx9sVmHMn0
hzdBm/pQW9n+anaH8XzEtvQaYTmLv+91MhjUPmlyMz5IdLJ0oJH9Cew0Xl/fdVlQKrSrmuflzeO7
5NWMq5XPS5Cwr8SL6ktIkJBthgJ6+quQniGdf4G2x0oKtA9BPiKRwENJKdURsYJTo7LMR3hwmEPH
rFbvdurUKj2GYY7GdkEF1eI6DQA+ffqMBt9rqw70a/YSbK1dKp3nPt7p7X7+OvwZd46JD8WblDIW
VrGJY0Pif11QMOYh32vhZnrcinRKRb5irJYrY9zSCbEYCKGn/YLmSJk0jn8a1RHQeqFDGY9AfqXS
3Yq62y97MqTYfw5ZvOHg4Ae1gLa4gweHCEJr/qI1Or7pC/pteRM5kEevzKRC1sXizngEx/wBfdPX
+xeJKIHfaNWZufcGI2aWjAVqpsITQBtRNQIWTeff6tpwfxN4FrddDxHQMTGRgXmzCtmXTTYaEgA6
rMyjLO5rOukp7lzr1VRy0+CY4MKS4HjfcyHBBWsZHzUo0o9SleMXW15EfAWPD4qtcE8LAyRkh+El
QspWdLnSw+5z7o7b2RJAB/fDcu1vozUzoEBap6CNrVHvTmkalKfT43SclQg6GvC1PrjuYJQxLuCW
HhJwkXWLcYJ741m1z79gJIXnDjm0Em462nAx97dRcSQA0dm/ghQ4laFpwddLup9dF/GPJdRWfg+Z
2oRvZHjCpCbSaI6cnzd+7MIdaloi71qKn2/Mxm23dNVil5bgVQs+0zL7pyJLVs/y+n7UlU2IxPqe
ixiO5D9tLIoaMnOZ9n9jD4iI/w/VUh6URDjswmu5Q3056uLBp5h+HcMhbm7nhgaA9ZePd+zGow6i
MGg25sLOlH8Cidr12Kz7rAxhhPNAyaare/9b1HMDEskABFe47cowun6FbrQVrbuVabrMbpXWvgbd
iYTzEz17kLCDt+iUk46pIZzGoXppXG6q7KnjAwXrrq7pFfsvTpNLNxNNCiKXWSOaHwh5bzL7mRYh
HZKC+U7q7dRXR3itqVi4o1HSv6z2rJGjAe+0aRuMCE2uZU15OU5W9V+0OhGoBI9oQoGLyvHM6Jvl
FikNADqNl2sPFo7PI29eQvMtMGEE73X2iVL1wLJCTNlk1AMZkW0zTgFouSXfcZscV3a82E1s7OmO
mBEL1qFBjoQUWxXZNqEkxiGZcjsMmAvSltf7+UvbM+HapPC2yMUjtGaCrlMfxzz0BBQ1JFr/Mskq
RQuCIo2PkuFkOaltl5Qwd4ZDCH/e8o73/Ur684TZCNZG3ksfeUMAOvAybnDAUkjI5mM8OuaXm3ah
blaPz/a8a77AZeVRqO6q7bf2j+fuv694+yDpUc1of/1gvjCJ4nzIX+RVB+iVBOfOJEGpmovTFPiQ
m/CllXHnti6gJHZSHnxbE2AHgHbCZktVc3HXDmRMdN+yWUuSMurqMVJPErGZstHSAOlsFrUo8e0c
m/5Fm++Ev8hb0fL50lms+3MtjnQJJpkHh7v2Q8jPHxpKrX2hu8gYarEGcSIKRwr2ulS1okB4lKwu
Ap+EW5UP/LruSvun4dUeKXb6avKGL2V7gMTNKcDqUYu2gqNWPISWQd/vZ7/L/i+bSJl+8Dj8doVN
0ZiJaHXbDnyDeyk3l36vSOTATQsikocTiLUSqo7fWvHgrK23u7LTB2VJadQ1ACGSEi10FcqvCg/A
iwWCc0ysRrKUMfs0FNedSIHJGXrp8mOV4pLzm5KwmeXlM/xii25EQH+M5hY5LrkAWf1KkNm8sqgb
bfCpR+2dFSFtQ+MwJiBN9rbA/qz7VhFrzinI/XHTyEDjdPJlP8NgqB3QtqRAfZJZmEbmZeykCbj/
7sdSnAmX+JvcY8NU0TT3duIN9FrBtQaG8Na32Dqn71BAs2hvK+cXxjs/NyUvXQM3aesm+J/CB/zy
9l4RdO/1cleJhPY0awFRzoeJrx4If71qVqS3YSbGozawtqPXrtthCIpmNFNVtwlEqUup0AVP5DF2
/8Oa69IAtFE3reRT3Yw8BpGbf7SffhlIJX/ua6q8KeUClIkqBN08t9z/ttSETON7lqVxV3rKcj9a
GgmCP1s8jZE0ja4rDQkGo1CmCFoIrIrT7pYmVAAmWMOnlfKEsBmMwYQwvG6ZMlyzH+MYJ18ykc8j
yWhpNkg/qhMR09uQ5Y5MrNHGE3EykI0hRSWzO1RR4HW2fqM4XxBqVoQtFWPDjQeLC69qHO5xQOOp
G/Sbr5iAGhQ8Rhhx9ogtX0JoEJZzDt63p3E7OiTcMPvFR6BKdmbbpTkg2C4gW39p6fncRzMd5nus
A/MjmLnCLPFEdzLa3herDyIuj3cnztYnScFRtEQK57/vCUpySl1z5pGLyhxvJzTcoqKeukwbqOn3
mVbNL8GtG5cQQ8Eu/nSNus/AQuXDN66fjSMQ9S3UKkLIxLFP+w0dhW/jek/0gsyk6u+AAizyDXmD
bh2xSMzyK6URsfU6dXec1VD+IUbqYmKDF4nZvE+QShzdDaDjAlgtbvCO/ngigrVlW0QAkUr5ogW2
aLxEO35FjfNo0asU/zTbRMVuLs0lD1WmbXsrJaY5qusRQ4b0oWJ225exwl8HPHIbecVQpc0xrBTL
cbAqkaQ17x1Fu6rmd8bA0yg4KbbAUNMlY+I9JABpGnnexuBkrCApIwo1HOTBX0kZPPdE+K8fFdnC
4TJXiQoI/SR5yNt9Os+c0rwVMLD3AFM9FO1IYSkGD0oSkpkVp5SRpGLMRZLe0VHPGShJ8xNysH7e
N/keY7bgPyp716b3L21hX4iChveK+nHu/lAePpaa0CzFhbA1V+9qqvlYG0hxsxs/afalTFvRT7gD
Wvfz/OmgI8VFmV6xPwrS+F2Y1c1P3v5YoQHwJ5zbn//0PBjY6rtv9Xwidw6a6zgom8hbgrASC50K
Yzj802GnqqK0AK/ATJ9Y3V0k07qLP69OuQZUmBecSjU8bpRIc/mkB6dWM3YC6ofxxjbJz14VaOLo
dns5NcudXdfsdYq9XqpI/c55UeN8GotDvb1wWZ4yMafUrXFftI/hyqTYrxkhdEWxHG/Wn8v5Z+jU
DblonB2Int9IbvBuHZoqxLEMA7xpj+80BEm1a0d5+GXl32bCpnnmq4Oc8nbmRwhoddr+hy+WQ85D
t8ZS0WceA63sJZe/TEo1mAUfClxGFuFGDBHFczWJdeJs42Vn4YvOSzz4fJNz4tT0dmtlwBjnuRho
Zwp0HYD2kT7m5+/HgHPxpXWOGAcHQllfyvOSN58zhoAapmXVZRIFRKGzcLHXDMYUvglIRM6GLEfe
+SHrjd3OoqFNvjnsDpOQEMLKfYv8orH0vHo8geQQAaeGI0RQkrnpKh6/KW7hLq40+YkAS//dETxO
2H7msY3fa/38eIBjfIMzFUU/T+1U/4LGzmesIKOrF/pxNDAUrRvXOpzN6Y4c//OSHhxUeNeGiPGN
VYm9UC3hbitLXwqUkthJL4rxDWtxAsbghu7RQmFcUSjEMGgpHBut7AQGxR1tMxKFsFjX7N1/Yoow
4Zu9V4rnPAMkSNUV4NlwyOcNVUzJb2iJajD7c/B+IOzZ7Bg0tbhu4Y4VTe+pz5jVeJGHyzg9IfXh
VMI6MFaPjFxcsWvNolioeomylSdfeGwzodtoQQz3wcI9scSYhAmbbVgx5ScwcHInfQFm19Lu8q+b
n+T4juFkBhreVgH0ECt8NRhnkbAlFKnnY1BLSoLtrUwPq2hVfFoYNEEchKl7CJ95X7wJS8jzkYG/
yytgVo3C2dXJO553PR5DGSiyvnskZdjEJjCQfVfpXEJyqv4XvBLLx/aCgNV6dp3GMp6rQd/ZERFd
dZ18vIXBpoqI+l28f/6IyDf2hX0xMvRvTFc3MJIuyCHr1R/vCHapbLATM4TD596dBJ09D2zAyJs7
CAsrlWKp4Z8Hp66ER1ltdYqx5H9P3SYQJWo2TL3sQf0s5oXummYnLzZCS90Gk6rHGnsxDL0xd94W
14TDPhVoPK3zPsoSApEsSfvlXeYF4dROc/X2ZUal41dfE14E1E5QvTzNoleKj4D1wE7tHryxsXVv
sQn68VaFElVBp5n9q91HkvO00a/l36oiksfKk0B07wPIVKg3sIyBRMlsuK28Gn+ILcyieCEdU4Ve
WSRFWjApjIPSLOlDrRiYdTjorSUxKTqjUhKd5zuXCpit/Uloy/lL1JdvolsRMzJyb7Hzb859Hl25
o5qI5TvAwZ8VwJdJX8g5hR5SUpAu+L6eLeINVY66CF0zb7xdHWnQzAz5GmyV0mVwu8nzMxdLUcuF
QazTRnvcU0cf3KC+fq6YD6FGV30KRWEJKFI/eKe2lvXhSYGwyG65lZ4CelgtFs4R1fndIklGrL65
STCt9C/llsEYT7p1Pg5zPlQtqjrUseZLkB2tbclPwRWNmJliq7QAj6uXtGoNsMldXzICUu9f6zFg
mYjFHB0MWO+0UIVGSz8jP5eOseJR5JO0zRC1ad2PwdFKbWkv+59GDRCBCLIreSZK3TWQoVwZKpWG
98hT6Cr3HbwL+lIJUdTDAEx70KuHkjDqqx/J0uNYqcYgtZTT9PcG1MqorzX/J2jA3q9WziFtTeEj
Ie3fdhzJpFV3AUE3Xts1vTvPUcppto5283Xl1zk0Am+zvVOnr04T9z6SXD+8y+oi9Go+7klZJB7t
+h/TYsIk6WnzEhlrFqxvvnTAiYk+uaOa29llF9C5qB57snarxhMZYhg+Jml64wYSLlPJYFF/Ibgl
joean6m8lu5NGZflCu8KGWkmBQNx6nph4nKMuhkcAmBnOYZLo5bIvnhDLq7e8otsnWJD7mhUW2oc
YIvZwPriapMsHdjLgQ/SMpx/Icx6vxvaN8M/23s2PGQpm/AE5vJTam7DS23acNm481KZYJmlP3Z+
fN68VRbfrvenLPYZnHxHjMS647my6xZjMS6XIhwRC/9bW6CRr6dxdM7jkb4lDX9q8AHmhFHTEnWP
SBApUwajttOgDBztIdIIWBbghI7K8pfNWo86Ygl1PB0hAy5FmC3KMNvP/w5dm5qXiilbNoLqewz8
HToWmXChSQNXnplDtRWbnNhTPIadQGa63eeBcgoLuFlAZIstgLSVsK5ZDL55XW9b5XmpW+a5m8cW
UcCaBm3lOn/LN9KhD68pfZVsGT690xKxsJ6AUkrwgZdxw1elP5H+pKLRcM2Q8rzqBgUNVOkKdT3e
SBf1+X9bRQPzia/MqbhPV3vuSUj74wsScZuUIv+jSL44WaY4adwc/+ed1Igh+bc6MoVKIarv9psl
Nj4QkWuR096JG4pNEeULoof01DlnCpEV5mzwIgKVa6z8EAf8O7Gp7l8G4L0wQ65D2JqeFDFxcnfI
Rdm/O39IOVeeZqR1YbJvMs4/xyuB2XYwuqMXwXOtHsWwQ5xIcg8/o/dHzSpMmhG4H/XOoQtRc1Ga
BQsLkBQfE1i7DmvAJjyPcKRJUr1rZYj8FlufLIaHutfne1Gk9KQcfeaUeTPPrMqk26vFHvzJTXqO
4sto2mYDYDwslf+ta9szGxS+x0XiJsCeU21oaeYDInCev3sH6/No9nZ//J+3PtpaIrnCjwkP5Alj
WPsf/X8t8W0KTD6TkFFf6XoM4ve5iZ8Ji2dR4VkM1Z7CpdmcfWf820KJGQQ5NmzEQaq4xT9y23ic
LOoGjSiVbSXBHKx0MuJjtiUfORlUUJ3ZzUniQbktJTdzLgleznj5dgDF9gdDID7kD0392H4wWNbF
+9LXUZjjToqLOvJKajNZmwxutT1Oh7uUVc5RG0brcsB8KBntWPdDdOZKGARM/k8Wx4xXnNIHUFMO
UXCGxAl83Vq/Ta9rkO48AcdR9iyPLd/v1GpprouqFmZ52c3ophGPFGwO8uMusKUaaP2KVCnlVTUI
7MyGMQ4uLDFOx+SdTIcPPRqTjR7Y65vCXnAaKV7Gdlaua+/E4VEJ0FfwppgQOzoWidXSVCQXBoiC
EGh1B7EkLREGWqUVGfN44soGozNgW4Y2UaQbSbs/4i+VRhNm5GIuFspu1DLH/UmGRRg+ayWFaOmA
svKT5dl5NpjGaXm/oOY4OYemjM3KlUoS9r3Md/dFZ0CWH9beUwUR+Jb/HI3GO2O3em8y2ev6ytBZ
feBwKK+4OBQmg8zTvZeejyBLnSrLkjUjvY6xSicZWmIrFiT+RwBKvvd1ULz3B1zJ6L5rhAMNES3s
Vs0ndjAyDCdKgyKW2vqWFg09hT2w5E89GmuHo/uueUxsCPAU4lMa1xqUtK3Ti8UbY7m893mKzes1
QsgsbBrtOvKOTilD20ew/u4rUIV38W8VGSNKrTcykIcPGob/T03oRZ5aIhITdRkpXDZja3LkXmyt
+6EDFezeI2U5VF5GI8pvuYslcxMOzTmNu9z2ETiPDup2R119dGQB/i2g7LjJvcYzMaJzu+OID6TJ
sulWed6Qu5qHM5+6jOYyQwzjZJTmypWzeHKN4ZDz7mg8Wn2U6L63mBBwgXqbDSott7MqyEBxCp9k
rmRQilMlmuaeDOZOUQbUfJgX6u7oPEMq9UgdCnJYt+nosciYE0eQC/vE9wyN//xrpzy+As8xixIk
ol+Z6Z4r4G1ROQNvL2ewTQvvCOxtyKgcU/Rv0kTjbY/nskHCkjmHT/tLDtX2nekQsMj9Uue+6Mhi
3u9LwWP6YMazm2tVmg0riRHDW8tAzEBPMlYCJ7a0Je5uyIHJpiV2qMAFmjWcwyNG9lyc1Um//ahK
cWZJo+7u+GHN7RADtPtB1JlCYg44ea0313qMkd2d96YcxmQBRMULBo1rG6rN4xMYB1Dqhik02uv0
2H2irQEhX6y+WisS26yrrQ6FFsDSzdLH+kmzOKWhZ5o50c5yGlGcBeumug5QJWlJCnn2+uemNu7X
VE/H3h4nzipKu5z3b4fHMPLihjaBUnOcIo0HhdDt6pr06scUvaeR7JNPQTthBoxO25Oqvo8u8Vyr
x7M4MQi+JBvwF0eLK2tCCthqrY32qttwhREMAhstp7nG8w+RT1Dqd7g/kIk6arW2KRVbT+VnirnE
lEN6cv8vkOLF9XKcpWAgp1emCSgA3AbS3vXlCEU2WbuFVpVLZgZzoRbn8Yq0SPe83F4EXHEJTMKw
fyHet4M56oPYCOd7j7XDcE26smD1tyDQypB0Yxd9hwR0lqcVRBHWGq9XDyBT1Rm5kUGfIuWqN9Vz
nF6pwbXeH8bXKP1EpJLwxmNYxvZnm9CYGQTETlbf7OSIClGrtJZGkCH1fdxupRxhZjIbn/T4RI/u
rrX2Xbn1c32TewxhloIbDRZTsu9OFcBOqtkmHz9SkF6jclvl+R6JdcRi26kOodlPj18KfOn3wmzf
ja4HuMYJpwtZK7i8In2Zkcz52IHVbNPNWqDSTm/i0lSdi7LMlElKLRij/COboq5WKsr+6Kotz3x+
F08AK9ihRWUoXY6jFZC7xBYfB0uR9PTMoUt5XWvA5iT2CAG4XQIYBBoBs+yiveYnPyx+2bS2FMHl
2LmrgnkYGpuT+6q8WX4tfFyLnwA6AiB3Lp/Q061r0oXmpAqQEql6bSXJipag44LG6QI2cw17otIY
xtyoWZ75O70eqjcn2wmys5Qj7+X3MvfeUMPebQmComRPvoxVol3UEKu+zC9bm+/fvGZR3uNwxUpg
CjTAJAsscwyN3BGFPFdjdTBtsB06E7TWES7G7D+LPDNyubp89i4oZK8LRwYPl/num78khvovx5Gi
1Ky9rReRWSWQJ0ZqurECGJKvf9ziQMXDCzP+wZLvC+K+nEFkXjVTDrsimMuZAqn1p8d3HMAgymJU
gKkH7cjLOzpiGu5L4EJLc0d4jtDyVh5Ex74+B3cIcW+V/veM/BoyJoLSjP8laxktE7ttoqnFtb6K
h4XXnua983zpqQTdhOuKvNIQcB3lu7aPtFnT7TTBAFO572UzlMCe1YGqENJKQuVY1TZypRXiVNtH
WhkTwdYWQF16kuWm4B5+l1pP3MM4VV5rssUpXzW87Yh08G9xy7xJnYQwg3HIYnC/AXb0OTPETe43
VvlTq3BcN0VbS3PxEE3Ci7h4qcJzTJU6bi9fR9BmQ/r049g08GpWWS8j3K/jjV6809JOzzt8tmio
X4wKBQ31fPZUKkU9m6FtBHn+6ICyQjWYyEc7bpz+0PXxhkggBxoqo3Q9lTqU7DuQgktSShYuO9zG
hm6vxjc1nBk3cQ1Dhvu3LgOmy9ltHR0UOtEZIvLxgirQUnBAzEabHaQl82sRwmSFQKy9t+BUXP8k
Q/myKrb/7pBE+T1TgzkJ2ixymzM78tZd6og6KivM1wGVisqdT64xtnj4D9n4rfJwyp7gd2VPURBF
nJ9iSMDiLkR0SDdJoirZI1jL11ELxv+vyQLYu1QrkWm5fefAGD41N59r1liHS3JbC2/xTAez4tag
mFYweAmF2DjS8ITcD/rOkxI6+Z0/KhckU9m4GwskQqGVdfLsUn0gTeI8ABNDA86tfsQ2FnsqC+tp
b+o5RkxrhqSLZgCXXZe/AvuzU+/1q+njhrbLy0he3UaQ376zz8IbL+dv3L5Z5vNcuxno6uJ7hMwb
LrVuurJbKtpq6QulhadYZVSy8PA3UrJItKlV8P3rOQbpVL0mF5EzXmCHAm1KSzY0CvM3zXNFci/j
Fb/Q7lX+k75qEjraJ3QJjaSO7SkkG3eSM92yA6ssUuUHlaMgdsinjG+GaZ9xmp0G/Ak2KrwhZ75K
N3CUX2HAwLfY8uqiRd8bMrEFhGTZSphlTjNeuPx7kigpjmBszig82J67XkT80CbjJsBxWP0sAqBQ
22pFoDrpQ0Rrpk/2cV2YsnX5yZiBOR3Mvpq1PgQgn3L3UbGSPmrJAcXeubYKOBnAbMqm6eqSPCnF
Sv+AlwWA+YfgEyGLNbGhQgc9/UjByJANLJEbytqlf0DG8scf3iIAjfxKOtWbhC6O5BMuT8+ZyL2Z
P46pWQVRIyjBkEhJqE2+X265TZTCeRq0n5OAM+eZzpeo7sguw8tks9/wxc181SpDN2Eo6YDYJU1U
SJMgRqZQ4pOTzJVg1eI1r03wkYsEeTpeGTClZxo3B+KxFx56PUyWV0wITT3B2eA1uiicXxXwnTA3
bmC+jvCLCwYxAprj9OyVRCMi7rKOvfP6U+FUk4m2eNdk96YdfWancWK3bt1yx9EsDkWfaJo3YBom
AQb94FQ0o2Ro5N5xqHonvSC2cIeVygvizqhAQaUzb36YNfsp0PbyDyq/i8ClCtFmiG0MqSNsy6YQ
jw6r6aBpG5+XDPLHSXMyOGKIFe3LcO551xHdch7PTee5E1glLRwS48ZGGMSlpZLQYDEiFiwHm8lJ
FItMzmOByZwdkuz3Ffl01Hw0COOH7gY6k6Tqg/8UzB8KypMtBi3b6Ej4RJoRF0V95qoudrizeXaC
76vt8REPgwuSKjCJqxKOo1PbV/9IB5yTKt2mpQFba+KLeIZrL+IQsFx4a/VCWha/7U1mSrWhXGnU
Tk80CdmTA8OnergKrp9zB4i0vMerRQPCLFKktpY43N+maO+QvA3g4954ksEPvxW23htNuPnExn8E
Y+SOoZlxIprkxA0buNv9knVbIDqQrV1H1H5Ox58tmpCv3V1szsseW135FUT3OVixBRi4MFc67bH2
PDWGjU+MB4CiKQxAhrC1meRfSQVP4KHlLeaxM+fCY1Ee9JElxcRO9zLIGSuVDiLoXJUQQcizWjf6
Hp8jCYL5ektjAfrxlxZsHCUbMQvNYLY04IEjN5dnEMJ3wLuK8LNlWkdPoGJn+IVEK7s1i8l6VTNV
aR/l4ricYW1tmHK9+9EIVXRQj40vsXka8BK8dt9jVLgG9hxbVlt5wnuph4msPArJ24Ef9G3C/ULD
GVxGuPug8fwyans0ZP73tE6j7c9eL9PhN3a4cLMChZGErRjevlf28lqkLWlMa+pqbGGZ3wuEz0Sz
MSgWvrJx4vbn8e9lI7y7eMybkXIljLqE9PFaT67G6tb8hmN3VigEP9BAPCUu5cml7AeuuTZZvqFN
Dikv828CZUYRegh9RlR4oBuq0e40pxMvNXiPmUvWmWAvQVGOwGjxAJhS1ihEeiixt4lh9r+B39kQ
gKh6mwtJ9HCQwZCepnBiE2DyWNrARJ4Z4bz4b/XjmHlBl7SrYN8chvKmQZkL6fHIWCHORNM0VIWa
LfUQVbD+O2hwB4FDhkMWG2GKEZkW2NxPqboIyYM5QT5kRZsoKvP+lqJKYL0BodImoQerCwuSj/Za
D6Y0yCNuryxLt9M/1ZZhGOPhtGz4sgwxrcuz208u7G5Xce5AzO8+ZUXQZ/NQajVOSsCbSMhbVUkY
vnW47lVgxj5uoVIQVL8mDrDNB8fQ1kVrVmdl1GopK+mjFGMkXGBvfitAYcDysQgx5knHTG0t0y7R
LtENwoMPXaRmIiTeutO9QWqi2w2nmnQuoubkxQEEsnBrQmYikOIMCj/kruwoP6MJqeEwBdDjSHm8
8RmGSpeTL0soSPw5ddx9O0R0UgRxPQ9/clSfDacFbTa4qgDJgTnejw91iZrI7GtnYVzss3d9qzvx
ytOs9Rq4I6R1uUBXGtXOsJqrUSUOc1C0WBh4g3CsLwtXZGcz5mOwMUQmPNcS3TVgXrUfy/3bzdi2
H+H6ah9aTWdMWdN3TFOPhrm7OH3AhMzV6dnyi6cinJItG6KLI8h79ZOMgVLWv/NDGIybyjl8XKCB
Homm+H96nGi6EKQB+Vn7MGhjOF48mtYl0lpE3n09YS7bIdWNHgpXDA7hPXXGxGXxiDVLCSnb8Ztd
SymZdnWnIaBxgo8HqINl93I2LcF5Uye818GEaztrP6V83UsXTJ3cDiZTLhMKgFjfFKmqrmKDIpOz
JCe3ZQrVlJ2jo+UrPiRLB0x3eF14ZsLCcx/WQjTLzkHVYiL0sdYcON9DqdKYeAN4sphZVAEah0GT
oUEdVTaefHSSwaLBGUL26bNofxRFydHz8M7YhLgHgD44wTMc6vCCewxmF0UdPlkFWdypPPNCIJmd
PSfh16tTxi3LVkCTwmYxh/M2N9Hebguscxqj4PmScSO7TJDnE4TPU0AQpp532/9hEqqtofA/baD/
HabEhmCIkNYGiyKDZaqjlGKYZ7T2QTBYKekkCb/pHI6xkqHzeOKye00MsbnQVQVU4u1L+IUNaWU2
XVuBOaquqIpb5Q+6esWjMEEek1yFyDHLrO8vDMslS/1KxDYM/F6OGqIKtzEAp+abo99ODD1clU8p
xjK1wCYbajVBBGIB70g3fUF5RneqjVZgHLIq0gPhkuq9n335YVVhQO5S+UwKJWesAPya8G1ZZf27
7t6d81LzSQ9FRwas/F5RcDodD4178nM7d3qeIVdUTdVav5+e7usklLyBbY6I2uHVr9JvOWENryMK
kLX1H4SqrW+Cooa1gXf1DUEkvvXSQUMVJY1/uHkuIlD1kNk7DYZ1zwGVoo6cokAMc5Rx3JmeYR3e
ilmjDotioboa/ZBbBUzUXoC4s1pABY0hBlNr37JpIDJSboax5q/oXFsiVOawE0ouQ63+/JkZmFtj
vI9xvku0oUR00Vp83+hkqnH1aYC5G8M6qw+05l4nuchae5nkzcn0ugimVPq+HtA297BLdQVmRi+Z
1NxbRBkm1ONmTNiumfGJT46j6BE0r2yJD7jMN8YkdLsFFLPIzQ4F6djCR49KGqAp77zHBPG2XSEc
OdSwz3iF+Rckyykr6vjAQ6zIbXJkrizw5ggilokmM3PVgtvNTk7A3fH1FdYW+tHE6+nO4HkwxOKq
3ODaBQfk66rTzFQYp9TmHzZ02TDpak8ltTlazWaktu2JoDOwuCOkQ6DwOZ3QcbWtQX6GUthLGtYz
n2uCjtgaCjSXPSqniTdD4KLWRFA261haQKBVXJFnnZA42nSnst87jR8KoAkzlLG/lLR/dnm7hlJt
EDF4kpJB7XrL7DteUKxC6QWuGIfPXY8AC5H2ZNPNOPWfi/0hn1lMAVj2wijq0ZtXbvxV0BN6ii0W
w7xztHZ8s4mVfXTMUHdAHH1yU9dnw4lv9NRcHQTuANgbtiwWkfE1QLAZHj3paEzxHfIpSTRXF7Va
6nhuIU4Uj2scAsJ9v4EoJQH2jDDb7VujS1xqcpxq0Y5JWHorBxZCPL1WVRoB3HJPE/GgfgzVPOGs
S9+S21/Mb6taP5ZBNSSkYmajoOabJSv6UeOO+n2Y7kShoD2B4ha9r1SS0yroTdLgKc+8hI8RdzyP
qxYNrCKvUBPAYFmoQJ88ih1v0WrwBhHw1SzmQbNADP1qIibIMdTt5AOOY9kQMaCG+mdVI+zmFOv+
s8OwTU3n5l7slsFppPAAyH+N0Thna2IFijoFxmdo2znEkz/9nwGarKRFp9adB9qX5O+gsTpSLns/
J904CcHY5pSe9GznTxZAjLsn33evlhGZ9z4QT0ruUZWpWInpw5pYI9x7Q255GfdRaMWrwspRkJGx
sR+SVYLcNvlxpAj8sml63Fbgs0Y6tDjHkF9Cl/P06zHmji8hzFGLHflNiQLZqLE1VhL7cLo9h9bG
bwH70+NtTGi42hYrh9AnpzsmT5WpsfnSn8vtxLDqE0UBrHmV+mkZkIzwHLV1+1oJZvta16MXyqqx
ioRTjRkNwOzZvWDe0n+TILoyqUIlYtKaIGJD3rrdJXMVnzeFZ+TBGBHsN1nfZ2ZVbt/AGfklyGOI
UW3AE80lkswtetBU+l9Yyjui4g5eKDrIjlYRHwtNPWdrc6QkG55v8rhcM7pDWHKsXr52IzKzC+Kv
QSO8mV3HW2G4gDspiO58SBJU+dw8Izl1xxxZtbkoBw1sRm/ptRp2RSwL8aYGI8yusdH0d3j05rS4
O1XqsqMKM1BaQ05xk1PzlRgqSYi62Ap2DuDQ9Oj9GDPoPTL1kaQ55rf+pwfpEwi6woLpUrUuWYnC
ei4S4Fg+PMCQpFxPRZe+88xqQXbC6k6woJQ5Odl/f2vC4xSv7s6m9aXnykxlFHTvszqUKtVwHKAr
OiyjlwrAgdfh0BmaBnizT9Q/mlRND2669Vj/ER4mOyb4sH0xuWKty8Pfvsy0ogYqFylCmXAskMvz
+XgN+Bz8//R75lgSLpcyiDw9vrFTC4ZnmzrepXjrCOvmYNewG9EqPOX8y4HX0CyKcFZfkX98XtIe
iT6Y0/zAYbBdcoKLvplEb5nclwhaAT4VKu+giD8GhEBGdL1RS98kboA8o/htKx0GbTvPR7q+aAjL
NXIs+5rUiVduBHJQAupa4XDK2Y5aXqtSmvOBcID90oiAZBwSBAMbe6YgXd2PnvITKkyjbfDAWf9k
MxCAQ7Vq/r+anaKpb+V2xTLJBCoGm6GlNFWO+7ocU8tAE4Tk2gcnawbThjYw7Twjw7POFfx+Dh6/
YH+FmmncG+6up2I9+T2bu4+5KJN96VFvqGz96M8XbPUYyuUKa3JTqbAOEJsRbcDDkpEK1SXsbixs
9tQUOhNOzOxwVVBaXMllv7iFc9MPyfEx3swhxE0TPCupQ0CEg5dZFDG44BNzw38muBDvpNSA9N9m
gGpy6GUG/uHdhwn23wv0bgDs5ZLtQmeaAWz3Ogj9x2FpTB69X/DknFtDg1JEiWkdWZbwPy35mWV7
hLIO47lnOuFVu7BJ0UAqtAeMZBqKIPapBhXtNsrrEqs8MU5ZfwfMRuxZIKEiisT7ShIpFtqBFQga
CZ9YJCpKUaLufLdVczQNGmQKF0hUER40ygSN8hvQ3G+/oYKf9szAX2mG4hosXTmLLM6R6eeCFgCh
I09DxeLPk1hnnnl3NtjYaU6v0m3X/kFfWNBOmwzMQX4YiRegY+whgxEyK2tkrYoyvBVvIdNPb0g6
YIBQoCcTbqQ+cpGZiE3kIWwMjD9oDm8XL9Dl6vNQbRahtEvbfvcQERT8QMCNSFCuQizoxiL6ZevJ
1Xuq1EMAWiD/skypb+xK07B+/8FNIVLfBg3bxSLiXy/09nCoEC+6WvTE0wi2dAkaDvC5V4phK5gg
r5USpYFzsh78VT5mErW14KeeffRy6D1agrQgZtGsSCaEkQiGCS476v/txeh1rtMTA1GF6PaBYCL9
giHyH7YXKp+55FccDWNXQ4VyHVeNqBoOkCuLvW9/QhOzJldEDjjuAWbZ7SyhCU7jipji3+GY54YP
N0cBEGWWrJg0fg3iGg7l3ZkCM5PqO65MKIiVYmQOm/a2E1uNq2XeJMY63n2A9F9lvABndLGwsJ1l
Bbnk/1VdZB41Hk0pGA3MihO4Gbct9ZXopRoVesSBWRVpL9urMGv0dMlWoay2Vb50PMzKZC2XiCYG
HV7JHsjT9uNQxsftqgde0/2XZhbHKfmoXa+jqbiaLeKbo9F31jW/ij73Ef2+rKepuAt2+24X+Qjo
Z45M5aZvjY2IBJwiP8MckIJ4KwtXbZwKye2QH1QGt6qM8dQgYVFzzg92QnsPoXWRl+W3tIHJMeo4
HYHr/9Zzvw7F5otZMtsxTLo+X6A2SOudRh7l5+j5BdGU0+C6EwY7Z8TqJE8S23cbT4IY2JtuzN0j
ba/ZX3K6q/wniMef6UwWdW2dTw0GuedTIO/rrgcOzdcmyvs276AYhcz8AFsLODguv/Y9xc48DN4j
1pYErJwVLdcyzbXR0I7Rj6lvDX0JqNkdpSgwEJHJOWleA8dYaiQl0N94FTsO7+44Lh6BgUmxYcxK
zF228YcP/ezaXwsu8Z/T/fAn3vJCe/I/bBORkJNtbpd8puDZOMTcgImBSiJwBXXWT3BfWhDhvW6l
Ih22qWPo/iFA0AzFTgNGcoYxj5iW11450sGwI+bKb4hNtnmgc2AAFEqxBAnHlAy4s+Y7pbo19cKH
HrpxKIQqdY+QEqXNgNwUWv0XY5yQ9Bao5QphzpSAGpeou0yWXOxrsEqumdo4EU2+f6Q04+tocnWp
eBO4uBqCH7ZOwZn8yksDOKz1tlBJm6Zb+7cEOdCzBmhv1+xIcBtPx6cDvmaJqLYUwSCOsLWuUP2g
n37PrgalP5jIjNNQw4WatUPVp3XKFQJ8WbOpLKMf9s4l6tcFHgPWWDLkx2YlhghhE58cE3volTCa
rdoHTKp+9jlJ0ogZg+X2vTFT9wj9jqAgNAKXrgx8oH7AfdPMHf628Erysv90PxyYM916iEb9tmcw
LqM6i54pAs2w+KwLts3yso5BEpaoPEz7tUARoXpCquIcEniCYSTwfx5EhJGqX9r7AyIbDgP213Hg
rDvwnBpay9ykZ15do8iZRgWZCer/Vv6TC8I/Ky82q0Y9HKxXP+4rBkL+uSDZbJvwAxAKDMl6ZtZj
CuQeHjKyrzNGt8BqOL5XFz/yFk4JwAcARToJ/RkMczI9l3puKwydwtw9bcPQ9yBnVeDbsyIZbZJK
lEHpQXx6U37bV3dUfI3XU+Ul2u0CBBvp+S7C0TkdjME+kPztfgmBzYiYdfWAqYP3/OYIR4a4sMjL
pZWJTOj6DOGJamtZZECGQE5v5zj2X9T3TC+nmBF2/EvF4/jB5k+W3/GQxThPOl/hGq2MByUVKGXF
bSxOsO+g4e2+9STIzqAkWjIT5Ml9d51fyFz9ThpQBjnsara7lQjZ/6cCs5gZ7JPCSBp9+h2QWNl6
+iPsJTuin5n/NFYeMBr21649sYT/AzNRY/+MUfTuUiBmQEiUvhtcTwM6HHhcVi78Si4x5o9Xz/gV
YxbE27O9vPk6jiB9CF5IfZN28JfealAK/bdJdVTamemH3lUUFjTrvwPCFB+GCk18k6eWCCXm9wQm
qb6YpqIQr2H1zSRjYQcZV4wQBhgi1wM+qcIPBeW9TuXpRx5oQwVM0g3bPpPhVzlUWHgYEUXmM+KQ
wQE3q/WYxIk5PfgG/kCg3EP1GntwXIbRhHayjd5VfO/QW9iA6rc/mpWa8C6Hcgon2Mkxe+EXdHfb
MjvS5qJBK3l++zJESmdPIDQM2pH/RD4nfnfU18DmD5NgYGE5DLXtp+7bKity34sFmb9X4wuEXMVA
W5cyRuwrM6Jx8Y15QyJ/2pW+HmjSkk4m3Pu9iOdTVoQl/k/L0VYRkoB/IrQMks9HbwT3Q5Zc+Svk
3LxM/hL22dch65Ro+pdu5mcjVksoZ0GCcN/1P3f+1G0W10XUO4TIIqxbxXwHNbs/MTsJRvxHYB6X
lODuAFyP7zOW5w7FDeKq7k3gXOyILkev0ytqIpdG/ujm9xoJGTyi72I2aOA1Vo5gpVqxf4Fi1Gkb
sJUwtdSTVcI4l5t8qelB0JlbTJQuhb3tHwGiRXrjPYnqMZE1+VweieXNYbNcbHKk8pNoeAXUvCM4
KyU17RLXvSqUfxM605N6s98i/fawrHT6aQKXCF+V/l0rlWM/xDmtUbUdEF9wYEyBN+cF25A9I2Er
U2t2yQFR1gASm3Ya8v9WPSaQU0p9mgH5EpxHRRd3E4rPs4/N16tPTjTpB91ZOZLDDe/8fqy7EkR2
n5w2SQbtqN24bRcDYLUn7sLVrEmkZTkrbaO/jv5txp1YDaiq5cq68EWaQa21uLDCS7/8VCJ6RBF2
hdSCMffL/HkY3WETlD60fiC5mrd9G7pF8O8FArm6ISal3EbK+h/E+HKQhxjge0A3NIeAGI1O9s/R
cygpeemVAYHFfX2KWj1mV+F9RGqP2a6MtAD6ISVois+wXsy74ef+uBOmApXBj/2Qum4YGmC7lQ2E
QM6w+tHXg53Yjqu+YjCra+JGTi19cKcwDmXNDj88HF1O2/BF2eZcqNbKzwbs5gz1G6xD5G1H8jl3
2NS9suOQQydS4dGeAS5X6LMb0frR0F6cP1SipvrvRAaB0e920RRy7f9QUl3qs+jq592DQnDhCErQ
Nfi3/pz01Erjt2R/hzwTng8TeEcAOS58qtTh1zJpQZUTcJuQ1gTzWXEMel0X6rU16egI7wjpXDPz
+t1sgKnkhekQqlPxDW47OdsyEgeImm3E90ZMo3fjaerW423apQoXMKXxb3Ty6oJ1/euICh39GLbY
aleABacFlG7x8KI7DIoNnTbjtcqnr7mDyst/UK+gBTP7tiLhS9OG7cJGmGBCBUi4x7Ly2GWDelt1
gba0SnOVDKz8VG9n2UpWzOTH/UJYTS387+vPtxBeXHzsmoYFqil0bTFapnRJ9CykBGqpaNVm5+JX
2hydHdmqnW1Pe4v2XaEOKg3iEB1Pp8BdUqNkuhvzhEKgPLeVacPqek5z0AqpcT48xP4Hv66XDIBw
JXMEopFk737N5LNwjQda1idEL5oiXO215JtDIXg9umLzhpGJgcV9oqoq3Bi3rlJ1Y9Fpna02nDyV
rtHufacx4hgHlrZydB2ydWmYXxUT1mt1n8XmREVrOxGqCYJ/1ToGP+sP4PYmu21YFQjwjnwhirFv
3AyXgB8GvgnkFAuptgmyaKjBucQ7a94Mh3Kg8KV4I94CBbz+gFh9sAHX7ujLDvUgBzD+YYv27r9U
Y5Cepbt07rGwv8MJFMy2Ak4LdFuMRQReU4Mrd06MBKgxI1O/SCPnWZVBSR26IfQRHDVS4qSN9cuG
q89A1VV7YOK0m//oLCqhe/LYHCFq2OAADkuKFDSl4L+GmVWggnKB1C8byqJh/dmG4wMEvtxrZFC2
xDBFNlww/CcBfFhmb5vi51nmBYtkd1JtPYKSXgs8nVpxpzWiL1zX9wZmBAst1f7hwgDcYrsAsAev
0ytE2JiDJWnarbQDuZWqTYb+buAdjMIWvPpiGEah4FowIMN4CwU7T9qevlA1vpHj2tuhz/GXcV1T
pp8v9Q+TJjfyEJ4hSq9ogmis8dn8NfGVnlL4hbLg2zVN4zCE650LJ7mZEB99mXh2wLUo2141jYkC
a1TJxxzWI9mcERqkqwDLT/OFm3D+qebroXz5kFwhmV7GpIiS1Cx4sYzMowYj2CB2FTNTb9wk+3kl
Xf/OncCq/z4FqWzh/kVy7OS40pSP/XelJRpnHdRPANYy4VP2yO53Mkv9FupB6rSJRjbVp+M8S01W
6lpMRGsaauZyvo8qL60cFbua2evcrUKC+ZXgeSe5eX2GXYjv2+rq7JZnV763GMlSbzrfluuDJjmP
ZR/SitdCdlTaRoY9FjvxWVKgCvphzoLYdvaxZtw22SRpN/ZZnc+ZF0ciKEEl5ULS1mviquBFoPXq
eHAyIQz7qWHDcdiT1EFd6Br+0lgWIJuRqRumkTb4PsUpiOoQjqZkFle1XzGSwEqaPcd2cll51ytq
EOddCR5pnN3U1rzlI23P8a26IDpI63XM8+DVqB9u6YuetLNAuPo1gcN5Dk8XKwlVi+mWgt7JHeaC
L0wcJRzdtIQMOdj5/muTndTUSO9t9BpnA6Gy9ADKDMIBJH7v7LWG96HySC48h1elOmmgPpW/2Uqm
NVtZKLn5Bgl+dJ/ewzqc2a/sQD9WuroDfG+Z8jeVIV8zpqwN/2DnxOyxexknHLCGnF3Q6VdK8xIG
ZyoejHGzj8mbR9S5Nf2hkPmsxeCfZHcHcep7Gx4nLKatVullrN0G8sRGSWm71G5acLvuCGKCrgrT
bCdAH8hLz1bhuTSlwHOmEKXJ93HvHsGuZIY5CamIYWEt7t+B5LoRou+ySYbB2ftxL//4emk9AzQT
Cz9zseRehbIKKDQcG31/Sx/CaH7UgZwKqNDcSsqZlAj5Zih2xMF9hmfpg06SyWKSxmFpBox7NpYu
7VColdIDSD8iZW9/7vz9Ue/j9hE/hMe7rDt4TGXDjntXbpMTvXwfC6iagOzeoqomZpXLGW4eXYYY
XUxrz4ESf+vKAYAB5wIBIi7W+47zmyzgh4JrjDHH5nEVg7sg/kaA5uU+OqQcUItxKBqzIl5U3o90
wvTAqSh0iKhdNaFT/rOToOp2RFEhxTxOowVaau6KU8nHm4XmWYsPz3036US3QYN1IScHCpiz1g0i
3GhZG+3onMC0dKWDYHvYeq3Y2MYvR3HdSjE/AP8UJHNyREKHgokFxTRqioSuOJwQJToaJE4g8azf
hoZGM6V+klhM6xd/aDdgbNgHqq+paIVJEPcsMjEUnsY8VfhUJrnruYnl389IjwuJzURqSYPf1pyz
6c5QAjSvBCmOEStMNMOSYboYHMosFJFOdeErBwaDT60RL/HWkYQrBqxFxz2whfR/c2HEIMjMhnPQ
0j0sY/90CdinrvDalWmnw9acHznUYtQH3zOz0PTuYgb5ItVCrLiKQ12TQ42F7YegXLck0IkUqUy5
69jdSiSg4CxsdklLtHuF90+plSpASHAMPkTATX0kRJGIefmcYisQ0Fy4Bd8CgwzF84rcA/AoIKZu
WRtQJnZFlKKz8Qdm2oOB1z0Mm54z7QY8V9pIp9vMBsSsGY9u9eDWsryQePxN7hMN4VgU12YgUl/c
lAti0ZYvs65xAJvpGCQsSJzWsLZ73pAsMN08ghr5m/QTeSPJ7/p9mGjvAZQDqwoXiQm1BEMA66i7
yiHP83Gp9dkkSeyLRhFizbzof/S66f8UOVzE9svct7qHjE+/zOm4AF3AJL5bxI6YhjZCZF1mmq0I
u0VPDCo1NYauhBsQVQ36C0HrUnfE59eJ8bUrUOm8NAomYnB70nc8KMmxL12yrvaozGlVu2gpjME9
HfPuLMkz7HJBiswbsDq3A5wMA60jkgy67uKzyRRu1M2a0KRYDb7CLqE7WPvr1GQJLl34WJHzaPfQ
KQm8ZwIFxbRxZCzaps6FdrCtk7zcOL62lwEyeYMQgb6GeytsmD/bpBYqX9QC95ohaYvvnAPmG6xv
m7rsJlrI4J3Om9UaRHiTKazrR7+k6WGjq0uj0h6mcszHn+LDjDkwAS/37eCNznHmpvsOorm/qwVk
ueTWovIv6fcmckNS5v6IjRwSmAEkVvzFcFnko2mu9G+OuFr62p3X7D0Xgc1CqsF/HBus0zza4dcu
21eHVHVSpoPU74mkG/S6W6THOemeajJF8ZWSBHyllhGsSGKQYDn8YH+UvcFi5QPrqodUNr4yeY8C
RQIXp+IBCgB1nG57NQhdxbt8vs7wwqAJIBSPWP18o1BwmASQ6cUqzeLcgzu+QCh4hA+48YUR7Wbp
vQaO3ZMog2eLB2FkRlttdxxRoiPYXJQioGk+44RbiiyuZC6HhJP8cjdG4oBv2P6wiWRQBZ/JrzfQ
DCzNgBgc1xfh04HZEpvh7Pi7VYI6IK0UAc+Cham4wijj0kq8Aj5Bm7hZfNP6CQQsh3cN4Zi/UGuU
Ohmb5mAZ2W0tLbs4zNbMeiAfNTRzqq+WKcr3bJOkFFJTy2FOcM+tGBtU4jTqUT2VNpmJAQRBrHhq
qbIfaUifi7hLieRr4D42dDB1YlyZlMpWRJTfCYVxAReEAawiNus1NYQQamTlKCSCmBvw0HAMzyzg
4+lZPUVS48VrJfjFCl+/ToUYTRPKf3QW0QAwY1hKauWIAPbj72wwUvwwGIk5V+8L+pI+zFXauEOu
mtY8N6F33IbMSkBYbuue5VKFAA5moK5QmR8RWZ1fsfUoBpZ3UCQwbghuDCZkRJoc8G+g934e2ujr
ye7gxNEceuEPx2jhBqVZwo9aUTAswOKNr/09q7hZWa/Mce3EpbHskc42pbEmptIS3NjeqpsRBDf9
HvGK3Q+P5hmrkV6pNNVYSZ8GCBX8YAp86CTXTs0v9sGw6mfv1MyYIRevFfM61ttDmGtj3dvmN0b7
BWcYMnKD41iWq5uEJp5hUg3V8oPSqjlbGF8VbDV3ltQyVvRg5SaTpXSNkg0cm5rkkiqSKoN5+Ro7
rqqoIaVzJJ81MvwAX47SkAYn3LsytRAhSP4qKRWoSxOFECTK0WJ83nJBN6qb0z4BHyCJeKsr05Py
Zv6PO6cvck87ljqwJVKW03gCXNQ0ti23GHDwy+EtE7nulPzkB94bPIipHfOQ+hSlwB4eeq7KlUN5
aW6Y9qTu2oDzOuOgj+sOVwOysDp5LFrhUXnpzaD5RpWpzZsmPZkd3ajFCUnOkejPmdqC4kjdqf+J
bAxTBhmcMlXH+pb8ahP4Nu+XYYAlgh/DF3EE34/POrPrLsPNXGX40mcaSP++auV6mvgXkDMCyISZ
qvNZrOChSkMyDDrHgNq5js3FcJTSU4U/CxHx+bBFLYpRp7lnmvuC5wswF8NNmH/wpVRt+zvg3Nf8
EjtX8hiW3ZkKfsI5cLMvNmF8X9smaY2IBri750OR8RlB4t+eryKybWkyKpHcmIt6Bi9aqwVkMPDC
C/G6isSgE4jUlR/IUrpLkjBlupUrQYfUAADFxf/djiy9uB/GDQnv3mYnR3A5Q0Y4+3wZmRpnLpuX
UScM63nVbHwTxVdbeCK4DF1b523ynfDBh2JNkTiMGIsNQsodnMw+86rvvjFFrlGndeScd+pxLE/d
TUTCnebOBUhnadT/4xv2FGQDpXGEHdCmbSBrv2U9Md+FDqUSbm+f6CnR6jiZMPaeEwQt5wHI66RX
lvt5jfkiNzZhj61CSl3smjgNlGH+cDSltQ4nBiyNG+RQFk64nSVshmQ/A36rRkpTrRbiIXNS4onx
aAsMdmP49B6m2CzfUemzeZkCJZ1Kt5HqY4SNgAXXsrTtQ5bBDBiUXrIh9ko3RTTteHcg9ZcrXirV
KudOq+f/SCOupm4OCL7YV5NXRyH2/Bc0pjvPDH2OIKPkxc7lYEPzRzpOxnJ/igJd7fXlIJsYCGSu
/8KAW1+AQJC95zw9/rqu6P2SBwxQl37UFg2+511raDYa/bXNFnEnr0heAfDBszu3FThkbE6oYMHq
mZK0dAvyL8mc5Noe2/24oGUMGjwLL8FQQV5yalVakxrRoZbdq0HcsWaMvKYUucDp37rFOxmP4dRj
xeLbSSrPOKTg7lz4PFmg12s0DFdkkPSN6vllea4QhwCLAta4zYyF8p71f47/7nl3dVgud0VNYJRW
inU1TeARKJRb1LM9wDfLSpcpsOxxFqLdl5vADlwxZ29TOw0qKcmr9TXA0JOGySBUdMWGxlq4z4e8
NpAdOOuU2pHVZOvWRmFPJ4OGBctUEOtzu0Daui5k8H/TCbdK7JJuKDzndH0v7LVv2YJ6+AMJF3w2
maS6Qtqlp17Lty6hVREiBEhzc31UUhNNO8xnmEtnIzknTVd2LRDfsLGXa9VHO6kJwaF7H+z5qnxA
uXzRLGll6c5VS/C7Fp2Er0cY8hlWOda5zsXb1Jgli8OAihpP99AY96U+Wz3iLHK2pZB2cDU6Em1B
mQWXCpXBcBz69sjg6TEezCazM7wHDJ8phoSk/yb3+jmVudBqKfoGDQfRHQMADDi9Q9wwScS+q5nm
qI2rE0COXXEicVqo5hDpRSzfmTcLueuCgBikJ+wuD79vTnGIH2H8PDjYF6gj4zfMeCm2EMejWIbW
cT7H7+481mSyiqlKYnDYt+e+nosNJxnb/KumB7cFyFkqRLlFisZJdEKb+e/jEEp0HLKuCJ9Vrdxu
I0IdHmLYvmu1Dv9vtxDozzCp4QBUqiI2lAIlyM038o7vvDIZCGKOknjsiwKRnJbl5MsOnXQ/nxQv
QNPf5M64Ph0LAKdKYlqfbxWAk8Qdo9gjDSuEKA9kPXL0pKRolTt4Hjd+i1Aq7+A25FiUCUUA9uCv
FMBxipWs+0HNqQ5HX6dFqP3B18YIzKYFTCCCHqEiI9smqq2NLv/LMJ0ZTLoqRqbxsp2c7KnJ1Xb5
J/pyZs1X4uOZCrCLwEBKyfJfLmRIKx2Z0B3NFSnlfzzLJF5TKPRtAt9ul0wmAozcqOEvDqQlP66/
+2zh8p9fqeVcl7BNINMnOpWkLdm5UNSkYWEKzjjiCVz1W0SuL9t0VTihv8lZIR9CCYSz50gcdgzg
2U0RBFX8aA8uEDqTixn3evvZBG0XH3aw+NGB+nEcFATeSTKuOs1BuamXi8EBhTFVh+O3cJNMsgM8
CH365OvBCcHYr7TbmQ5wAdM8x3t2s56e0/8Ni57w8HboGD1ZyMkPUCK+QTKkvJxmgnYUTvQbzt4z
gOrst7ZDFfFeyrQ4ek7FbH4zhsYWsxu5HVmEER1jfhcv2HNKENTLTMFTrZoT44C/x9XE0Hdrjvo3
9mldC9dLOp+XcmbnPgR7JvUpdbyCBngq1hhYWObj9PXkglXiF9+2L1Mubzt7CvaSjx+zyXgu8xT8
yMQUDv7NYCg43J+CLFSPDf8fmnYEEOavgbD7qfgbXG2s3dWkO5TY7FsUNFNShlMDO5ZVXzvdS3oP
iuajayM3DCzlQ3k7XdBL0kya7UC8uNZvpOXSja0QMExtwmQBFRzYpLEh9NGWFeDTA6i/G33rp7G5
29UYBTGoUCzzhlOCHSrPTpaKPeLr+IaPgoHnA3jPl24EqzNGUckh4onSlXUH+w4Lt6s7y/eGc8p+
mxcXVbza0ZCBeG0M6673nSpipejC6Uxu/cziglIvleJ5mP+CQ8gOaMvCTbX8957g91a49DeEWTHH
y1zM/vwN67z/amPtJ92YPpd7A5WE9qipKLd7rKR27L33RHaRWVA0TNQLq3Pz7R3mf3F8UZqqDqNP
PItQTDq+hK8JRv0khPX6kTDi7bIQZQzDjhgyWS7prrFkeMUzmVgUJlBjO2r8v4J+S16fOAumsD2H
0Vm7QD3trgh6vV1CxyKz9EcbobPWlvp+gstHzGmX58EMUowJwhLUEUTheMdNmqOU+bZbAZh65iBp
MjB656kpwLqv4Mrf23jCkM0G6v4jN/FSQTkCFGnTMqzZLVLOrnOkRdMOoU/yvUlsjcMno5E397Ts
L5ledJ/7MWCZbrRRy5IwUhkPBoj2BS5lmRtNaY4akllt37KA+LbawzSQDHkrAivufX0p4s6Qeb0x
3ZchN3fRhnsFzdpOB1ercO0K/AT/iRWFllh0Tgj/1Xo5egqVNjPNLy47LXYy6T0eVo2W3tHC0KWm
wrPSWN6p5ONZQ9u9W6mpu70SYnhU7hayxkQp9Ycyn05RL3E9Vl/Rg/+JQSgUzXoqaZ6KQ3Z6GiQP
Sad0R9LjWAUJipth9w/HjfuyYjBTtFyfrdHRgW/AhjeccNlC96Cm6wdEoX0xg46VK6dXhyUmhY7L
97Izlpdv7N1uyE6W2f/kVr2KT2BQaYppFFKbUqmerDg9S8jiN6qbeButorcxq67KljtHUMIcbxiK
54C5dfmKzHxcdYTNheqDdI8ICojXr6qwIyE+9FKo+hZHYkSFVg3dMryNhHPWi4RhIzNzWxG4CqYm
fkG0uZyZxTVLNF6aZAQuytZCY6ILGzoLIQEeljUfryPGDGO73t2s4DYGi5o9p2ydKGHils9KpGAA
3jVTlMi+5yG0GPv9mFO3EkWIi7z3ZL+CP3nviqdsPnPih5GHo5aYY5R1ldLf0+vjviw5OZeeHElr
cZrK1EDbX8VrNMEgjGFn83mOAf1LDyz84vu3YHykD4irStAZZ1fgB1Ra5EA9T/AWFSqFf3COj1Sq
wciqtTMU4iR4iyboRXvE4OVDIwSA5eAwSswloGOtA5L18uNBNMCNfbPK72PCblGOUyGLHgeA/9O4
u+TVlQiuFMDc/kzjk0JGpO/+oe9RRKvrjiKVhcajF8COOpY1U24Y/U92KJoCe8pSnlzN54UMEo8D
+FpKbzJgc1M90N/fCaai1FNy44XH5GucIA7yjFE9ii1Ztvl//Vub+kFSeFEZ3jvFvGwtdXhD5Uz9
Sd2oLl9U5249yiIIyxZRkTDjqFexrnGCiuJZHNNpbPwRfIm8NGX6vLAeciZIFQRHdz02ssCdexAZ
ejjbV9sxyBtb41GQyY01fSpkvSOLFxvRRaDhl/sx4haxrEEiU3B8GrEUfNLpuwz5rrLm5nnYwh2Y
us015AGGs3jLFm+LV1jdkZJ7kf+GhaVA54AT7ycDNOL8HkSyPxOWKAzLqnm7gk3o4B+Asp4OOUea
r1feiSZ9SbRqwxUBHV6rLD1AUeiqz0L/BEHUp8+unKJa4nNPu4KW9MW16FlmNk1jEWDDuUJamf3f
oRSeDtXuMLnRP63/Yvq6Vi2eBZM0VO99dlg+768g7sejrMKGV77U1qK+aBaYLkVQmvsqh/6FPG9a
GdOlmnA7bn0WFuOjN+FNHl0GVFmzDEvFDHuL75w/gp8rtd3ED3th/WeYrF+UePJwN8Xn3u4D0eum
WacQXdZC41L5iDjpX0M8VZsuIaSsrEoFI/IhAvwvVtYdetBtYDb++BdtpU6oSpm8VH7zJ6RuKlZS
ZR17nWaJ4pBIeMy6kM30i0RG2TRXMh/m9InXCElIE3FKBxsx5xsA9HWcolobV4hzfGLIhvTXx47L
/J9S/lBANEphdT5/ONI2B4KCwxWe8Izzr9YNzDaPCFui7nfNghDU6kzuJf05yOTw5Yeq4eBGM7p0
+e0y6A39iv4uCUQ26s9J7ztd3AWYusuWg0ptMywhucTsxg6fA1lOEdPsomuRfOQwpRuED3a4A4Qz
GhH8P3u+IAh3DxQo0+E3O0Owm6TvYKnd3X7Yy17Hb7Y98uut6oxo6YfMjfh82XrUrVYuXqa8Mw/h
JQcpaEvebf79HCLl/yuIP772B9z8/dAhm/W9ma4FOWyAfot/i3C6s7Smt18knNjoJPCibZKHnMGJ
uvlOiNxsJ2iito9ZVMTQhiglJGWU1OEA290uSQVVgkiMPMzmibSLqQfIUTgv6UB+JpoIkKRn9pYw
bNfyubBuEVaJ5Za7x68Esl2d+w6a1w7iXj35jjYOk5utAlRgqYkOuLpJc2LB3k+GK4q77hTMQpS2
E+OXeU+pMiqOy+yRsSdv5y4lnETfldIi65wHfzUmjnOQphv/daVJnvdRqf5rSz6iwSTog2cN7fif
TWqU/PCKsaJ+JzJGwc8Ci+4HPZazgbdM8RCbFPCNyOND7SKTATxyuozZhGsezDPFiPjn0wXbeswc
Ex+zQSmKK4j2uzDjTbBrZmjEZqqdSLmtFpG68wXpCGoCqb0PKWZzK4vqg4+SgyUcKo3S8xFnB5GD
E4lrC9miUKukD6od1IJgSixtOIjajk9RZvKaL545nBCNtA6stBhQ77RXe2MJoOjRsbrtI2SrZEGN
01lkKCBxwz5mmSIc7QsoGl34t9MMIyreiL3AQJKLtjc/UAr3rznYFDtAuG15zYPOiu8SbWxwJKaE
LQIDpZTEMUprph+q6NKX/9eGvdCkx1KIhsOZsCuDYNc98H6/0jb6wiLpWxjacJjAgCDd8fLNVu3s
Vs9yAnv2R+wB2J33eEoIQ3iPYDGGEb0q3GITJ3SBQYYNK2jMv3QvzLhimrMMcnww6/g7s1OFGDpC
woVyPjqeXzR0rRk4g6TRXcTbGqG4nhmzhywNF4spxipbGSG8ForrnEXgaSY85hUvyY4Ch1qJ3cLs
Edoe1OI7IdZht5OQJjU6CDrW9CrJXU258Oj+isCK889y80+GTYozzAIUkyWmUzsoyJF52n6uv0wG
wW+jHa/XLWq6y/n1kfhO3gGkFZJCIzpbuNzxhf83hxJvGS40YcHSdg/ZWVeAFD4LvamjVxjlN9BT
Heq1/Zj2Qc1YFBQgy8Dr3HEW5xxwEmLWxHqxeSMwyYKnj+PFhC5fBJLUcqR2LjmKcDecMGUz2V12
Pk0d4NAXlAW+i1j41+aG1cPgbWCI/2cndkBDWKi/Il+Efonu/uroaImEeoKeU08TS8Pi74TjDZv9
DKjG7EtRI2I8hOqKZvXD3GKRuT78HZl3Yz2BRQJNx+2ThJTPGBtUAOV1a/QUx+OxtMFVaSITcQOu
R8P7A49MgGVmWTpeZVxFSfOBw+ZvxRlQdhk+W8MbkROQdEbXbW3KMU9BVbpp7XSTxmSu2c1wlCTY
8kTGTkQ4T41a0HJtijRKBhNMH6eguAwbGDvQOVeKirbdBThYdaF4wJiLvYKVfghkJhx9WtvffAb/
nzNv/FIUT90fBCuJVEP0hGMZ3O2BaLxmw3P0LetlwXE/aMpZSyOXw4nwfMEzPEUIJJyDE/SprVjh
ivk3qHfNq44VgC1MI0LUDr3Pzk7FObjPPLYrhVgRq1vZZY2upJuNoNJkY2ERFXUezIEKvZpa/cVd
UlQe65+pKLrtSutlQ8nCmNonE+oHTaiZrKw3r5OzloBwVJnpYbCzSYfoyg9Ydy8sRHEawiscIX+P
Mpg7FPJwgQlFxj3IN6UcQw5ISjbzeXdd/bIAGcjAzcXaomXJ9P9BaReC+UTDXL3I55e28XBaGFNd
xa3FXLcrzGyvGAE2+9934b65105DFLKS8UytpKtPt6660ScNUOo9GTb6D7hirbIWngj4/P08m7Qn
qQ1r4Mhvps/64EUDjiwp8i4dudR4HT1g3ZRysuhG9Sbsi5yy3TmDKXMZbtmqVmvh7XWDNlMzQ+Z4
RzW5ArbrV6zjkJyvl3DSm1vRZcIPPjEm5TYEUtvqhrXKX8JceCxYXDj21z46U5ta1vYGP4vttQbI
7dBxw6oSdo/xATYgPMKL/YN9tnmoMl5AXoAfCHHcqnJDtIGHx6dZQkduUaPNhvqY4985TZt78+Vt
0gFYJe91VDcTK1ljgMCoRgQvulS6tyeRt/L9pJYZUxQfdWEfLNus7Upbg+KUWkkLUWs7YUVwzrUK
muODrqJP2pBLrJxBXdF0MhBQSHafcfKPq8cI/tLiZgNHIpk0xHFHDme0EIsrqIUA3wNQUBXAG3wj
KGo75No31VVI2FrQ4M/2FNrw0T9C5kB1wsuQC7oOw1g46PG+WDNegUb+iysLS0ppkSmaxY9gPYnF
ywhHzgQQeUm/7vSnYHAGxXORncDkfFRIvRIxnQygNzPbSP28Kyqfbpq8ahYAi7Xs35iRqI2aVY0k
7AsSN7b142zyXM31wOXzFBQm/cEvTRput1EcKIv2+An3yWm6ikwyDyJMlJsSgAarmsq87nrymCis
gSrVpRGWDCKnZXvr3UDrqKben3Z/XE+oQr7UJ6Vdu3c74rz5arPq6Ybo/KMWLM1OxmRXwI2so/UY
xClE/TSxmUl7QBnzxp8ltITNLV6Zuw/h7VY/2te24iDLhJxDp85ZluzoZ9ULYryzovjql4o8cZD4
yIyVS+Fo13KU3/00Ae9VLo7SdS+7T8k7zBn58tt8sg79w3xZioJOtV63eHrfLS84otgl+1F0oErg
G9Tb+TLLIstIfePgSAmwx4GDZpiluw4fmSZ4BfVqqnfRKiR1tLGOxxVUWui/boyhIYGo7sgJp2du
Y5YvcyfcvWWRfnNoFGo7z5QjFmRXBwNBLPkB2cgVe2YLtrizTyUBQF5YlI/yUciPiYXaW6hE54aG
f/Ff1njAodoyXVWMSTX4Sr6zRsXaMzp7mTktp5XHN9YOFyhyK3B0D7wMPKLAtVjQSiQWMWrE1ixy
1IgKSkmANnLfEzC1q+1lgd4IzMtdXwO7SQV8YF5XkjEWAzG8lXdGXe8jNunTePucgJvdvPqnPb+N
+vuN7QEkB6zsX6KgRsUBV1NOyIFP5j2/eWOe3xUs499C1wzg9qQrOiizXyh71hW49+kdOzYMtwFL
wLIUeDIdDrZNKkvhhzSEV1/uLUjPz8ThPDGhXT81XuOC/kEz5YQ35McGLZC39fASQalBqVUY/JyP
MQB06L/JPBNcehl2G4lTXkGExzsbq5KPAIH8ZMbmCzFhDZGg3B+fTD2/6Sjvud2ODWXlppevZc1J
LKR3/ZOkIO99lrYY0sdzEnxAZMb0RWYQ2BwRIogLiGsbdRbHmSpe1I3D38ZOtqQxfrufgtr+/3W4
9fUBXL5aZNEkhEoZQ9fQBdsjmauid3JdPLXLLaGFBGuitOtmzVm1kbOj0I2hlXXBdl4VwyWscYYt
Xgo2tgA496Wz7MrnCYshq5PDfugnFkRM2l0TrAsbyJW6osSNOEQeOBi1bYBEqRBf5rp6EbzGHcdk
yMrDf+dPwJdB5MtcsHmwPAJU2NgL/02z4zs585LGYMb0cp2BsG//UKlnZ5eUmjKo7wGz9u7qDLc8
jCQ+7OEJGiXAzfd/RJvnqi66sqG932viW1U4N6SKLNTtDXyy1Ts1Q1JQIuQ0taqI9cMbmsXouyoF
lk+/mDFcC9XOT7v0XKlZe9sxi8AKyF0m//aqFz7vHesz8r+bMtv9cabSwXT+Bhvut1dfawD9366w
ChVStAvuQYTfiJE11PFst4BgKCeEoGwKBv3gY/WiQwtN9O/7oJBdoBOISfCI/MxZ+KHjX7cfUVik
FPROnIwHEK+2vkX1qGtXY2k10s8/nkJ24/XEpwXQyvfbIWV41mDD6Wo/3WtuAf0y1NmYi0JXDpdD
lctmxMItBwe4bQSmNesVfEeyTB6+GKvM9DysMI8buZPNXBFhZibyNbcuG7RvR7DixwLdhmKM3H/A
gmxbkLbx/5VBmxGs3F+8sAKUETs8goutT1K/4GFqR9gTqRCTU8kRnDDf8mj3bWv2tXCAWPiZ2qsf
jiUmDCs5v82i1bga+WMQ4+TXvBGe6WIqNHUhWmt9ZFYPcXHVeo05Jr8UMVEi8SAi+2erC/iMgNAO
Fcuo5ZDk3ufFKSPGXV+QBXVfyzIBKujGfZwLy18p2Je/tJsn74gkjB/YTgAXPfu1fPW7R1fkVo6J
aFKDzv3tq40KQO6pBawqJpftGVGaf7hJ9qsjGENoJF2n9mkMwjbLp560CMxuoyZZDaPz3jw1w7ve
X+XKDVEIIDKbgbzRJcG8CWm6htNDOdjM3WdBBp9csjEBvm12Y8H4S8p5UcZuriDh/4C5DoHUbHPI
Ofz3YrSaYbzd1vD0VIv6zD4whMHWkRbdTtKYQdmCZTwxkyphfiXJUmQSenZr2gOJ0V+rG4SBZQpl
1MVLEaBqzSBVGVeoUpzd/3sfejN+NkDwiYJaromsrzoIuwjCvXZ8ocy8dlOp/YVZArCCgcvz3rQV
d3O9B9pgKm4tjJQU3ga2R1mySJRAbnIVwIuYr4SnLzw27uAPp/XtlkCFiUTbXuYo2k3MQjJG5K7B
hOrmq5n2V2Kz39SboJy9pT3EK59plzqwC8atOG1TORxXX+pltSkNYZGCzgfcRZtUtLRdvPo7sHOi
s+rvOZAlolto+RjeqN7W16nEt4zOGAeGEmyf4GTcjFpiIIFCAwqnik7AoectNx91q2PkzEXfGWyr
9KQ17SjCKLTy6ZuZxOl/tbRN1gw/i6gJDXPne/HPwiFtTtr5mJDglvpKqSDnF3QMFpu9OOu+xQLe
EQ/u8tgZfR42iPLXEG1x4BE6/E1+kmooPwHyRVwxEBofWm3oYl98tqQq2qpoDAM/qu+CwUg6hGyC
sOsO1dQKS3wYQG/1yxLec4da5H/hGx8TS9WRaWbbaUgqB1PicbYq641SbIoczhrR8zJr/RLbcWe/
k2iLm66YbemzvyRBrXLYPkobxBpR+pcRK0nv5Q/+gV3+LV9tARg0/GexqLM1+q+Lbnmz4KciBA9O
XTIMbIF+2Bc4wLU1+865kmyFmJspYOn/NHkyKJQeWA1+wN3uLn1tVO3IMeEoN7OKkI2crhm5XhzB
+D/4IKlmLIeB46yZjw9mFH2vh4B0PdUSQ+KktU/0b8Jc1k8scO+fqJcKvCoBy3nSLpFCwaryMROE
veYP2rxEkwGVHer6JAWnz1HTl0Di7TpjfvmI9wPiM2RKMMCUw94aqX1ZT+8r8QP7E4Y5/4dIm0kY
tMVU7AieJZgoXrlP2SH0xNf+UUkMER5wCWbiQ8jTA38b/mkGo8oB2PHbEU2BCRoQF99+iHbNKYMh
8nik+r433tqHYlZ9aEnjBvzzbx9J35z/InIcS5sqloaHMSRJYb44jEWFttDAAJ0FpdCSaGN/Ytx0
A6ad2TtFVvoVp5WHchZxf2d33Yhpl620Ssrl1f4PUQMgSLQeS0PrQKmz5ve16uDKaaRnKOxWOjus
RplYKh4I4/B2Y92mfZg/3AxaXwZhc1jkCxroW9ta0Z6Y9JBewRbLol2q32YeYRSlzWHXVcMRfe2Q
zNb5RawTr/tFVNCGpOJjaZhVsKi4u4EyPWKFnjbA5VxOhGfiJu96qy7/5laDV29gh53kDhfb1Gtd
y+C0cw84158M2SvlGngz8kU58Uep10HqY43iOI4QukOpyjS4bV/Ur1afjUDfSOoISaO1XDB+RbZm
z6zSR36Nktk4zX+3zJzw6vRS/rezYFCEAdzw4fzk4CYGHUGd4xppRCFSuEayzL7EBO8TrZ6PP2AT
9OTdNDrKjsWQ+akePRLYby7BKl3sDEhQpUNmVmUuLMfhrpS80J4rd4XAKq5l+0FxMkILMaVWzS0P
ugOK40S2i2X5jdkiadZuiES3Bli9BiUnuSSNU1/lJHYjaW4X7PV7iYdUOEr/6cY0ONljkTHF4DIi
z1dHT/+rvdItaVwN2cZFHB5OwsYTSuZXgTvGi24B4DPQTCEWgcVNzrUj0dsS9upvhjMmPKmGCHAE
H96xIPlUaHqja4siPiWcbNGb4xzdyLnZOOKxKy0H2ydoHlYrig0uMdWp4gMPPrrRoueT93qeJgtC
Y1Vu+Da/8jEGH9a+fbjGseweZ+Gz9rRzuYpfBhxbbHP/vDMaQqWXjpwnaOCNUM+N1SlaDN5mjUVF
QeYmkp790LIQ9V366jjCA2snEuPJ2hkMjl4wWgJVx39j7mE6EWQ+69vq3hqOulFvIbuKxMjMuxbP
559VR+0Dfg/JdgvP4eEFNzaskH9JjcE7ldE0pBPTcmNFsTUtht5k5qkwQ6MitzxQ1RJzke9e2TQm
wkVu5SmJhXKBLevB2NspxusFHGa7Ycz3W3hkL48/+By95WpMr1vbtFP8y0KU9vUR/YZUOqhW17c9
ngZipsE/RnCVo72N1VXpv9bzsARv/okLKW+1bgnnqOrJ+93pDFUbjto1jdnNVTIF6Tle3bzQoMMa
N5XT1IG4JKUOhseyCkPemAZccUk5VZx0ss4EHBCDgzzsfYjFLLqNJbxzO6bjAXSXWM6gepNm27Ws
Rb1bnsBUvCY2HxrRVsvBb12xsT7LvQJZRBp/JJFUCVNk2BPZpxDVHXzmZsh5wlpYZ5UsymEOzrgJ
g9zBCz1yT6558HELijfD7olZbBITOzVviEvchofBzAk53CbZNucfKAwkzVPjZTR9qh8DCBnTtqAJ
grVO0/rir8YdCmvpG3541mZO0HQB4J+dKXeImJrHMm7RYQNzQqRmoZDYTxtfoAgLsS6K2wnWQI2B
M93yMOzktXKQ6sL8rj169mxzS5VpppAJx9L/S7fGtiNBoJHWrsS5kUzVzLvVb9QfVZWpQKr3Fafi
RCGhrUQnrJJpdqFLyok55id5t9VMNq1bGEytEO8Be233FqTmw12Cq4956g089ESZHZTOxBGMeqK1
GClw95UXpYmeA96CtKGCU2kAxq1EuY+gvOK4h5kDrXa+LUYVpzYlg6JOeeHqKlHiSpNuCuqDi8Qc
CDEEicLYSlCAavr6fOoIfxfOSNDISGzvYpHeoln7USkUeCUY5+zqXef840LYh4F6jrb0tGL6qmqy
VfLlulFHJu/YJEEGH90aSC/kCJJTDFPd8pjYlkn+nd11d6IY0H5ShUcS2OVjYxUsbwXVu/fnwetY
UDVO6lSwpJxlm1j8RiIufVM3CBOjeuDhelRB+W4jmiQdj2dqXbBkH0q4UC3yBIEUseEsRdLTh7db
e4MvlrUYrqc4a7+eQmvY6xgdBL9A7cnMNzsRWgCljmr1NsotYSze9J0C2h6zrNsMOtjq3cor9wQk
q3KC1qxlj0KwV+lmUsCZBwzNDY/ntgcF9wkx6wTdPVjV2AKizyyA75myLgg9zCHGbJxAmUiLfVq9
a/p7reEbivYOZewn2hQTbtEK1DYCbzV4upFjgH0DmWCNHQE9kfptSEaNxHoUjQS0FKQ0VorrxWqw
XMB/jdC/tdK8hZY29zWPcPCEn8wxqOapgEBpBtLonuTpSNPiWrhLYJH7V2El1i8eFnPKx+WxkONn
FeFFQ7DoQ0PDOvC0Zhm23SUXJFoxizrdUHCTj+OeuLgCvRbOw2TCR1ZAjQjE8GpIcup8b2CeZTod
1tIywLSEnMEjXgkpxsGcmlstPqfO0AsCUod3J/6c8T8qxWGj2w6Gp3Vjnq8y570XqmjKr/RwsAmv
BfoIWyDF6pKdweWgBOvpG1171kaKyBSjkYB0DoGHRJ+ZSdmJ8vPWuosCe7YKuMaTjUDbTnvtsih0
Y0eIuSF4A3G6qwlr/o8EEiweKGOUzEcClEDiiEHHAKzJgDNXQv1K+5BeU55OddKRfffAGLiGcFq8
bsHtTD/x5dO4xULAJu9gzjTNSdhBuOOFWqkCeeWjBu7pOR+XRn9omwdPe2othtroVHzCZdGnNTTJ
EriAyHHncsfj0D9W3cY92cHfsauOfgsETOo5oMKkpoYDoDca2y1Xz4z70HrS6wndXEX7Vx1x81qR
NY0jMrO5j+jEkhtLoHp8OcCWxtV9mvjUv1VHTXbduimIAKGmMHvedMldchYhmKhO2T1RFTe+pchk
oVE0Dm20bYNYcJw5TOdqob1uigBKkA+ac4A3RCBua6wYcO+N5VzlH80fQ+IDyEr60JvlPsMRK0Z3
Oksr85R5ByJAEqUENy2im9VhASCMRsCIago7oajwMwCwN8EwpYvwZoxcZJD4Tm8zNJhiR+jqls/u
+t7yMy1T7/RBbgdtFjStOeqUY7x/lhc7Or81+gXd/tsaI6hTVL9KfISrC8H4cW5PcfZu628NI73F
RO9strB1H1PCntiGe+rrNH+S0qSlw0zekzBG96o5JYThO74yjjnFnyFEPxFER1UE4vYDCUdgTYPc
dlhIyYEWnnp8RWOsJEGRvbTSDWySsyACrUVZ0d/L8wtwg+gL35yAuhEYzD11eliKpvGa69Jt0gjn
IqoBqZmfyuVcRLBL/jgbKPLM+gzZaTQe+SDl7diaglKbxhokvg34s5UtCUCQ2rL8AYZPPwD4pHv/
6VfbL1Df6uUYPK5WbSsU/N32KR3Y4b7wAjIPoLt6XoxBSpDhFTbygXog2RQG5+avXvC4aiFDkWu4
XgYNBx2Y3KYqceSjBVYRIYYDbbC5BYeiNTNFtS8b5f77Z3Ma36s1gOHedVDL+VCV0VH2HNdvtbtK
qKfUMtFIHRB8XZq31EOzTvbY9jSgFB70jSZ8bbxVDk2laRk80Ab2ZfpclJoSUZo7Yqpc0t9rZcmh
SNMtSUxzSjx3GCvRzD0QkNUsIcO6cSn3EHLL8Q6m5E0me/46kpOMP3/6hVFOAQCsyNX5wEe6kvUb
hwMJOEpCD2fvsoIyzawHX1P+5aG7LAL747p6OZClfdICDl3XGCe4/mdXSJ7zAHIYbsZbYiOtbTMP
aaXkjyHLsYKKzmzGYwXgvRCTIZbaCY0RXQAvrx49GmBJzG6MrLuUu9e6+xc6sFqMTLZItzyu+/uO
Dws9iM7s88XD6+pfGQOLekbJ9bm0Wi/03QoC5nRhMOPmwRhSNnyjHxgDFJ2QHt4DmNp6TpUGKNjt
id4pmN/4TBSMm+8UVu6RvDlbJYfuxcetVt1hRbNHl07IFZu6iECRxKcPGmGCW/VPKAogULrs9QQj
afIoeOkFwKVgmd6Il+J/wUHGugb8OnRExHSKrkvcW+s3yM7pokQsu52zTNnSVx4ylOUlR42llx/v
tMDLn7cXkIX/EP78hshRZBUn7n2UXVce8Bhiz7PhmyCPPPykHqT9b8unFbD+0yfFVzBitPAR7gj5
4YHOjEbJfxIUeePvdtjMXq/Y7GY/lZn/kLJalroJV92Tpby8xx5mMY2ovO5eLFdpuSvCRghHO6pG
EAmmfxcSQFXUT9NFgCUrvZmqlPqmOJT7tchIxwtoqg50VdeeXPpYDf9l1jdAwaGqa7jFemwnRkg3
1p8XkcFP3vAMx+SWQfKn23Yx6ZB1wwR43xWD/FWcNjf/U3CEKBDO2gDlsWJ2rqUB5DVPouEgK8RW
rBK1RNXoLvNSoxxtyW0aSAehNH3pEsHB82HPYd1UFAHpt4c7yUk4InvJO/mLfm3C5UK3UGFRDT4w
SCv0/Wgnc1J7xzbOes0POr3MecmhzVAadqvpbs+xx3LDNgFEvQ9KQZwZQ1oJu61/wfOg9pDhaR3A
0+uGov1So8OCOoJc9/8QpZQ4rUzLNI8oIl+Epy4vhou+aXDkYhGCJ4wNvXDIgzHoItCwBSbumxxy
uTAhjbhdZpSuIbavq7vRioXS5FSO4B7wtieGQqrmKXr3AH1rRUqkjzYPnVDsIIGX7JNaal4HWlR0
wjKwhpe9OYPdfLrTWdVvIPRuzs9PZ8mZqXs9y6S37MaX8YrOgjN6QcpvSRUuDiHYHdyR7aLPDAHi
NstDd96UtnTsPhZ+UWrpZvsxH/H0byC8bYgVvWGiFhWqb/EZn8cReOESF2CeIy01hgapti+D+XKn
QuFIs2Wl6sZJEuJe1mdbxOc/ogIZdtnh3yk0kxRsbSWg+7V3L9FW96XZvNUkCnxM0ADotr71LF08
gx9G6SMFV3XnZhh4bMWus61BPjHg4Gjd46cRury+Q+15Zu7hX7/qyeb5YI+gy/OjJSkX1UjDr1pQ
ZnlQgFpl+WRyNdecIN9etKlOt2bal9xpkGqhs5W0eCj7rXzEpvWB+ETn4Uw0LLUC5YG7jAqQ9ZT1
LGM2enB3oPvAScmw5KoZRQtGmH4ZhFs6BrXzPQYpOKJBlYR8MJmNJGQHzYZr3U0rz/OmWgcCpxG3
raXIQweNLQu/JGeMB47Oe4ZwPGsGTN1rv54Iez7FZ5KsPza6h+xpG0/DcKsNHz0XoyFFZsaHaQ3V
/bI71niPAx4rhe1HmkA2EXdvTL2z6pjPbiaqxtBHFzwHRkbub01k0zu7MuCM43zgVbR9ImSqt3ug
Tyg7W3l5G70DjUek5BQ2Zw2ucE+MznjTSUwiSlyfevyIl/AGLv2rl4O4+8hs8ftpc0H88Q01i6xk
YhDClYEICcoOHUaPmlq2xZEC/phq2NTHXUcDLH8n4RpAlz2kOOnuUeserRO7jXiDFqolDj/5gZEx
GgY2Y7P10uXJ3IwfAKxm0dFTkDDMgdP/UYMzog5LTV+7c8EgOh1+sSknJU5sUW0SbPIEio7y5A7h
KQhumBShx2pOlDky1wVbO819t4lwoQMfF5JWZBBPoqhvnr6zoUFIx8oTeolvFx5qKmTCj2JeeiTC
oSvjgiy+uAsiXyxjeH+nZLF8Bp8oLaZgXPEtlNbnpdsDmGwJkojpzMWuFa5PStuCE8jhfqKk2ZkW
37Qed1rQ5nejNceaR6FhovnEndeBoewBAa8wSaxscbAyIO2/eW6bmH+1tCaKiI+aHAOcoEiv6s4X
AEcdSa9V2olUhOEchrMqinNM76IGOa55/y90iQncR8yp6MR6GlW2ZCPjKerZPD1cW3Pxmciu4iqz
xv4eclJERlS+dNPLwFKhp4ohIaQoM3xXBVUqUIdpHntydZwbwF5liNlBKt0rDWUqiXys0MLzGYN7
JsdUs2xVX9uJdfY7CdQ1zc8m0+s5CRCPArQV7QPUQn51/bglu93nWvqYO6SS4EhcsjoyH9M8Nu+n
SHkKh4HEBbmUXowzumte7CEq5zgiQnN64dDnxPQk+5rwmbWlOhaqktsOkm6hfrRcXHu2JZ9j/GQ5
IP40pfna24GeG9LBDjMjOEjH2gIZuea0CrzMVBMzG/n6hIfMRXhUaP7iQ9TMoHQ7XoS2bWZ35zN6
eVkrm56X+FRtsjKa5FXGSPqMEQOmP3jrD6GNmA+TJWtYw7yIxZy2wbLJ8OyVDCmgSPORrLoL+dXh
sDeXcYq+z4Xtv+cjCHNEfYXR6wZzDT58OY4oPF2wmTefHetDGBJsBlsmkRyP40bo0oAYEzps5vsr
VSr6lkkd3P98INfbXBafjyn0xEPdmoh5tqVAt91QDLLA8cvyeH9nSEwTPBkA4redAsLDdiwLcZKm
TqLcXmECWSY3pSFAstQwLKFmARmSluPDTnPeyjdoCTSRmuOrOg6Bwo3Zs4/1cjp+sVlgnuVzjNET
J7d3rsQuiCYV889Kaegx4E41S33VKeuLDo6tJBJisqYNNKJMjGstsX789H409W6NotcPnsC0uJXo
6I4getx8iHVcUz4RbJFFDexT12Ee/NioM1uvHgu4NvPZqYv9Clzh1TvCJphN3siKWH6G0T8d2Du8
J+DjY6G/Chp9j8j480uArllEDKlxqchNsfo0kIcvHC3cD2sMuvKR4BgM8UEtkUkISkr89vvER5L9
kwxmZtVlmcKI1wOLSdEkufxAPtJiZWU122APuz7FmLx1ZV6x4f6Ni7wMeq2O6EfifwG9HeFWAA/3
cPiaLN4z4CZQHixUXQ57xV39z6cCEWvqpwSxLGFlLbTc6Jy2tuTBB1Rga6u2bqbMOCKbqqEVJ2f8
w+ihT89vCfzH+Rc6UCVfYQbxTRUP3EWmZZE8nKu+dv9j1vZCWHdbpBN4k2lp57/Ah6cG5k+1AaP5
+g4QweBBruC3E9i8wcgeM4ysqeVy34cf67dIDzkDnerEk23FpyAXJZQgMPueBL+hYFeTAla2oB9e
Zz0kQx13voECCWah4fMGXYlqALd09TSht6L1xTQ6iUSKOa3nezOoXfkDH9NHeM83zJWS9G24wczg
FLs2tKluRHrn89WM81H2m1WXaDcDieQ3Af0gpwiByAfsCJGeWVeK3abdMd7aLRDZPEyi516HsC0D
Gxge3UUO/KS+8ju98ENX+9sTVKFJX5EWsD7Ge/XflC+HmJ1UTyjWl7Z0m+8l7ghNewflxVWNnHdL
ibZDjJA2SZNHFN+MVgEKZPanlD+3lPQhyY6jfASgJ9sYRExHsysToVLIhX1to8L89G+aYDXksYpD
XQAKgM0KwCj0p+uV0zQgTUbvdl0lI+Ab0z/1fnxb44UYx36INufMeJtmvfAd/wjFY3+BFZh2yUOg
fFDA0tRDgtv5r8NWGkxbP+AjknUdD9u/UrioDdql1D4BANtOVtD0Q+TdkX7YPP6gT/r0TCXYXeOM
tjXA61UV2eDIPc93ktRU11FSXXryBxMPyIkI/PH5Bn00s2zaJMOhk2oMef7JnUdTjCLtdqrk5wZh
pzW8UB/LvCagFOb80RiyEjSWwvQaY9G8dnajZrl+3I5+j2HWgfw8iShUHUAPGyl93TAZnnWDxXc7
vMoHudPDbIhvV8pjLnXpegqNMsqYCYm54uWrs21XnfvBOw/nPUbfJPLF7naZp5AouubEvB2HFg+w
hPZ1HlinHBFw1AVV57PrrQRweYj5xinstn21hB50kzcxeAmj6Ar6lzWoFNtkhKbxdyMHJ6lCQamD
yw8Yohp4URthEFvE4liSHMXr4fEnnuDCV7hKiFX2po0wDciOIA2MfaEQoXcnoggNJzAH8cSQwkqz
nQtEom34snv3ng3FkOI2PAQbYCrUIzl1MEwsjV2kwiqaHsn0oq9wC3MvmnqFuB4BjYhc24hFHXWx
ngarHdqsGLToW+3OY8E4B4LZT/GaJgOeXXgdqKoPIFFdWdTH1N/hqsqBE2s9atHygxBNHf95G5Jh
/lTlZStv914r+8O9AVswTrJJrhrpAWVmfjmkPb2/PaezKlVpyBQL/gbLiZpnONdO2I+/iFVsn0PP
jdoXyqOD/UDKJIRNLjX2xH8EGxWLBjeSl/nQLnXMLeG4DVhSrlm2OU4hOgUnJZdXK+7+ePB+XvYU
7AXSEXCzGJOWTGtkvClkIQZc1EE+JQSXYZbw//zpU2oq4J0K1ETtVciw+ccGJFl+T8kSqeLnSse3
GUIzrm7bjFZE4ud2rmDnoXlsjWzLw/09HRRU8K7Q19YnGsG0lJobUcdJwie7/WZ/vrVhoCqd+RHs
hvXp9T99CiWnsBmAjKz6qMjSWGuPOa9ONM+BU57Z9AeZ/BjXgkX7fx9eAIeKbWAAeGw8E18qqIDC
H8M1KB8lPWrQxToorPyo5Z16n7WjBXXTL6mmx4+GyreKeNnQFNr/G3aGSeYfBlvIponEeXmdFX9N
vX+e5XcQ89aVxAjRBKqICywBWKLE2IILjC5ZE7lfpnQFBhsvZNGJkFVN4dY5ZWFDExAyHB0wnEIi
MX/b75TUSRyNvTtdm2NKFJKUYWaRIGPF0i3SW21INXy+VxeEX0Gqj2Nu5asAE//DX5v14tr2qwev
LFS9z6TVyDAblHXaqgk6scOoOuf1rABXh9KZAIL3wJySgJ2opDsb1VuDFoLdt9uOdqTM2GGEF0FD
uZh3Hqw0+3i7sYNjCg/laXg+7pI9PhZ4LcoU+QbO8KrsWZ9sehpJEIXLww3AsAwZDhEQktlEkqFa
NpzIGmM83VGp2XNEFL228y0rZsVZrbYa0yEkXqTKpqSYbnR2XvTte58C9TVu/zhieC14ZOmUPq1U
HdbmNe47psAWeLxqHpD7gYbEI2Q5a4Dgnl3jN79KpobMyUF/PLMUPuKP39577GZl1gQBDF3BwJ1h
0Ds+fsWZQ0z4RjRY/YdhvJxAY/vZ+P0j5VlUHXP9OLWsgu3V6MmMvDlfPE6YubmVlN+mWkPClb+B
V4qqyd6HCf0OS9RRXM9ki1bhw7tfTtq7cB3F21QGSqga8vNBSoTmAboRe+s76tbma8xlq2itWBVr
6gPzoqsEXHdAhNge9Yk/90UJoTnS+X6lKso1YQm3sAb3iTSrdwFCFb0RmU3ctt4mXecMegxNKh5a
T4AX0kGvofgumqBbNlLWjjLIfHaaLB24ICEn8aaDCepof/S8f6vqitsekFfe4xCWjIDlIMkXGAgK
796GGM6Ckvq13smOTGJDkLwoV0o3eHEzrJXBX9802G1bEeBC2x2Lvi+S5hw2+fFumCaeHodYqNAy
F0jVDJi+dyi0cQFIqOmVnFhAaLP9/t4uSlIfn5MDgJ1rkHtXBX+zullmP5HyIFffRJIvtAZAKQC9
15XV7GW1IKUSQEdMshPoAn+nCtk8N441LF7aSpbAE2q09Gr6YgDMWWWG+TjjavF6Vm8WG8jmldrE
MDG86y8LxxkfxhoqYjScLmJKTZjhOHKWUSkDRLjmwGNuW00+ymdw/9PNrgE6Iueek1Piajd5h5pU
bNZq1nGawoiIHU2lHLZV4xoO9heeVW2iyS1V0LlfFkGlIkhCFiA+6ME+7HrI9dn9LMqdmffjNlBE
x4pP2a72VLokZjVTsk9nfkWW/B3k1IXwsdrsNwsqTnPLQfyqPmP4OMQXi3GHCF3QnQH5aaRErZ2u
/0+JIVC670Vy+qxSaVpmCBOq8c+srCVpHmO25YpGkQXE8oUDZ2w0wS9ppPLMofQD/dS625BdKHRs
yA1ST/0HgMb/vSgTXcV/ZSvIJ4ZBzvF5lBiJxeDJ3+Zbhz6ogzyQaiXZkFDCWWf+raQzUxgQuhHL
Z9x1x1r49vFMc4lgai6F5y7EELMK9TVwaqakx3tRwzfuyh2Hb5oIsqsuTwD0JOr0b4D5f3ANb33A
T+RrS0AlvkCnTJRpctXoHXpp7zI7sDf78VZ1ylKgoJ+SOad7rzjFxiKUEpsWsAR6VoIYns8Hlz7m
hUnRhhcXHGRyubxTkybAmr8K+OB3NYmJpLLwLCBkAnMgmUZROnjd/jEDQxzeX8v+ZgfpJzZQqznj
znRm+zr/QGxtIJIJViysCvuGvhssIOrYe1kDw1qG9j73Y+AZpAyEv5rYabfLN3FLvzjuiVqX8r6d
CtFytn7cZC/QynButpBXb++RCvxOIcuKgrHs9QBHm86Fp/xGKv7E0wxnHAPYlGK3GnGiTyTwkM1t
f7q5mF9SQtmPUlkCeOsD5nl2tUa8+MSIri/0MBguv6tCik9pW4p6/+o6zbUql1Dh2UOdyOzYcV9A
xn61+94oY6BxLQrMNDfsB1LwhAWorf/XafqaRYTfBzH7Ugvaa135mwmUSYNkwr/lsrxby85yDJXS
qx0/lakZzOOXx8e8sw4biY7h6dyzcwxtQM8HR1jKksUR/4YsUP3TwAgSak7uBXMn/hh0HPhEVxRp
pb5aXIuEPqgQMejkCpLb8rwG9+F2iwtHHxyeFzs8SHySVcoXs4gTTaRx4F8KH9Hrr/iRaegjgI7A
wYycwRWFvOJROUmjHAkSqIazTbarGWAISYzUIncYkhokk58f7CrDDtnXgPbRMxOMSVitqtc1X04f
VhgkMU3DbxEFTk6vJLsvRQzwKPyXEzmpr5zsUqJiKoaC6Gf+3T0FgWC2KjeZ50Kxh4E8JNgZLdkv
Z1VDDzh5of3TZ58hP7+AzZ9C5AhjJPWQfwhsFfXvmdNR8GzAEt56XSGbU7lzgCGiz3styIeCYYdG
tZj4/4WDN82r3QID0k1hQ+ThGl5Y0QhSyxHEsmo/Osp4NX7y7FvR3QIhPjJFmLDL0qccMMIjuan9
Ol8PwKdaoExfPwGhFAnpM/jwiNEdUrCjEYNhx1nQNjaZay8hFwhzqNkRcGmnKbfAAz1mmDDCAXG4
UucftsGzbWCXiKMm3vyBYfrZ8MEGACTT3EWqHUZiKdO80JV+FyH11Jvn2hb+cc5+qUqjvJYmjdtS
cEkVG8WbeCEGtOnOZF0GK1wOY8Uh60uQr7t0h4WUceMmHmZ63TNbqvWLdZIQ9fmF/tKKIBQ+6k+o
7B+dUcCBtqANSQYRzcKaziiPMF8Huv4WTSP8vHEuvr+Ghgb+B722i5Q0jGIN0MbJ4ZKRnsvc9/Xj
pbi7OKzvtzv8HYxFdqndMQWFakp292aGdCf+jM8kn2O27yYmcjKYfhjOImbi9MXfwvESPg195WXb
P3aDJ9qKr+nRxqho/E+pFrAV8NTq4eoNSt0pls6i4MhOQ89iNWXvFs2c5kRzP6qddsfkosx42EOo
O3XkQ1RXwQWIxKKBsM0aaoVnMW6r+MRHSFSlfMzO8B68/7oVz5dalk1m07XEf0g1SE80ROOXUAQO
GtGMu7fNHiZy2mRWbK+rlFArI3wS1CcLwA2nm2dBQ7QaT1QOXNyF/3EY2H26jTdKTNP2yCoNybD3
zj/SqnBoy/4vJQsIH0+bPyLHdavffaG2lzBaQ/IDSFEYzAabV13N08mH+0K0DTABg44UawAqg7M1
SYpaPF0yBP8TDKr7VK4p11LGABR7xv450u7bWy0nbMEetJbXXpgGv+oQ658Xiy7j6P0WEEWrzFBN
G7h+StJeykY5JoPRbXHmGN4UgovA6rvzY8SYOBrsHjxdEmN7T8Oap/tUZfJY+h/sqhXRNqvva6hy
APw7bVFTGihXj2b73ydv/Gj3D7MZN4G/P8SZ/KwaiZFlSNwZhb1EsjflsoOH2kPM9K81GC+ZwYNO
yiBvKvESVp8iqeIy82Kge3GxcbicpY3/Sxyp0db0AWVqU7l/JXv2vFlkP44JYS3zp6HGCnboT/zN
sPMdDjCp0EW38QGoS4vTeQv9tRJgJVLkNA8gc46aLWZcuGgiY4oZBPYzHVopgiSa1N88YQhCf7Vz
S4eFxHR3y5wovm4iJrxKOPwFsymb6UEYJAfOJpn+zumZ9rezC65w/rsX1cyIqACO3p0CA0e3j2yo
1QU2Ki9kWHfY4OgAwSRUxSYT5P1nbnkbc+MKZIdRPMUZJheCtC4Xs7rrxOFAh+D3Elv/a8haVvUP
wje4ZXeOxoYEZ8dZSHP6z/bXu/mg/CDJG7XSq+GvdQvd4hoaTkjJJL4pLuRZwSOsPtdURxzjBJyq
RSxsjnQ07NJC32GLUvMFRM7WaRkpNP0fE95Petyj70wAOKnL9ANh96d9K82tv1ugmzWGxaSkNq2U
06ACP4B1QPstnH5bofVwnEJFGqPM6y6wseglCINtRd+f0t3cQIGm8jOY3sPVqXCMr3np4+IVjSSN
lPSRKjI9AxdmOuEWicvqzwpOMDBcN+HcOVQDb1wvE64iTfQ9P78ET3d11CsHexo5LxbjhSJt/kV7
s2I/WawhZqngsAbVnm2+MbmR4yFJ7BN24/5jTR88w7JqYc/aRf1txQcYiWlf70BRy9tHztuncs5L
yzcYD8UYsxTC0ptEHIMP/D2cJ9Gh8R052UP/PAeq25weWKQJ+PqzRJAy57rhtWQOJqwwW0Y96n/F
iNJEQ6Z5yPV8gewQIxQvR31/11l7VWx8NaZUGwO7OOJ0f179D0hGpPPlmnWsfuUFzouHXVDecNXN
zbz66OQFfQ9JDc+vLltoBdS60hIRrjhVc6W6PbhVoyJceTQUzh8BC3dT791NaNPu920ydX5TC+3G
PxYySF6pqqkunMIkn+iXcocFMm0p0BGBnuQ6wwqSRluolqIvqjcNx3vx2GZ45u72y46eAw4yP+PZ
+GybNRTHJtxQqqkVm+P57GSaIXdivztZPHU15UeKjHYF54KcmURlSicXppHI0lbIuPlgFW/YN4DQ
vhlhh6RRPEKTvJkSYFl3CYafhygKmu+VsdRG/uChH5udKiaCo5jdepcISW3PlXx2qFKkN6jvsgOj
wNcPYFgNFNUPHX0jIYIfLkJKMPt/drwRu2ASpc62C7eGaIGPbUzsuHUl/VSzI32oX6sPbzaCCAbO
esiFc3Zjmurz+T8GmqVyGe0Fm4abJ0xvd0OfbxyeQIifm1yMpddIlOUY+fWiK5CzRcXLJ4Sv9DAZ
hXdvfv0YpPsqYIpPMcaVkVi/SUn0cnxkpFleRuY4+ybziXDiKji/zDuKpzMjctsz+oDWnEtgdSoR
DHBGT8vz8s3g8VS1Gh/DyQadQtxWAWyRFG6flD/ZBm+MkK2R+gbN633MSzMbia0Ve9BH52w8OWR7
58Gi8o6ZITyKgQWX7dTeWxz4xTsy7rHI+E1tokbiJ9+H6FnSIeRC+/9yM5i1TNroYx9+j4HUts6p
GPpGv0eH0QDSOeZzWCh0BNUzv1COKs46JgaGdhKR/Cc8/lOW9rqGcttQkzdkf/bxMGZ+gmqZ4Sc8
BNfQ2ue3tonrJ0uxXjqrRL7onMAC/SWw21UU8otkSdd2rB60qOYwYme4pp8F15RyF37tjK9EdgIa
cAgbYEy1D7ncsH77GTELvgfq5O9Z/+lhUTuMAPqz85ZHWXjvU4I4v8dNLkv+DYN+madmq8uhg1Zs
o2tOosTSX8fzd+ZCbPrMM5Smay/f106FFKev6J+cfceHXYQvDVNqBcEU+ovg6jovw+gYK5sZyr4s
VxtxMsWsTYvs6Fe1R+YGIOO6ngQ6+fcNNKuCRs3QS7OXIEaVOysCjSkT3VoAsKKkvGrQSLRAwrlN
Jw3KEL9r0mbC48s2QuejCdzQmSblGD/6ElX+zaPY4/AG5RKFLz6RSzCEPx6g78g4JlOiEf1HpxBm
hczKz4urjH1QQmIvikxcxNI7Cy6WdaNFaRZW6eStw5YUJgJB6jrhnpP9KCEdwJA8Da+L/rFMxF3M
/qwCPKzEGS2aAv1l28MhM8DOFKTckybnWr6xyv5VkfQ1htH39n9KNz3XTW3ewiHwC66iUDX7WrUn
ktjCmY0cdpIZd6bWbcnhFLK16RshlxrxBoYUVXO5mDmsKicjm6NaPqcOzPtqM2WsEi9mcRJ1d+18
4sW5u6IEgoZ2/deFP+UrEzY0UrPTZ4+bwCIP2EMSRTqXeHTe7IgzAXmqKn1ueqGJwPIFLzY6Kj+E
qb9woYd0yYClERpjGQb5zTaETY2+CXJwBwJNtgn556v8GE0raNw/bZo3KA0tR2fUccs4CFu48hCS
Fr8DgrfBa65/D9iN3lrBH4mZob8xsSLEfI7sJG7AbIlzQYTTmKBOcMZVhWBwWrwvr3AT8yt8qx7a
cy6tbt0HWQxbmP8VDYxeGQAWubG4aPw+/7YdteInCkAcA6XGzZISW49ZNa0HMYwXCAOrEFqekIo0
D00tW/+Br8zQfBX2lGiFJwTvKct5CEEUmqtElpi4QAZKggCbGOX4bO+8S34cNn0xSwf9cFgG5Swr
MHVr2lJB4dFWRaXNyfzmfVJSUrGzWwkACj7IPNzs0Jnoiwb9e9LClVZbUYW1CGi7KHrfaTvmwvMH
iq6RUlcWEIqW6P4zl6PV47Jxb4R2Dniq6x4HH2+ptQKvQOgbHY34Pk9h7zLgpZjb7GwCsoEY74Et
WAz+qyyWAg+tXKrGrP/Kwwqv6+/69P1cZK4iKVtSBDrqenA+C7O972qcQjTh58a+4o5E9IzTT8FU
apMnDoFWpmHhNMdT/YwZKIU6cHYODhJ+E/i2a58v2c1KqAqVWjeg/CdOwy+p4g3PEmupJTuUpc9Q
YBLu4m3XF+Gyv5ESGsGf8NhGs237Rsz4prB/7mss6TalPUwcYRXLrAMB3QJwr0IZvZa8xYSjLiUL
/MWv4pKsHtnb33mL6XfIFnkHy8yod5FmAf/E40JykOIy3sCBTDfUsk84tye86emhhHVv4K0pLyw3
yk++dozYkRfCb+FEyJWGUSmHumknT33z+x/qJuMQCpXHW/cbTZQBcRIVrnnZaFy/cW3Qjp9RvR2A
Ej41xhi3LODlRzTGgH0m9filEVf9tf6eBs3fD2kya3hd/qbPSPv+OyhsDPLYFUtjhjRP9/MbFtN8
rP4f02II9DlDLOYTOwx6NSKN9iXskC6Zz5T0Ev7OMiiryCoha6sqj/3YByFurOdCMtcHst4kuBGe
vFukTqPt3JkFU9Ccq4fCFv9iLP0rEzyc9M8rE2c+68V+vj4Ho9rTmFe+VN938dl4Hk5YuWPZ2U3S
PHmhEyhtn6oQE/yywhF5AuEIsAhzVGDUs74tQf43FBA9qXkhWxkWmdxH4oE0OW/SvzLIJFLSADPW
x1ggrsMSukXovfybpp+ekWBsUOdVqlqHj4Noiatyhr+RBc/YTkad3QHrBFUdH8zUzi+6TIAvPg+d
hkQQWPouVxOhqhIV0d1n1flkQQJIryOj3x+xu4SFi9wkPh2CDiXRh76KqkfUhE53aassUxMKXtJ9
hTGt6IAmN3xlfCxJH4g/TE3+fgkBBGcj3qiZvOScTiybIkR377OAdW2OI9pbWrtjlIn5+3lDLyh4
AKUDWvR+OFbSEKx1RIrYIb/Z38FETOuVkqDO5vvayDTgRNvFiLXnA1faSLyNxNRpCZPTcPkNanDx
ChNUAF4y/g+N/3CSNQz+BBe2oVknGrMxxNMwV0djgXHUlhBWDQKe9z7TRx3RJ90jwqsYDeye525A
784XaOZblTvbcNHLuMYlmiWfDXFCVBuzwcmhrKxF5VQJerL4F8WNVVR6y7rZZsqIu/45UNSUwXhI
9WmeqZ7bAASFIVx2TONcD1JEVXeeUSHZxfGFs9STeqPLXE1Hjdsf4RPugA8r4H88VNbg2nUVXc2+
v99f911YV1suujClaj/7Hb2eoRiEk7VgVOJUjCek91AlbmiYWrdX9/zdLUh5Yy/W/zg2jFIpM2Qq
chT4rRa5nljGGqHX4vCzA9NRN3DKd5RqXJRLMDggPZ6WcafoXaykv1/F7UbeD8Cvf+2jvZTO1f7Z
0eQ0hILcTTF+3XINFWhuUqzUQJoFKwUvBqHxVBD9oOX7ogJFERJCP6r2ZKJ8JLuotHpay2Z1L3MM
O94UPBf1xQO5A00WAHTQguVMdXGiWUQHNpVVAI9ZCDVkJrhnJrFGyOx3AA6KaEFxNt/aktV8oKtb
0WlUVl73uB7SiEC9F1rAVNEhefMYjgKtmfRbvCuYfWCxx1CMMNy04HMCq+LInA6lAwKZOmM2Px0w
i2ALwyKqCJqkLZrNof8wxY0CpGdbBkS8mkEfajNL8gbO+VwvJ/kigaROaPaKpZt/i20ryM+j1cZ9
Q3WiwcUaXBm38OOvrCdYzGALuCl8STeS5ti87dqVfSFiHyNgbry35svkC24yp5QbXpTo/usPtryz
FactqoDgkGyEnpEOyAV0ts7XcqLMW32iinBzya7/qJgqwKsfeYDWnK9/Aa3KLfhURyRYT7f3TF21
uIxqsFqJbMEyK/GSS1nkp5JqP4SZYemDqa3GEQOJvQuXLA25Z83/BHhZhmOuGgta87IFwVIR+CHy
qrtl5u46phybg+hZmtVRTnufYBgpj1Dwb6v7Jn0nfU1Skqba9OsBxPE6lcRyw+p/eKUELzzv7mPd
yqaGDRN626cxS0vd91PgO4ruBTt2La/3UyZwP49zhtNK7gML80k0yGHHjAD+MO9aFI3bxYHI3zw3
zk9ZSmDQWYlipJEYRYIVgj7OFRHKkxHyBheYKu5QCV3Ng8f8TrKdGRYO+v0+4J46dmwVJsmaUe9A
wGCVFcmHvZefCR52UwIPMWLvF7BrVzbF9TNfU8EsS+H80jorP97QWcttWimhugKzYAbciGrqmuuO
jtLZiUijAA/LfW7ajeanRHRqiZ24oJIPF80qHAbXHu2eeai6QauCtu1csZG0HsW2B5pG92J4fIbT
q/ltf9UqxTHT3cX0El8CZm0Kgh3nDlHQnc6L1PO7bz3We0bWOtbwtYhGvuUPLLvvfSlg3n9CUFrU
1nzbR6WkdPXA7Y6HRRk24AFpE8TA/AmUm5+LSwufQaGRrkL/y+QqhOGvljnsh9TDhmHVuvomThe3
Nu+RZHRNsAbk41clSqROLWDEaY3Pd2vbSlrg0mT0T39lKXCOW/qbw8MeiJRrcDPMekqZkakfGlyi
shXpsWZmbMQ3L+McyehqFxw0KrXedghcXpxOcxgsdTgqJBQHV8TmJ1FpjCT/5m2401EI2jDbZ5Zm
RrRKlkB5UjEtJLVCfHrnC2/l2ocfU1PJekciy5yQFPycyRoTx1GNacGIaYY1kO4M/hG4oOeul40m
L/ntToiKY883TajiQwZVpMsuddpJ1Pkrx50IHhvmOWiGrb7JYKgCOlQYa+BCkQPwqs4OU2SxU/i7
3VrzhO5bhr9QCnYLjgHr9j9+LouhnGqXUNJ+DCHj6tONxBBHKWKNYhFjIWv9pb75UdxCR4WrthDl
bJh//7tC9GMRTNtrzARJ6osbl8rNAHpTv60GPrt6mZscMNgbLOqyPJy5Nf9yt8zokahfOC+Y8SZP
DwbJ2L1wQ8W0RsHspXO3msVgmx4mJ+dIHtjMOdS7tqwmKx4jMFueH4aDCauWrEbnPX3Db1WqPcEh
J55fQHXHtH0rEW/gd6J+sDRhdppnue/8Aa8fRxX7pgAzomeWa6Ic6Wqq5DU4LjIhfOgWfE38hpDB
5tW9iVxSugjkmvCbI7Qjc/VmN9+r5T+QIJa3qiGehV+tsCTtjbEQvqD65riQULiNRuLDG/b3ysoi
v3iLPkcXNV3Tl7IF5QqEVb5/pealvthBb3+Q7ihJAvRUf3aKwR8HADXZgXngREpZXlg9HCOKyGdA
sVZE07HQUMy1gvbdwxU4fD6vFAHbUmHrMG1E+IBS0QuOBzP1zObantGi11R1gyyo3xL8/S1emyXZ
UbjNwg1GRRrA8EPr+PtjlrHd4TuLSKNJMuW5ALu6Y+EwqQEcLHpwCFgT7HzGB6tvPioFm1cnq0kI
P54gUUsr24uIhzgFlVXNWuM4ozz37nkKZIT7nUKEQlH9y+RQAJ9qAKx3vQ8C/y4XYVHuJs5MFgV6
t9aUBqAEDtm3Ifm3A/PcWQ6ORODtUBsSXHUD+n5lsjivF9s6Osvx2rk63Es/4tU3bqHMOiS1vHCG
Sujam7UgFC4QVmCslxwBdl5QaqUXz9/MYOgEmJ/ph2DKyjdEIClRz4qEN4MEeJu9Ew7f8ZOgDaUf
vFVlOd5d+gMZlhROE4BKLdmKI9PvAB88JgX/yKd097oAz/Z0Red7K1m4LevpVxDvSqVxBwlgkORG
2FDTFnc3J1HN2jOiW/eWS+e/wqU9/2kSEaHaqYpzOVbGoJgxmlSwrX2sfrfKLpysiLyrxJB0I+y/
GhXARRX3TESjYKQdZYMkNXj59x2O7HPP3m23wcImnPILYDVq10cwDVbyA7eg4wzuL2b7maccoEhl
8gqLd4juhCvnng932T43aoy4Z39iGsUsC1ghgl4yyrjQ94k57dLKBPNTNQ8+X+Mx/8MtDj/T4Ose
5xAcLQex/BNJeLWomNam09tCAiOGOseOmXTlfmOXLtPqc7YV1FOBBrrsTwyCaJxanL13LQm4Q+mz
oVPhHQmziFc4P/3tT5LNuY4fJk0kjWP8dLMLTqmHa4XjElqUABGz/b9vhFbCT2yD9nreO88Wc8C4
qc5EEz8ADniEjdFNFZ8yS3T7gr3/ZkcztbxRKavkQEKJsKtF2exP7cY3TrFbMoUd/BTiv9sPeyQ3
6BUOE7/+TeTAP2StthMivOOEDwWZEqzrW/nKnp359Rz9eMn4Q/tzaer5wdWCWIwYdCsAveGyKDvf
C2TvCIMkIi6qPxl2W0JLSTe2/QQ0vn/LXAYvJI9FqhvP/1gv4H0lpDB4roVDtAbV+OFZEBxgMXIk
yNYTtTb8sFA82Ls4rSQ0YCuQ4BdUq4l5D6QlLJfsXfPzcPanteu8L2hBCVqM6vqwPteqW+BpfQCr
nyh8Ufw60DFrrn4krVEXl5irkKvfrSe5p4krp2Wb9bhb3GqX/sqvZu4u2vJf8qgA1TDDdi6KQcwW
MwZziZEthoQED3RxPfRikTsUSSnOUWfHwoGLYE/EmTooisWquzfONeUVgajToUcy6UWPCG1pf0/t
yEdV76O5A9Pilr8XF3FG6AhS34IxbNM+KAvP9g22M53FSPzvnEI0Zuo8UAFRqu1ibrhwBen3MOWF
4tjr5x9OQ5PuAQX3yRjSEx04Ql4BdtNqTZZDtLTrFMdfVQMWHfcGMZaMAsoMTZ21psNQ8ozoQuCa
jmdvoKo2J8RJgyo+NonbvcbRLooKM/Vvq9oqdo2lHmuZO4ZS9SnTmjsy8jAlsHcYUdVrqTfHnZIs
vCLJZZi1ujhDPWgYp1q3Ti4NSoBwGQWhPBamIEb850WmKZZ/HkEc6zGwwl+qplkbmn9cyUYW7vpT
R+AsGZ4tdb4NFmKrV2f+0JueLSTER9ht8oKNXTtJ6e6pKzcroXkb+JBS0m3QEA57Ab0xEM0ynD4f
l6XVQfQ+jMC+fMURzyvBO8hOwojUuXJ3l7CZpSS49ksQtRg07nTZkvG9P1R+eN5gu1AQhYkNxYMG
hD6+J31LNs+KOSlG3ViLuzliY6VYAcjZDy6Ha0sU3qiQUd5nJLBz/MKKbUbIrDw/AzFnsakMszwH
yPTryduhqmX1IHrEQR1ufHj4j7IeNeDC3dBOXkBNbqc4reRo8p6T4S1L8gCurocfXH5KNtTOJrIL
JiUN9WW/8TpOB+ObIUCkM8NYI4nQuQWvBFx6Vo+HBsiyoPgaCuPqNT/NsjO+5CyPZ5irKNfdrVhw
u46G43HSLhGysYa18hmIJyz0veyzuvH/YrjvOn+CzpBwn0e+f3rYJqSfvy3lNy7mrJJ8vXLwBN0O
IOOz2Q+goi/3eVOmhTGyGaN6SGqm1HRecQYR4XwFxduysGCyCKdABwV62NATEzIFxXlKJ6MR5DIM
ONIftIkbsDPg9NPbFcWJJIOgJ/LLnxCNSOutKsUVffRDoSqU8Yy1hX2p5PkBemiilxEErDp6U5Wo
sAQ3IIUfuGtIW9T+7mk0VAiBCWRoG2TaADWrzGesoGusNU5ojmRXEpbkeQEubR27Jw5oCqiHMLAN
B6cue0yjGjZMgZV/1GiInNH/AQOlOSR3Vt6GPcseuDyYcb3b6v+JdDS0BdjzWfSQaGj0eGAfYpOk
UVVEMIe6BYSgkmjH2r5bqWPnVynpr/S80YSCul5hHDc91EinlWjLLWyAI2zvHWvSmXT42ozgDmrj
AnkQFMBupJACNwA8LGDBX7a38LW6omN+3S3V8gOBgJW+SULfLRthqRUf1zsOIIqxwWaCN3OA/H4s
1+xn8eTrl6N1ozjuLWml4NOPK9MCoLThahv2fFR2oOh+qyQ1xpji0nl13famRf1I8AxkCnD4Rd9e
UJ/a2HG2V75K6Xs73fPeAqMlKw/ZWyttrS+wXIKFXADPfxuoiaAKmZ45WxoqDrUeW0I1V15HubV3
uvbB3jy1osiw1Idu4d+eJWEpBAFQ7CnDyooP5kg9eeX3qbRqICr3v2GgtmXCH2K9vhKZqKCSOT4u
YvSAlAmAKacaE6a3ureOzPAzN/nl2U9WG+7HxIg7glP6RpipAjRWOZvZvnhxt61SDY9OyVBfaRbb
bHR8PFNfXGQdC/ca/K1yfCvZmwLFaH8jCBGrlV141NjQiL714gPn5e+a4C2Ujc+A8y7JnroE0rtF
abjiDpDLQQCJNS53gC98dr10OPggbSbPbsT2r2X77wbT/dVNwKmm0Iuoie6kbbLqJsIQ3ZfO5x2Y
ioFD57OaaaZ9XmCTgrxzYzyfB1tIeMtk8h/ew3XzKwzURPMpb977IwKOdTmiE6iSIlxn+GSd0Sh6
U6ZnBI4CAm2C4LPw12jLmxLQjAXm6PtBnzlDbsa3Nd0QwPQKSsutrigocmOXh9yXyIc4Q7UCSrsm
B/NyURM0Rlzx40VgRw3/JXOpKIw4XVZg7XPyX3z67GYywT4i27UgrqAXpxrSINbzEKZUjamBOe7k
/85OO5rVLiVUBKPgYw27xCh6IFJ/mZfbNo7TGUoYBLwbi3dfPqJiIxyeaEodith1i92sadedDrnk
fxMZiSOR4lKRh5ofcpHXruodl9hj8jRKHLSGdAxvYRC2sQiUHYkjJ/p259UKPWyUln+KfJB2ufti
u0rDRKGd5l9xE0c4m2bIud1iwPebg1OLo2wkcXqgJ11KkSeK4j/ff9o8PrHT1Oc/Qet2IZxgZXA6
X3atWM+jS9L/EAVIWpS6WVCepvbqkPayBPGBICgEz241EzYKFE6H2OEyd7mSj0iQEmqCpMBmaz0K
WkRqN5s3fbYagG0ySrKGWTCUklDVTJ5ZoAPjDdAKXyj4JDB/j6F+fzxYckN6VqVghs6mKp60tpOo
5PNv3SZftP587loZtEPmfLLV7PTuZke3Jnt7gBBaaSudyedVIwhaWlkU3CeCpfeJ9htLRoC+ucWR
4NSsTJJlFNapQrWqXUvyLsZRKfgmjobg19VlTsstZu3RwfFlAZIXlkphmSWPHSTwonTq4IlwR2v+
NhBGEhwum+mDp4CwSTv+zJm3zlIS8WvOw9ZFUJS5yzfpgsOLAUDZh8VUXk7xEWS3CxV+KG7aFh7K
Qx030kisilkocRwlVyrrtyeitnT1BQuLSs3b/O6QkKsJ3mAFKvGWQXEdT2COmpr58unVNnKymoKe
B1sfq0ejhx1spO5F62QMmF7uc8bmlw4OhSWqZujsTLk1gY9Dkw21J9RmyuhEKP6X9gWd/lpx17LL
8v9XiqjUl7t/+Z7dQ/Ph+nzgms08DC+LByGm3IqqFcrk1ZXVc/p3LEMAsGdLXeqIPjB5HNRDqA9v
PlPk4fzQx2m3ZJhA2aecIqqfcpVZcuiaSJF9aK3DA5o5SFGBqzT6E5sVFxfX1UU6tQpgNbnRZc1E
+6eujJ+47Oe3SHUB8NDR81aLdFU0aS6rGZtXYNv1bd2jNibyVeUUlZjzSMGPGJ7WkzoANDg2mDFp
9mwMM58moockdpDILEu9cnYwgDzbAu941ChEWdXAA9Ip9IYh8aw6bWsfdAB+V3XV7BwHdBBE58Wn
/ldlT/L2AzvubVTreWzKO2xi3b7OczX53m+GJFwe+7xyZHjF2SpFa2x3chzXiN4ZSBMgyVMzOH9Y
1OJ/euP2XoJjR0vOUX7IglCnJcm+6P4pfgXwV/ghgpFlE5yc6E5fJ57dHxpo8Ex8umgbkWxcoBcQ
D/WR0gXnGsrhlFlzg2NtAiwFFrSvAFfBSWtb5QLXFLy3hFEt9/t2gxOujPYS1tMT+wxM7A1rPi15
8tWugHGIEm4NGeCARiK3pOof1XLcL5jlbL6gWXnvqHTyhkqsNnPSx/OfR9i9i38rTEfJCrhMdun7
/zrNbNKCIcIjuAvrzLNt3cDQvW7sfUErNv4V6UZ4Zw1onVjiZ2DIGZsGYDMf3p/SD0vcEqqDAzoW
RQ2nLL5Bqs8bt8Tblh0loydXbWcFPVY3yaZRk+a8RZpo+EdKD5D0bkCViR9pyKsIF9IMrsr6FhuX
v868EVg9TZ3zxLYGhhN4LMS/O9LUYOcHXE6fCKFeA1MX7T1ZytorJrntIDfDOrykPP1LCxlkVhtV
PxmKVmIsYkhD5Ua9czL6pum4E+5uwJygl+FUfvOqk2wefvwOUzIr6bXtkdtSK5TyI1iH+1NExiO+
p0MSjK81yxDenzk6DMMABvsUqLzKh2nHht6s3ZfYgzoCUovxzbx8O/obKvSeyNDAOb7srn1prW92
h47BzibP8hdOMwk50amRTEOeN73jlCXYvsYamnW6LkeEjenxbln/pGOHX0Qwtq78ZCTAN9cBxj5E
1o1ewMAn1BvybiewSO5XG3oJzZ5YoH/+Hm6fHUBn3Zl0K1Caj6kyMO6A5pXoDFMOHMynyUOYZiJg
aocCT84xUKRfdQdDF15A/L13aXzCbZSjPaMuOJdV3nDbZpTmG0+yIqGobhmF1P+/kAWHGWBNx+YG
/ohw6qgh128ZM2NHo4g/Hnfv/r+W5ns2qyzqft0IE17d8Bs43YgAOWw49b9wzxYG1Tj1Wz+PRvsP
QR762lUSEyUvbw75iuTsVkR8SrwbbIb10IjW3JhBguyMUI5hwpDQpqeGmjlGa6PAeP3RByZewWsV
XwJPbHTaHEfpMTZ8ipQ27YV2kDJ8rBxKichZ3n9p4ZOFfLX32c8y3ImgmxYCuWd+xeWfzuf0jjqS
MUv5JhqRGAD0ugaa4wBQcg1ML6HJSPzcjRQo39gW774ULtx1rgpCSQG3Xl8ZMDkXyxHZJN3ykg93
y1EGTykzJBvBpdSDTIbCiKdCkxJgo7fAvgGngbtkHe1SOvsH2czytF+zZ5hXtjI4MMeou9CSI72x
vIzQ6b1jxlhz41YOtQR4qygOqBV+WnxolybND1GDfnpanVOrM/1vnD1N7Wcfo2HlJ8YrkosGWfSb
eYxOXg7VBZ92prBNVCsMMu48Qojqu1yEU7llSSSg1/Moz2lPfkKxD5T7EVd0LHOaPkZDOEvEyG9R
sUtUdWJCmkWdmkiUstWLPqir+psonvdsLaCfV163fyTAKxoSHglLKCnXW2oho7nBA68X2whhYubN
7GVwi/mMeyknH+AkB2VTiq5/+jyRI/3rh5Egi2HClO6Yvss1VXK4oFW6xDv/MRvThQu6SeyVV6Me
SVrQZi+mwBIJeboZo3dC3TZbGSYoDF4lD60g42N1wagar09wUsvsxXY8BdNtP4XmVWGtTtwVh9no
fHP3HRUCpUGwwPzyJC2aF4qewcKuTLuC+l8UUG2t1dysBXP03bvz46muXFVewEi5LZku8boLfag1
PveL104b3agE6Ln9TkUUJMXsZOEgQLGYv7k6Nlgz5bvavz5OaZoEewiips3bvhO3+X1BgKGwfgjW
a0aSTi3Z545qcy899B1nVVcQ88HAs5sIRyJSMr+kQcDG74b3izudbHgj/L3ScuRKEgQPApBRwA1z
Luvz9+fX6Ow3XxzGZZOnJDJzlno3DL+whympEvNJLTVlj3o95jPcyR/YCdD+PIHhrpCs7gkwe0+8
uTpEXLS8+8XXLIC5F23MaowactswHbOnycurHs9rGs/V/Jw/w8c0de90PEhRDhdZQ8OqoI4Jw5TW
Tq2UPFK0p19ItRtdJXQgIEffsA3JIeEbRQfWZSJb8eFZmHDL2kw+BUuIp2/XwpIoKGZCfp/7DujZ
lqvH6nYriKeXtaWpkB2AC720XIraEq2C71iuBTi8PbIABgat7En99hG4cVYdZZZ0Peo38ahL3ugC
/qSxqF0Es0RtXGLmynmCEbWGKE3I0yD6jQPP0ne0Tf19Tt9UvTNd1f+U6EfxD3gSPEOD/k7pKvuI
4qa2IaIxs7pWlUgzKiNt0lXLdizcdRYgNKtbPKPA+zg9xb1HBuo0457Avgz/SwQrTtYzvTGa3+7O
zYSQ8NX3RfepX07qo3QFIcPDb/X/OAmQRgPNTQSD3Vm0JOZxLzkLj4OCYghkCYKZIwzB586GbSFa
+6AMZ9v0f3+1hUCeM2/Lsd12Lq/lR6JyhoQvWfIhjJ1kqLGWF4WXMVEU7LLF9K9rMy2eKIBPH+lL
mcysjOktF5OupD96mGEw3/7QTrHtHa+4yZJxlr6w9rNBhQrnVIf3TxENrJHs7jFsCph4ImT0DkTA
6v/a3kfu9SNOe8JuV2xfWTfZJlH0If706pY7bQHoq7eBxtR8GdZsmy/W2/Oa8S6W2vAEjJdysAnG
SisiKYCQwG3n5I0chOVn55ShJ9l+dgDC7pA8k9xixsICJAjJfIuliZrED7iiVGZGL05hKGLF3vb6
YqKMvO3t4yG5eU93BZZy4Un1WRfACjIHaOTN8cBfaUHUUDxhIs4ukMU3E3f0Yz+2FVCaD7bhKteB
fpS/JaO3bYkhEEySh4SlxyekN5D26Gw9Gg2whpRI1jo52zx68OfdED7G0/OuTFd4kubBYsYVyLGt
1B7CFNQvPCZv5UwmvwcdkbQ2u2ScHOrtRLZtSmlVCBxw6wyFturV1KUjj2j8Yp1+SjbT0JApuCKb
V9feMTb+RqRiL4OSCF84rYJcMjri5DBi6w+nE4Mb9FmS0fCPhqNzH13TPJSdDSS6goKvq9pqY526
SiB0QEV54JRSCH1Fbg6AqZL+7wNSq078bz+nMxFBenw8034vR8MH8klf7esEtrTA/Nz41hpesJAR
51O13kYTEEPVGhhX4PCWQPdKKfkHxZwK9/2uADWwMmnj6bvVtGw/bcJogZtBw7jHIJKQuxRYYDHp
+uvCb6pvOVTUJgjT0grdUV+uLfu7no1KMWYepi93hAqF7D6g7JguvZFO9KnBV73068B0raC8fu6T
0yNkwjPuceW+hAXPr+KVPWlxKtiQmcVQYiYdwDxBTKYB5jak4WEb7qT33ubvXRw4qVte8mjYIM9k
z2hmXy2eYDMq/wOE0QALGdl+qAXIci5VWdGTL2boBbkJr+PgPaNtal6nZM0g1i5ggsxYy0UZYIAH
J6KPn7WxoaORgWC6UQUGwPyYR6gWYk7srlI8X76YNdYUVHOnGzE530Co1jIHAYqFt2TAP/p5/c+y
f4gG+Q6WRu0gvvDrLzTUVzaAurlrGYgK4grhOn0tg3NibStpXfxQT4gbdM5G3wctUn9GOlkG4o1W
bOfA7iWLsm2rPWYxsHsVJNKxhb8DlpeX4ltE2fdiSBPCks+Do+nhsKj8CTeRvjOEPpJcZrRh96Mc
Xeo1T1g6ZC+iPHzLIX6IiZ0nRSwP1d4AfFSnQv6l8KJdBnmilOK5yD0Ai98Bc7Pt/lyOGO/E8bID
IQSGuTvVtUX2ai6wfGNn+07OC8U/ap5fTSdwseWJvprpaOfYGCqlWHiRDB2iGS7q55cG6HI5z/Xi
DOLNJdmk81qala8d2A/schjZRZZH0PDnGPCCPsDEPfXohGu6kuDNWAb+++Kpx5xh4ODE30EAshwM
tm33BuxPlVSxIqn16Kjoxrju8HEouR1xA5C09oWnB7V0JX8ucADtPJ7qif0eDbusxfb04HFFHu2e
D6HlrAwj9EORPouOew2FC0O6UykT59lEeM6L++77mB8LNDt2vmTL/gzv6toGCHoyrC5eFK2mPZpd
QzoQdDfBGlWmRqDec4inxxTU1U8gBp3LvyHHDWtn26RapfiunNVetZuTZTSHFkwwaz5wNRv1ZRQX
S//hnpV/q6LnmuV5LlUfQXH6srJVjci+TGvqsV47jpT1XRkwMCS2NESLt/Z6SBzqg1E0EFGOXXy2
7t1QJbh1d9EFhMsbm7BERJyttt+ali9vIusiPONCdm8LDD0JilnaVfNkNVmEJc9ZOM+TLXG1XvTU
heQt7QKkQnqwbbmeL+sIaIfBobqYuYByN7LBJmSPXhtXhLOZ2ETM89BnXyBS9LzNVW8H2KCZnkss
FfrNcJNe71+D/kgCZzZUwwbckmuGcJaKHNz8zlHo+7KcFOxlZU1ZbGFPBe2DI75TFtGThj+9+3GT
0/DVRAvqB/g3wGUV3pXG8SDobUGfraj3LRRlAN+uLD+rulIQvOlgNMBVXHo6MrLzSR/qfT5E6O2z
3qlH/O2ibsIQMFygqgm9reGB0DwIyiZoEEJfduzMY2PgCrjxoon4yX1HvuDNrJ+W8yjSBOuRnpjJ
2UXyRdHPakLZ2GiLtrBkLMS+5ohVgRKdnZKrvec1izXeEGL4pdVqxdr0EESX7FCSLn+B4faupeOV
doTFncwxj8JWXJM8ceZ+9dzLxxbMZnjju7ruln1qIGZEAbCUcZrnoOAJf82Z7VA5XgAPwS2ow4c7
EakaaNfevI6aFTT1MAyT0OwM2Z7Lw/wk+7eyQ3JReNnWryUtG3ckFTqGAFIQOgx80FIkJ7yOVxzC
3TPYCSL80O2My4F0HcwpHN06UvNzL8nrImBfQuPHKPSKbll1OLzN9gqQkF5iIHkTRvHKza3BpdCm
3D6P87QYmmJ2s1nmzfdRrtBVFZdDAvvbckgcDedAiBbBAkIwRaR80QyThrGyMhWXUoNOyH4QU0lm
GvDYK5FXID3GM2GqVHLFLBPKb8QBuhVAVFN0ZEro0H+shHyuYDfod3aCYpXhZLpc7VIhEAVXNh1M
cJ3JK1u5lzqWf3oh24JRnj6ihEPzfEmHvJWq0rgNNv6HJo0fHoPGkttIWR5ni2odJFtqLPt+fcZW
0pCEFx4A3lZhmwlaEcQ8hAb8lV18BmGDf+WanVe9WqnlG6/F6yUKe+T3RkBrvIQZegdl+JFgKfhd
06ADv0OEn+ETpxzY1t7MbpfH6nZ9bSxcs1mdkmqoKYdCga63l45IH8Q9vTpkSho2dM/HzassUij3
EHJIi/pRh9rIuMafrebhuMu9w33tioFb042zApBjmwbqfUZR1SEYjTSTDASPLKWsQeA+E1vOxRkL
eID+Lu6UGISiMsmhty0sViT5pe+Xx3FxkF4Qhyi8sCt4OMoPpdpV4Pj50BQQx15c+AvzZD/0JXm8
RlD7YtebX0ZQETy1ZRN9IXChmg2z25OVpOfrSyp64EJlstc75DMBEAx0BTzVN8JlbFch1vBGecjr
05qsjvN0QG0sSoLEi55rN1wj9hpHCR3UgvdCsh8QtrcGzprLJV9bqd3ca+iWknlR7JusDTlADIpy
DUbQYQeAOMKnvuAcehsZnOu2haV/kRI6a74t4V8/t+GSvBqAF04fahcptIt+dBlLxI7L7Flkg5od
z8IN3+lugzWLJiEB/0zKKkUEoEndq/K6kdA55htk7zQ/Bi+hiOO0XzuxLGRtODFEfMHO1yGxaKn7
ASOWO0PaSYA7ZwH5E5hYyVOBw3XeBAkax1WCXEkh/sJbQiSlJIIBcNGLjWOpYWdCJG6FXsrakIMW
lVKquYcw0GUJiR0TdjU7H9t37WF/57oYwBplsjzyeMwLYZXoK/RBg+EUeBLUy9XkrQfpFKYIckru
wYLUHkeUC9of671LKohFuzP7FnYNDFqPY2WF8U8kVNrWtgH1debcSYsOAZmKmnJlLicPsm2rZ9+W
Upld6OnEw0crJuypN5LcSzZyfTG/XQBJKcaTWvS44Ry9mNJTwHIYgsWw8N/UA1wz8iRO9T+eC6bt
UDA/EoW1zsiskiJEO2l0QnhLCNDFcFWTQJyGndeAytsqk9o8xwp77b/VwSR9uOM5TUjkpa5ivDtA
lD/rUbl7tpq6uiSvEqLAYJ0tksouQe880hG1puC0DpyR09esMpRp+mLhOPKZwY7t1AcU2SqvtHgG
uj0lnLebkCJmbm9tqsgwk0jGn/MaagbL31ff+59ZnmZc+T//JS+DCe4WECVrk5dujR2IVGmH8irZ
2pPub82elmgmMdE043BgHiWX//nUGxXy/pRkCU00BgWKGgkJZLPBOecseZD0FVr9Nah/9kUla/lI
8qxSme+fcE6Mg/Wpxl2Xr4J/M9If9M0KEwA2U/b2nq+G5JX3mo9Co1/vCnWJywGJAqs0vComjzoS
jRf3Pvrhg328+lyIexcLE73ds0lcI6AQ8sjF6aRPhNTplLBK3um0zh55KmqokW3BIpPizfVbONEp
Nt9mnDVeigTvPkS+Bi2lFYJ6vzUoqUUgbUB03GL8qP42lbbTaeGO4nDCh3hrqlfZApNB1EQKRr3X
de4D4/2ov3ktm6HBcvY3WfRjeR+zyAnT8ykh0raPyGg8wYcZVuzUoBPV6LYaLx/ruhPeW0M6qqe0
QQemTEl7D48TxOzzVo2JKdMaOGhgVfIhiYeQvAOp8ro7AyrPin1BwWiuUaBujwuit51d1Sz7nwyN
4d9sfyf1Rvd7Vm+OFMUezKzOTyXAl6RDeVeB3LzNfSzZ9OQaYorIyDL7zMoEUeKVGi5sljG2fWKc
nOS9ibWcrXcytHbdSypvIn/Pjrg2F3t/KoZLuyvEO5+ds5aVya9VPTOrrQ3lnOhDFZ3ci4ybjoai
h+O2QDW8STSP+evbUJfpawgKX3QmTUzq+5ICbM56W3D+a1DBGgUyg+eZxTCgBNI+MCZCIaJ4KfSO
RqPUwOBSIau7fShoAYUQ66jpfg813PYVmr/dQuxpiBZuGBzOqmAVtjfkdOBZk6ptsUBtb+Lkd5SI
SxPQdR3Gx1/cmm+LNtRPUOFMPHaGGvqS/poTmoPiaHKlXDdo6IzJv1BjyFp6MkDcePSyXkiXMltO
9i1yUeQvIusHso73jI+tXVXzScZ62bHWTD8Vko/4pOioDjhrCbHjX289wwY7IN/b41LRRKqbU8V6
smRcPlPVYAciltNEupngtIyOWtVYjbb8H1zmNqEgY58OOvDQGUIASWCQoa9g5xdeiSm0vyHLQMyx
DDAHVQfuhpFdgmDd8g2SXXaGUKjpXcp97gsA+0UH5XYOExWPX1XoAhVUejhunO1iVHyE///6VRWf
giiEGIswLeTL7r16G9crlxn+rGdZklxWXdi6Or7yAE3Fdt6h5T6szkmtaKaovmbsRHYqFmkHnYcf
e9awm5T1poLGqeiv42lteMtgtRcjQ76IeccWvSQ49bw9FGtPfFbH5fIg8WSCQ6hetCP9nNynyBFs
2Mo4JoaMOw7Ql/msJ06eGzDUV+43ciZocm20MH5PO7hiG2aY4yG2yV6h4QK5lzBj70gYN5S2Lyrp
NJ7ypk24az97vhhgaaLasTV3jgJ/i2SDh3+TX+W8PLoRo5fBusDmIBJzAcuAN3+tbfcVICrH69k3
oBWqrK3fYfQAzKLOgQE6P7vqLuD+n4LklbVAXNDD/+IHM7B9g20TmIKS+A5KveyVWbKfU6RjgsFB
5H/s/GyRqRxG0PPckzPDEeqNNO1dzj/+CqAvo8JpPhnNiT5gHXXCl7v1JCq/ZtoL6V06yyh6/Zko
1aalVlsLugh+93gRfWihCAMNkYLhkNs51QXyMDZLkXPgbd0zrcSI7RL7kKlGanogxmJSiJKrbuik
LGMFaDNmBxlgPe0Yj6Jl4deXQ3Ztd6RZZ3OJuziYELsHvGqHy4Hqog+qFBpbHo6mEz0bqMRsuLiQ
NHLQiHBj3ksRlAiDL1tT21o8NVjMFO9NGp8/utvuq3f8AS1ObRVdsH8Qms3eA/GdUlDEGI3cg1zW
MfXDa/ZaEaAfpwhlzZtt9lSRgZ1WeBNrYoCFmZfxIFVOc9Gl9FuDluwBGf3Ui5BA9Cp5hCf/0cVg
Lw6jPvrNFAUndqQUoztJq7NlLredCqiSd9VJHRcdPXVBX3U2lpGimaUXkR9o1KlDIwJqSXRXdfQH
sm/11lOya2XuQPDXsGHwSersTrC2hmL8ztzNYQ7SwV9iFsqRz4OkizI7iUmIRsBAMEFv3gGC/tGv
OKMbI45GQhs+nw1VKNc2lDqV4EQHyc9xIxYXoB6b6IEGC9vK3/XE8z+zUtAplaoEongZl+w3ybdN
l/D/Yvh8J4Zz4G9Cqdx/F4TdTnb5oBFXKZkVVFJ1a2gxyAt5jGvivxT6Zd+gxOEw3EUgKaOz+OMP
keGdjQoXyxzTIakxIMK41WNlmyTB1yG7P64F1f4AG3lp8ZtThpYeccwYBC7Ip7o+W6bwWpIFKONU
+f72Nxjnk8KhGg15Z5Nv0whSaOfRCkbsJBpirj6ajmKA0JArJ9AVA83IKMJ8ZQRb1Eljll5BDCf0
ccDkkHEVcVG544y18eZz8VdWnlYcRrTfTuJgDwI52YqNh/JwMYrLXcKCAIa7EhSNmAVrclCXS1G5
cdTMwOBYquF51ksgxIxhvfX8xnpUF589FAu0KPTSucEG3LhZaw22TJBBo26b0kiuyMbJc2ZgHX/U
b5JrlKjUU/DSQMybEH31oIxXXFP46vcUSm+2NgaYnxuQqihm0Ua4CGci35Tyf+Yc9sL3kho3HUyK
H/xI2jD9AcAybnzmaJbLCT+NgBkfWvyX+mBCuE64Da68mGZUTX07D2PWkIBj+0lDSx2iQzYxC/pK
raX5P8sDW1xA4OH64MCcpIl8BgpCZL7/1qC86ylCguZy2DRLPsmgh9Bc3gz37TYLmg0zsrF2M2p8
pQG3tNsxIunRz8iuj3/zJ9TUIwLaHUMrB31TpKNRxsH9fKypf8DD8y2tkt/+rEKOgZvN9fUipDGH
oQt8a7Kn2caCCiVd3lYTTRY+8szJBcR122RQcNFmfuJSepsgFwCm03bko9WkOk+9ndFc3r6oSJF6
9XxhJPdyjgViVUek20oRFqTMO3Npc7SSEHSgRVJHuveVDCV4LMhq+81xZogdJVsWt0JOYZBixogf
dXSiYghPm3Xddj142K+H1inXDZxPWz9CW/4tDZsn6v8gwUigOUDnhnXSrK7oxL9rsBr9xRxuKdSG
3tqTSQsp0ffzVECuB9y4zA6RN7j/3zmth0QmzagaFNoTz60FuOj2aAlGI94KgZmEX+Wq3id/CrdO
DEcE2nBofSQu+cxfZEPe5wf0UKruxpYiQTRgSwhyoxyoC/cR5RZ5wUhxcDPruC7DEb/H6sEsKtNk
u487TggsI8f+cF/tmeqOhNbouwRXlJNlJai7Lm5LAdn3gXlypuCcyXspABnv1sJQXDKeUlR4Tndt
L3D0yCtq6hv4DqK33JPqIRCJ9UwlMvd0N0jYZOBfLGApMHeoBUztReJsQD4NaTpDTA/PKYj3IlWi
E6s4fYsUyFYhDxL+R7lOYcbj1Wjev0vvFFwj28Yd59/wai4CCsvEPGLHqX1x7ffKWX7DEn+FAG/x
tnsAvqwN4ppBWIEv84uWrYbFOPeZBSt1PDOgWGw38oNSytnZ3IXGZ2D9lGqp+okn9ZOkzyLppppI
tjJlNLnh06pzN34K8jy2Wyb1yX9HeN2aDi9QuUtPQOhkokSm91AvJnHRZn7/oFTgRtbVxRE4+6ZB
tUmqMCpeTg8nSXZCxScDWCsGpYrlILDe9C1Hi3ev6h4OMC5L6RTR35QTZcNqPyLzS5OB2QgMTzQ9
NKg521w3jBiZnCCtOC4NSYpuu3ZkVFxD8pnPLNtjkRqU46KVsoBQXFa+TEY5oNuYgW5tNSqcowIf
+PvWFfn02nirvTVup3+6TdU1IgS5rSgxtDb331JO1zwrecP0oCjc05h2EtJw3DrBmzFmvhNaQb0v
8lllnoQQWJ56T881IhZX3SJdlYwwrEavjj4Ivc/d1QO/ZvBHi2jfjanhX5ldlntnmwXC8z2pdqrh
URf2ZD11CAOuZWSE2pMv572dDi4oPqWW94tGrDqA3KHGtkbi9sPnzWRUghqYdl2fuJsgApJa395k
N8gYD6zYLQsOLYk9MkG3AiHpMhcKRT42td3h3w8at4kuFQmlrechnui732hVvryD4xZU7oQL8ll3
yCrGyiomcTiChxi35iepVHzAgeOeclINpP5dvLKIy2Og+7tCbfQsWvAnMilD4Uy1LCBIRrNhZ8hY
9CQswkoOdcSJYd4JBhd7CLRVOTCLeaiMwkum3rjcNP1RGTE8hDTczoZG/MX/1cn/Km3peAJtO5/Y
ptaMcHIuwiOqe+GG5slyQHRqRvKxNYXBzweoUwbFdgqiUC9UjqGYMrKKC7FzppNwrlS0ox4h2OS/
TTLx8LkCc6xvAltBdwROTMble3mJ013DmnVSlH7DYsX9idiuafJkC9LdsNKQ0Tc0QgF1CLyk5RjR
jOYoBzRoEcbZq1RHFj/Va5oqAwknblKl5RTkw/LCapQ2f3zf6AUnHj7ZAuNDBJFUxr5X7o3g9x/E
qfWF00Y8hsA9EdD/vdBwM56eFzQVecfhcLkRDeLR9ViltClORk1TnhfHft2px/sRd+X0GcTKFU/H
keXZ4Gv2gd7LLgTVtmdw4A9MK4HjK4ER6dOgSnDngCiEY3BQoBetCc5mSyU08OwVfDmq9qLeq2B6
g5cQVh8fGtEoCisAk1JIksKL15p8dA6Sz/ocYwndBBnh+6UYADOcyPYXlFCw6NjowfdqzafkFTQJ
rT4K5Vcgvb2evRhD6u/G+HfGuzSmWabX1bYLzRy09lu5SOfmps7D4DgGHLmZupZA6cN850/5oi9r
HNUi4leJMrhlux02kGO+P4Ha3Gb5XDwGjjc5CJYRpPBRoBgTwv4U0lMPjNk5Ta9UNUl/wnzfZfiM
WN/Rz3bWeBXQR32/I9ujN8osaJ1XcH2aRusb9eVQ+K99KDJ5ijVbrBWySySeY7pq2RNt/krUrnkL
5b4zCyc+S5vWEAolzlbDqd44lXKXfcIpbJ5dEvBYmof3Ks2dZn3E5QNAM8Fvp8M7u8NeoM/MFyBb
uY0b0cX9w/al6dn/x8G0KquO/OeyZS6L8tc8FDdT+OWjgXlqErc6UWWmMcFlj9oJbxsi6FKZ/a3D
X+af0EWSNVdnw/63mJfdBkAWa6jo+b76tsmgJLdB9w5TUFhQWNi672r6EqKsECyfVL576T5Fnnrz
e3h+jHnGGcrhzfVcTbLDLcJIqrygr00A+crGN0s3KleZaxuftIuUadt2jJIC0uqIy+63b4kizHli
WJFeKD2Cf4Erj1A/aZoHIGhl9kmODEv7A+T2xle1TMc1+C9PN25c38iOC8QPC3gUHBowWZrwc6vb
0mmDCzJEJjx2O08pJsz2LrpHFI40HPfBsW9BydeNQtySU0ZoWhxJEsA1Z8U4du/uEHnxxKLtej1c
vpEHmGJB1VGoMdiIGDAJiQFu1V9c7sMv2Og+CwsTI9ARvQeucGMFUHhgM84DmYezLVIheMdJz/RP
SO9v/7JqAiSMH4Avz+u6kg+sgSP7tg+X60b4P/m3NAeHIa5txmrk/l+O2ODDXZIc/buLO5MPwZzF
q2tQ+OiqtOXLUwaYxQPrgpZLiGwdS4UHFLlo4PUOyzM1BW9cDkqolxbFQ9alF05oT+2mg0IS2SJF
lnGQ+oz8gt65oL49JQ3J9dLXgTpH5dfaVVu+3Vxf86i7B77p/j+Ozp70lDB0SZX5HgvSVBaGG6dS
VWFNl87VzD3+GR8YyeG/WB1O563P9O9VBplI7gMLGbY1wsBqgDZcsJ+XECh0PccVxrMx1Ns6fcHp
k3lyhBj0/T3187vD/w1OurhXbeBqtgwKha8Nr625MKfNy1nByURCX4TiA7KQktTV+bcDEimEQOh5
Xtrue56YIM0d0Xz8mAmxxE93rz6Ksp6p3xjVoqRET3Enmat/L0GW/Tv52QDIceyzgFuP3PCguhqV
9fwFKhSVZu9E9rPhYFMBk53nKb09o2YogJF/wddHpWJHrmC+meCcAi0j7hl8sh6eTXrosIz7uop6
jkzruTRKruAVA7k3QoXRm8ZixQeo0B0mYvTSi2MWyebNASlCT/o8lS3OSHP+08ZlLrQEb5g3wlIw
viSl1KrGZe5p+4ZTrwsDZBuc50jlT6xDSzW+KLKVBSPUq6prqyxnCqDywcjDQUYlCSv0qR19mcvu
4KLvzNoktuXsX77lU3NzmcsP7yq5V0TTYnjTlaVM0ZqVhfJTl1NlMAQ/IpE39sphWDR/TxsyOngj
hwYg0whGZCubiC4v46Gv4DLarxc8xJOkQ4lwPrAgw0IQVS9QTHkBBp9jcIqkl8IITRmNyV8LoltN
WPJP4UMrS/3UQO7RC3foYNSyzenU8aiH+5jWbVqJMcll4uoHpRH8qgYOW6jvv4T2+VB3wFOzfFZZ
pFw3f3dEBs18x3gHALVVSZVmYzIaijRWEvtP2/lRm4MqjQtqqGNoK3S7PtB/Hy4m8aLztj0+FWbf
Jfic/uqZMfn5vB4yBKvBV6+uZhB4yh14UYjYNXGjNZmajGZSxWOVe5s/23waL1A94SuBwYf+laVa
dC97sBsLrfdfYP2jHuEfTzxLNA8ItbQvUYV0kYcdN3WMad3yldV5ID0H00hEhCPtAyxLLy8cgNhJ
DIOFMksA2DUkv8yBwhe32y14G9kanD7Z2LRTaSLoDGEeWJ46fFUAZbLpNGi/2yDsA8cNgheMsvfF
9mrTjiBw04sJuWELQIHHhn71YhYdyDRl0W2doIG7wkKiZHzdVwoWWskARL8/BWuCeIMIYXsZNT1E
Ct7QsCKezSCb39ZlHCCymi9+BgHWgcZ+wD5As4q2b0SF63l17qHzJ6kfjLnipH9IneQhpj8qmCBu
vLgw3yvQ5jbsn54gH1JA2ck51uHWSebEae4S4eAV20zHARLV4fuUWzk1U5B7fRelyx6vG4GBE/73
O9GDhRjzWBtS7LByCIIwUSi0A6G1w0aAFA9Qwixenp5fBgs42ICI/OmMd77hw9rB8+QLeEAPile8
9j6JiQTR19LUS7ZwWk5FxAK26QxcLUOWZt9zO3jphmvyfLQtNwj663bNZ7fymoC21schSdSmQd+p
gyBM4wFEK/kvmPyGgQGondLK26rQt8o9UUS+4R59udyFV34PQaZQBcdPsD6JYtoR3qIVwkQsPOr3
cnki5fMrMg6M8X9+Sf1AgDJuujwGrSpGSBYRcF/dXVCrv0OMAffqDiA0KUYX57Lm5x0nh3Kyguju
OvhJbOwrDszDu+AsZEb0EXhPgYxBkgxSKtmWMTAm9wZEnhyctJLZB9HWVta+/srEST9J8A/3tEld
TYd11Q67ewuv4vYKm/squWO5McehjypbEQiUr8eXQhcmMw/bDOpcxXn4ZIS8PAGaVRr1iIJ0hPne
IBNX8fgntBkotC6s9yFbin6QGYt/OboextoAFdggL1ivUgDayE4oM3ODi6KpY8y1pHvIfQey+5sr
1KZKehvCUjwFBXjiSd7XP9NtrZS6uFbvxYZ0TtY0H3j5qAAEnZgS/mm/dRm3GXLGJ5affH3SQS5Y
5v+5ySu1rojIjC8L2LodxxP9RRuZ/Wg5uBIAftXnyXE4qKScv36xkb3M0w9kstHaCsdDswLxmR6T
tX5MOZ43pJ2wTsKlf6FH/ukT5GIijoMGswQPD/SxgeLBgW5Ows1u6enMLHA5XrfJRCuXKV+ELQIV
ZIlMFVd7JuoJDkb2mQjJm9JP44/P1QxvLZc1vAo1YWU/L3Me/llqJ2TkX6AUfSexjmgl81XB4rs3
NJFwohQRZJOWkRPbdN0bxFjHJYmrijVZF348TrzlgiBgKdzTzA6lBQipPIX4A7f2XR2UohDT5K2J
I+QqCx8KX5Gnzs8E06E/4nSPHZb1YYQEPROdOpFcyrJ0xEnB+4A5Ti6wuvw8JwxnHAC49Aj6HGb2
sAFavL5Be0Q8xOW32U1/lQd3XZdnpr0zWYPvIngJaulgiyQneSq/cdP6dP3sEwXyWzYQL1hOO8SX
Jwr5PoIkQT9XpcmLeT/5IV8qGuJuXB4+UvfG55iyl9HfUsay7kIhQ5+cXxI92JYwpObtxBGoq0pr
YkQKeIpt8Vc8GloQJ/uAehW4SMsVhijk5vcqormlvHlxI1hsK7zae1vZJePUQEPMuIuiE7RUzVA6
XCAZtWdF1OoOOSW0v5L7zfErWE4ZVVtcbo6VGVHA5u3bpbstrAJcptvV1MLjgYbESGIxBplNeA0N
tPDkJF1bmiSKMWdg32kAFLEEz/5enLRuR69A9Uq6zA83/F3v/lYsjfnWeXAUnzOuQhneFHTSLUXC
jk6kPcmqbmodoQn2saufB5Oi5QReD134kVNURvDG9nRwKg75ro0fyI2niwfrENqtS5hMP8N1j3o5
Aq0x0pb0kYX0Py5TdjtLLESCYOozFy+q8VAfg3ksAocxr6P0Fq8tddiJfNU/Z2EWLctqn5WB9ed1
ONqKBxeA37frtOhQIrFE8FWY/dmak1LYv829qTvyPoUBUiwu58VTDl9PqLe/wX0syzgv6Fa6CgDT
8VGbORgMh117hbE09+Xtt753cT6wg+GZfKA45HHIBBBOxAqssLyPX8CZ+umAYpsExb5esR9+CNxc
NPiWpEmQl1vy0h8KPaxrueoY+0zNN42VqID77TNYguK3z6mf5uO75TAjUBhJcJUh0dtlJvIuzY9u
K1DdKCyonb/QghD019/B1+AAKWG372Ctj6uz3+dTcyewtdDNwbErVV7/AeveBMHItX98tXbNIxN0
YNEv4r7GqtQdINVzatxVb2mNDd6Km3xxfBsKRRlmNWr2boJPDc9tLo7Wet4uX4ZH448ixVknYnqg
xg2t7VA/G7FEbf5kWhHY8yzwH9iTISotzpXjNvXsOyaE1aIfAaLVczQLGveUefu4/bEF5vfudg+J
Kv+l09Gt8LP089Majd8yhf1MhU91XrtGcbBM9q+6jAEA08jN+v5Q1qVX38GuZzwlCxrLSBLeIR5A
hfetBnuc4lj7f6Xsh9PofwNKCu9p+kH0731ImtZ2E3sadeBC1MOxBeb0e7tWS0G6KeI1RZM0/mx9
srKuZbec4zKQLFePhTahJ40uAlPkbDMH4UfSyFVGTbv9JFaCDKBejjyY5U56Apuzg9tyQbHBUc3Z
6PFeUlDBuUTBkZ4DHsKbowe309is2Sx6FkOZ854VoWF/uFt69SG3WvfLqO/ibCl+p+MwdbK+0vH6
tGlHJhko6qv0hVSQsTch9qLYKzYyeQTZZEBd5AQgp6fcqzquFxOdGFPPsTLfVvKb9gNA4gZmxx5v
kjKLEGi4u1IUrnyNilw2zPIilBDLIAkem6Q+rn3gmVex3sT0vGFS2RFKESPto5EY6XTzy/Xi+NSx
OVEJGDGTzQoSRaDw5gOzW+lmB2qp3/av43+Dsudp7M9DimWYJPvJShCAFFCerrMjjUxC4rLDV4O+
H99A2SKZB21MlvbICLCUAW7InbKRzIPucNEV57qHchciXw6NcwyQIyDojfDBK1L6+u9TvrtnbDHn
rpZJREWl52oKY1j4PVIbTMPEhRxhaQCjSXIzZzGgMd3KYzEAyHU8+w7CdRYLjD4zIg0xGiKc2Xba
r/Gc+K/lDjJLal6+wyt+Ria649RcfcWyT9RoNnUtDRdaoYxFMTzAOgMg/A4+2URQ+1cY1bSdMfqx
mJK6o/lhCSowXfTjIhuKaE+8e3NlF8SOADRACW5+q6LKpkjQpWRrtEUkSn9tF3HnCNeLndA21POc
yxJtYP9xEEP16njqiOPcUUHRp0ArOuR6M7HN73YG/b5QyuluWVmbizkPzBO5slG5YIcER598hh1H
P5BcmaVNege4BEPYSt3fvMBgfxRcWYUlBlVSLdK3FksqBPK7yd9B6VEVzcW7vPKnseT30icAQQdJ
01+Xt1RbBh34iZ9TuQLjqQEmk15MOgGX6bUDLxtrWkkS3CqDRc8ta13EUscPKTllmNx1C6xbFM+9
jjNEtiVtfI+MJ3FX1nOIQ+Os+dg0VlOFAVI4uHg/f71T7FboArPprCQJAeqyAlOsQrfeC8rCVVX+
Ho0xfxV7phEAW65Gol1Z2MEG8UmrJB6/q/9v41HQq1p2+O7If+YURLkKSXVkY0w1R5gioGUaF/Uv
C6V0dvzv41qWL0USTlhaKFGimubTWjJJ+5sjZkQUbrElZdbzWRmV6+o3cPycNrff7R+xG4T1Wq+9
O9gM9UnPXQV4M8uT797DbPtyG/3qYopUPRjH5Z7yUZfHZW28WjHUzaxCJIMD2KVywj2+zI/9bwue
rCcpbPZDCKqicUryGMkXnd2Hyy/auh/0X7yk3eR+WKAqa6MoM/P/9Pf63WDqK/h71edjHwGju9tB
49+YVDsV8PxrTfDqBYGruc7TYlGJnnETfuQSS6KjQOZplN7+yOSI4eCCTKTDMMGxfLiRaEH1Y7wC
FSsbFs8N4Socbo//X6JjWRdQkSOiYX7H6PWM3gCSFUDN9ysNqSja4N016qW0lE7QJL6XAF6PiJKb
eLlNbrtY3M31IgbYere5dRP4+nOdir563atXj5sUsrQceFdonEEKAtNPamPYy1hGoNOLhZa6NheS
jlapsgCcd1pZkhv+WXPlmlzAckp5b1bE+b9nm5LKSwmx1JuhSpG84USJ0B2ntiOgakGwJWRPHYGp
8OBXgtu8UDIOc0EXFMGrK56qr2q2OO4LyEdpo1smZLO51fLz0LMmm4z+dM2DRPpc5lBnsTIL0g/w
hz7hclSI77UAtLfEjp7WsVkxtR2TtBtbRB9jjMyM6zCYF4kB+K/UrcujrEioxZYKXrWd3Kz1FK2o
aqpu4CRssK8Ir0StfGYUfTqEyajkD6zgL9jSh1zEXLC8VfwZPW/idrN4dDPe3lLghl+WdaQZJqlC
bAjYTSq3RVX/YAUwDkHHdU/dKWr1Jwm72c5zdLRGq/TWG8JmaSgTuhZe/SKuyHtLIpCuAI9iA7q1
XUlXesymuJgcLX7/D3D9IFYkSsArBrF7sZzpSYMIhuOoSsUlJjzBVAbijV9NESPNesgB71LbIgfT
qfIiXk3mEwAmsoqTNs9z7p0NOYTg7KhJI7JLa50hTIpiGd8mANrMsHLt0xQnHqFH9C9xokt5CBlN
H53xAgbZ70wH6lj+1uYli7A9VrezSFD0iD+bXPXbV7/RrS6y2iDYImzIhnX8+0gg5Uj1Y8DHRyoB
6exFVw9vD0p+hd4fG9FzYvgCWRIQVaJ1jIAs6nsj3hI2PYqGKv6fkWXOFkOyjz5PgEDM6cP64s8+
uf99DmTianDKqYVhSwUtHrFs0lgAEWkjjtb1VEjPLUfpkHBgbaOkdkhPpWp+jgQfQzp04M4oczWv
rxkpA3eKjKUDEgGQpuyjN2roWH6tS/4ilHaxnQ3+QmyP/LXLr1XriiyiWfZCjcjfreckyZ/SgNf5
s05zogG3uO95P37f3LN5SR3U/LPvt7ETw8VOtyTwRSh/5qsnFsf5gTarKDriHGyvRrqibdpYs4j4
GCexfULp8B79JqJvve4vUGeLwfC7i3epC3WBAjIpJeYbdzKzs89zCNrU5+7MkV7s2b1+aaAMkhUT
M/pDFSe32vb+fCHbGSIr51wg/KTZaYX8VXEvkIeYX2AVzscT8snf+d4NlaWOxv4wKvTRTLTV+Ntn
kWagcvrNx0LVdVp9cg3XG0N10f5KoOeoWB29Dsv05AIz7ymOMWPLtnli1YqWVD6grnLosswDYz/u
8A9C0CKjznwDKrLQpAPtvckpHGPNzc4qSrbCnZzXquAC6/dvmckZ4oJVfgHHV6GftjhZL+NV0Y3W
tiE2tyumg8bgtgExKqwl7uYv7+6HqXMjqfcHTWLharyU67771YO7R5IyxlZo4ICcHYCMB8aOSCqt
iGKAiVZHfbHTyq4K+S9jJ+n0qvSy4ghVCy0WkAxP0l2J/XDo4i5xN2QMR4XuUgP5v1vrs52t8JTZ
gSOsTNyzw0JdWoXimszoZwKOKgBJl+EM7KkQQdfXexHv4ZH8jjAq+HZO+BhESWlqDvLV+ZR1kigR
SdPmUR9o9PkiOBbTpn4+FbXe6U3otOKOf+Nc7J63p6h+KRQYii0gNnugV1k5QShfnHwy3w7hS8b4
kaAoXS2i2PU5fW6/HvpUzNJ0zKN4BjmFKoqe4NR6eN57w4dWeiuyjTLFxoVOBBsyZmlHUXwTbv9D
epkdYFh11xvcgt29TzK9NHPMSTzzCRWdQwq2rDy2wCKxunbTZgt/6jyj6Fvrf+7QXK3B2fPSpHYq
KJ/d+TTpo3zJH14STp+vhqOtJ8vt61C6ixBUvMJy4QvNP5E72vBOgImTIBNtKP/IYiDqTVI2r3qE
j7mkS5pBsp1nojcGeQbSCY6pg1STtdDDq937CBNMtFcX0Oqr+K548XBErT9LfRTAxYZCdR+jYCJh
sIqiyA5gBdlQw5wMkN1ng5/EBNiYuC+3HICjrI1kTbCEvW17xVu3Sc0X+CA874yPwXth+XUKgnc3
mm6hyO1FeZ7ZJA3nbcZbt6QId4syuBh+WgobZn7XKdR//cyBXjRvwaTwqFu3MUYnbPsuhD9a9Y8V
q5L97QUqS98saEEIRjNiImqnRwusIV3FGIOxR2cddUUNdvfdPj6GvYG/6+BQpNjpjvjRR/FVwQHp
H2d9yNfo5ysc1t/9u6v3Mz2LpgGU78NEt0rn6ttcxcljtugQHBrY+v+tns1e9UFT4SWXb0xBcj5+
12GeMH0Q8aAf/ey4KGqkNE42GavBsbkbmkMfKlAGYzbScSbIWATRMClQscD3uevrH7oz7BZSQrqr
JZ1rP5wVTXuZG9y5MGv3ZbksjsgnVAarGbZSf+H0q2Q8NbeGbCOioout5pJ7R36GXcpoRv8e+ZTX
2IzhRM0rjHA1d1v1Edikm2Qy8Ss2Vjh3y99vM7ti2ary9s4mwFuhkDu1we/+jI7V54Y0VYzw740V
mneLUNBCfE34d67wGDv/C2YGkdKRDJE3bl7ALEyS9niapt7FP7RbxjgagMXiJiBn/L1BQ+GMj87y
2CAawcCJakSuqV5fRC3IEwVaRZHLHPG8/IoaBUHDlVKeSWgFsst/KYolGEeM+LPA2xRCrB4/rXoO
5xXPjBXlmEwFYRvaeLCIbIxm6sNDQmX/ulnmxEMszVe/NcCyoazvipCSbjHtuiixSNpw06H0XSwA
G6c1k5NLrb0DZgC0noN7Ug7El77Td2Wj1sXLCLp3TxQNRixGbP5QJocCpWIWy8UOIDuQazpIw+Jf
HW7aeaL3OJX6lm0gjfOdKbWcm+R0txB2D1EfzNG+Kf22WwCJDdh16SWulRXhk2ixen/I/ZiHccgy
EBIuuYcfHA03kkIwNFCG1EEZpaRhxBPJ0M6cQHoknKQgRGzA4XFclBFTqj3e3NB5HeqEY+5oh2kO
oo91cTp/GwK7pfoRk02NeoYz8eFgV4sryzbMDSXiRZhG5R+BtD0B6VSNk9MKKDDFti3fGHNT3gCj
rIO+CBS+CYojj21VDIo0QD2gdJDYBpN8jk4/XDjOsTEwbNo5ZrqMirttR6Rdk86EKD5dWBbnG5Xb
i2lWxlKivUX8LlkCUNT95E5koDnYGsCg1OgaGF99yuR/YNe5du6QSRRv0lIQpNdRomQQddGOCwnO
EU6Ym6qt4qqCi+NYdmgio+Fa3hYnHcNaddbUYfPa2Ah5KGpfGszUkD9lYyGMHtiUBgfRCzm9PwYK
XQ/bQQ/v2GtGbEskOeKmJXuWOxWKLbxSBzKICaY0MPzUPjnZ0XHUA4ZiM6lIRA1ilH8aN6WPAVei
TELANVT03aysJDXWoW+j1P21KeaZPzLk+u7Q8d41fLX6u8snuOu41TuWmQt8bLFnYoymZKcjhJCq
V2c/wDjvgLE+WnEAgaxBY2Uvj2GIXraCg27gOJ+lHMdu6lY68K2Orju8yrfuap/7cu/eu1fmkYVA
eF2jCHwP4rnVKiOIkC8cAu9jzxIIgZTUHx0vDIOoor+Wk97UVdtS0LX/IX+P8hNe97nt5B8dXqQL
0ykvUxnVeXSWb3Irqoaba/rgyWk9YWuVl0480V/pYpaZ1X55zhzvfTlUAm+abPoRav7vWKwXrExL
OSptB+G2ooZC1nIC+4NowlPAdbJDdJFeYIV8+Z6uy6UB5UlwYJpW8HMxKhVWVeuAFuQz3fuRYSv3
XpvOw7x3Lf2PtkKte+6H6uZ99jSJjHHRLq+fkDeGweZxuIPhZ+g6rw8C/dvd1iTuVTH85U94kVlH
QJ70xMs2A7gvFBIVfk5NNMicCH6ueVQFQpEZuUWgKu1CCwpoGLNMxG1rrjKTbzirpdrGhoyYU9P5
+8SEnD1GQ8StMDSPkxsLbz543cORutJiPiCtkWph563QzKZ7dURf6rolw+qMaCvKC8K5oLG6oCPV
iIjGsdy3YsH4yVIiIXE7A8lVIDcn9Fwkzo9D1bLCelD3EeSU/WPRszX1TpXSA+FNPzpJuipDvtUj
bMJZrEfzWBPT32kch0F57T69JGw/VjJgk/MvJht+M1ILqpItJbpfRqYiix3Dxo1TgOOpB97DS8tB
e0n86w6Bg1D7U3Cc6IlgcQzQwlv79Nom9N6nsyh/Buma6ULt/Q37gROUH5kSckvguHH6LAOLLeHd
6LEadh+vpQEeU0+NqHhXrNZVuIeABTfVQIFdqMJ2WwwPHQ/eGpYm2iJ5gQH4nOYSBtSe/GxTsg9U
Y3QdtJwLrvyzRBjhysAjofC0nz7SV56H86wnhEhwo6zQ37ecYzcR280hkNzXN6pYwTPGBLtPa994
BJD1kVcp3YluB0xiXlnzJklKDcDESAWgAVWcB6mHQSnS7GEU1mLjuQpllWvVziaKdGAHsabXL8bi
+mp52QGfuU4qSOSRMja1hHP9RGYogVIcFlJ1MoBs+2s0vH5HDL50CPK7MUmuIUjClwNuVFlWag2O
PeNMbmyGoIEA1OQse37l1R0Sp77A9pbhjfpKUPgAne+OpXy28aQHgZtSBr5O+RjUyuoOtQ5oxpju
l1i5OXRSrGVFfQ9qYmvuRfXnDCH6KKwUA2qb8IUr/nLg8ERyYHjB/QAsmt//zFi0KShcv/NfHUez
SeuYLJa2fBDjJvC4n761ql06sXRwR2NIBDi10BDHq1/Lnb2dav27YqAeTO/AglvqYPbnV5P6Cr3a
rA2FsOgLyPRmJZnDlkRaJG66Vf8AuTmw4+PDfJnJxLnOVX4c5kn3SXdF2ILev/PWzzxvNFgKXXQE
ay//gZBGHQDiddeR9VV1UWHLIcgearuFdU4Vtsl0b+MGC+eKGTjsJqe9ESjWb+bqtXCCD0jEJozz
fk2doTZG1TGi/V9fZX9FdlvVJMTiZDglbtwmlX0dUDmReHdBShnQiwgTW4FztgBv+q7syEFTqRZF
P6CoSuG2DXeVVuoXv3DMzsP45ZNfBJ+5Rb8Dr8+CpF7vHPd2NIbgfAMDR3YqMD+ApnW2DRGzptle
L2iNr+P6FuO+J1QZsIYk4+flSyg+sDlyv9HOpTiBPtPKm6i0ywPK4of7NheoBnE68v6qqwhotVMh
YTPkoa6ZaVF4dUlu0PByyM7PBaCxvWM1epCblUPmodz0wvr4s9jL7/TPCDes5Wy8VuHqTrDgVE+M
4rPnn88RTdIlG5Xc5GjSDUFYgF7jPGWwsyx8omMuezIHkjQul91N2bmNdHQswfgVrQ9pLiCfGXLA
4TPUGz07gB7NXvWpffW/ORFfKuQ5Y+K5JgIq8EjBHTr/F4Ws3/hTVhl9GcsJPPD9M8HGlkdrhkdU
LvfU5NVMFlymn9jNnA3Vrv3+L1GDsaE39ggkLcWrwnWv9T6rCiXwWGT8jsi4nVKinghZ82BozPlX
6V3RTAherLoczW91Eh6O/o1L5b2BiPX1qrA14fVaLHcUPAy9YRetYBRxP69mYzZlRst3cnKyFdaQ
j9ioOGSjiyzuVCRavkFiw1zVtpuQ055JruDG4LgfuMOTr2VJwa8F2UoN4P3ZBML/N2ZEPap37GvE
ENaD5yz1WLJgugdUGWmlvo6nZ5SqLegSHnXunJwR6EmWaMJNZwhwS5WSWWwuVQgJTlkZIrKps/TK
GNR/7D8BztkA56F2UuCnEffKudvUZrv/DGX57fkK8yGrEkx3BSyl41EjN2jEm5kAO+M/K/Vsow0N
RhDj/TW0zBuvNL+fyksJPloP4MDmNq3r67kpSYrU3ZILiYKFM5k4UE/UbxKb/rNfM7nR5tf7ZK35
VX6FgOp+NFSz119y/krtEXAMVsitR5NoZkwt0n8WsZDUX9ROi4jwP6NxV/GksdvgoZ1Xo5JW7IOR
9311F49VBuKCyPbxdsoii758fDC64LRsaS4X5MdsYE5xVeQuxZowMJpAfmh2rqD6jSSTQcwqM6S6
WVelLyrBV6TdSZMVss6m7L/fk8X+7wmQ5hGYmuIeqJ17O/knEn4cVdxq9b6rBKVIfHEP7TkaplMP
Ta7dQZResR2JxTyQyXr7LkdesAbli/wFfvqvxnYkVEcYlGbyS4T2TIl3dGTsQiEzDLaAHynK+Roy
oByYkcLINHy9vuoAWXSypbKxxbqlYkDqZcPY424Nu6RDhuuqLsfXzRA/E75gW1bKVfpJjbI8/GIm
JXr1h3t1bxNo7llFQBmccq3DAla3bV3ACdUEI9aRcreOY6tyYcw32az9QaLCiQ55b/cylZB4ODR6
dhyf509yKzsKO3Sndt3I377C9Xo53NmCOVBdYWszEmPMYtYivvt9l2ZA+zOU/H7ae9mL/GH24GK4
wQkIRBaRZBwPj4cnFbI1NDUv3puQ91poLUbTxrIhPiI0yBfonL5BTnCyyUHa5IZCnv+i0qyVxW8R
C+WQaqA9/TelXAIFs3XGMG1VfIb9LpCl9T0/PKBUmfVVWyRYTro3VFvL913dt8Qp5/rZhw73vytn
YQNTXmdA7HzsVEsirN1j/F1QNVMam75gLeOJl4t68caSJ+LQJyQgi7VaKmdx6+lVNp49IgS6gzUd
q0/MNOQWld7fBMlMEHdRXmwLRs/exP4Fd21CFSOHfrkKDGpUs9v1uIEjKZZEpofD1wYXSu9afJS9
8N7L90lQq4nwib1gSpn6N+4sj8wutEothMzlNxdIZl1440FeXJibeEFy5UE1xX4kqZwoz7AtyGYP
jA7/7GXhlTYwIO1apCXH/tO3/PNI7hh3paG/QbRLr6WGunnhKlTjwv844dMMuEKwFzJE2t4CGWdf
XftEtbZQ2QMloplpmzq27aSxRKK9T+0HlSAtLWEYD1xfAVLMe/QIXFndjPlQHjlmyEoScSIVmYQE
pplmZfJcPtkE+rPy63TI3gx6RP+S70f7MLgU9xMR5E1hNreM8JQm/Ci1Z+APkonfKOXXi+/jQF9q
WKnXxU3ZpUV+7HwQ71llv6oQ6ghFAnV3o2m/GQRDlSS5U7DGPSM8tw/nHr2M00idnc6hhMqmeDdV
Ex+EQ8otNTAEmkJZXnCxhnDCcayWzedQkTXFmNxR87SFjhIWkXFR7Ue3MTmSVUFksE6m1a7CLM01
mNXjoO3ieY+bl/y2YHogZ3Azkv0T8vUHyY7M4ohut+HWzlE1ZXyguw0AeEkNGNBf/nEjW/bfLGE8
gO0q/SETO0+8eCrDm28x3PMWsWv/+kThlHn/JgUSaz+TbBgsGIXPvZR3zp5HaK2LHLX8C9l46JXr
bxTcxlsFg4wLRr+egibjPDp91toUP5orqs1uld7S/9X4xTZcQcB3bTW+y7EWbipN3MLhI10+Z2to
ciwg9AKkhA3ZRcJXNz4MwsvvUVtYNM1GxHBU4z/A1aOQqbO+gs14R43UoxB1Cs85k6moWJbu7727
eB5MhLPo5kEVk3TevVBrhuOmG3zsv7C69JhYUUOXx2hm3tJg0FjoaPrnBZP8CqPzQjcP7Me38/N9
YJq7xO8v25mWZEPXqNJ3tpa7Wql0vQyct0hUGEB8Y2PfMrRBhu3Nj7Oih2kUC4PJEGVW553vHfcc
uROHAcWUuO/DIPptJo+VbMTxfEjhxQGxDuI5KonSZSv41XYo6NCRIfwVZ6TIQnr6+SeK6CdC53fS
0U0TACNRm8i3p/gRlyJ33O1rLpEbJbzijHEKKWFNWl1XZt+8m8oCMi6eZKyNLZQdR8TuD6YMc0In
5g1RO/1moOFa8KiAY2w8mc15MxBHa34rx7X07NPkc22NckWGbbe7eXfKLk5M9xl64y+LN9hsn0JB
ln6LqmIWMWjFbih2sqkLdwhJAHEPH6AVtvWbiyycowgNTLDX+Oj382o6ZpDijrOD55JpstBGElOA
gqbnIDeQ95JqIo3wsmuD6OP+LgSnOse/h0QpBDwLxxVb0/Ch4WYXpUyjE8V386+d+jJ1Qxx2n1Zc
zSoyhAbKLRBwrIwTE8tdUIoSRo/pfjoy6rzTpuDk+teIxNOcwiKWnuc+zqCkIPsv6/YkMyrpETLo
YBJL53FrWlKrfel3+nbEVnd4AagDCB6wVjZp6OKiyNzlqZEw/ddknsLS3qpvhqTGHPhr5IFD5I4+
4ta+B45/J5nWAXT6ibQSnjP5+7RjU2I5ejjG5chws1Rk/DhXScvLPyXk/MnfBNhHy2Vy8xEN5Tz5
r7BS3UZsj+xf3Z/cC2ZfbQz7gX/c0W214ryY467jmVmzdVintNduGxSUw6FG/zA6aj3IghubrssC
u0mP/DYANTb0OvZsn3zhFAFjqso7Up2Jif5x879jIx5KMYfRrZTv0Zu/1MTpP3rtzc8q2aAKQ0oe
SWuRpMqA+hUdlZMBCAocb5YmMhCLAHVwcivCAepVZ4CAhDy3uURtxtLQ9H8qgqWdpEQXGCGUoaPb
2yfQufo4rS7Owu7w+UesiE/NUZrckpnW2HjsfTePUJUdDSRVOj5zvlk7AtDgxwuAJnTSasSr2zbm
xqWVYr/5YfFTnlqoX55VMWsvF55zUs7cwGn3ZupT2A7bMBIrdLtrIqsK6fQeBiG+jqihxGQ7gLiP
vhswfp46i4t6+o/sDGEFqvY9GpsClf90AYz663QHFTpAqxZHAFD0Hlfm+2urwDZ1ch+/HFVd7ZM9
rLxMw/VzmD+0SIuhSg5Hbk6SRV/P6xgzjjQaLqlWohesjVksrbSyrX6USTu+eYODz6PeuRpjUAIl
gGckYZ6Z5zQI1Nz8clAX/8s+IUQZMlq4mvs6Trf9Sie/W1drKypx9R2Ob1b2Jfke4kPt8UMP1ssI
EDF+kdM6JOLxzvS3otarnlTuafpdk3UFZbrTfdVPHjPiZ/jFIAHL2CJs9WeyV/MHWoknIiQ/xQPv
uO48PaN/e7CBeKbLqsjTph1DbefqVCz1AZNjgbeiLv4mF8X6g9bAVv4U/HB3bMxcYkuGTd6y6SpT
ABwqu4K/l9YSMExv1yiiwLI2jC04MFHhXQOnXzawmZYIhyt3pAG+mTHyh8s2WF4JQhpyphMfbYxS
/r3ED/Wd91/err1ifemi4YJ3OC939ZFMDijbpWbFCny7Ew783bWDwBndFMqj98t+z89zvr8rv14p
utw++mdOQ+Fco8TQiNXDb6SY9bGO2E8eGk/fU4wUHQYU7bLs8GbeA7JjnVnJ/MNG6eKl82A3WmiN
71mQEdrWWLeDI+mZBm9xP+mh3riDZcrwwKSBwGPRaIxoLvRgqDqxTSsVF2v0wT0aLwIZuJvi3Tkk
9WuzmPsS7EsV1tIQRhccFKEQSMuYdSXwGu2+gBeEC0OCXPrUwzcu96T54PPJBXU0cU9mN+5xuO5P
FmzWg7FmEkjJ7SQCiBvbCDZwePQu9YZKvpa6WF8KLLnPmFnxfHrjiRTrR7dM/xhsy7zQnW9XI6wL
UAZfqBhZYcJNp4wnHmgNjzIU+gjo/rP6vETPO/wAL/c9ojf/dauT7+PUa2acJOVwyVDQbJ6/g2xI
akedgZk618VTKhLCg91DKjUggEn9WikeKhTCO83cemTRUzWLXjo+L372z4iF+8Fy8IXyuCczwmBn
RikYMf4KGRFen0cWc5UR4xzNJRMyrgO5fOmbu41yoRjrOOvP0ThlabxrP0KYcLTJTQUVTWJNFvBk
FYxqk+pdCE8GRE3dkil68+c9Bicn4gSVyLAbwP/Y0ZHx4Hs3EYpV+wCnnk0X1Jy1aA0XlU3SSkHq
F+6ivm+GY1fN6eIRoZctPydWvFQeqIMlFGvy88Qg1h4ytvDqlkEP71wxK7agIIWt94Jx46Slj9h/
fcM4rSAiQ0nmmsOIOwSIBFH4rPZxLUdZ4qeS16whZQHaZQ2143QNUSt/z1ydeeX8RCO/44LzeyLA
nhEZOLfz6nvNDKTvN72lZ3v0rODE0CCfGLo9F50LHn9w53KZButNY69/roFUpv/JSyQ+2UEqNoMA
244WngDlVZex8OZD4Ru7pi5hiIcYoCIhOxnVk9uyCMp3Y7Lfe7fK/d4gR8MKfj1emXg3J2WDdtKa
FPgpOp9aOGJfLRw0Meg4wq9MmL6j3K3sMzQcmQiVVXNGi5fOoulGCTf7KMrZgaNKSw/CqNHA0kdn
qFtuQB/f5P0AGvqVcYc6982ap1VBnsp8pwy6xcaoaYGOmaGHTqp6oLuzBod4unKvLlXxPgY3isS0
KhrPwyiDqbDUpUEcjEuUUpTyn69ogqdwICHb7eGaexjYRrNTbyao/Y4aFD1UUg7OPEI2JN7ZycCF
EMPvUzcS90aAQdq5tSgvoQZOEfMWX+1eL1I+7np50+08LEHi0lQGcUXzGcR3I2ZCxPt5Jj2LHmUO
x0HrnCc8r918eKkP9Z+CAMtL7jakRiSvfQTAT3eTZUkib684o2UOcdDEvXmKldpl5yjwuVfnkXPl
IQrrduciQss0ZToLXgrORfDlcUop+NaoxTujZeQjTh69+C8gSmSY203D0WbBnF7r4Rhy90uUeFP1
c9Ss5BGjr194iFSBkR85QIHmRZs27H71DPL8GwZi1botRKuetUVntY1pexUOx1Xwdj/Q5VNkrC9F
eEA8VL2VLpboOpmuno+4yFEP9r4TgzVJXKB290lTSBjtDgsiwajlbwV5rPliA8lfLUtk/xxoNtjF
jC9hXHe8prmFXbogZTvAskk3tAtTaLfTkB6V26mhZMTxAsxVnDY0Gllzz/v/cX7A5ct22sMYZMbD
zqczO5DhM7ZFwu/+1yU7rWUNK6FPP0DqY13+10RQagz+Ylmh2vOvaxHyhBs95Sz6ojnJAQi7H8z5
Ewss4FfO15Aie1LBTY6EJQ+Q7e/gzd92IzVYzMaqtNxBe3vvctvohbgBE2h25Lepequ1w4PE52lc
tCad5P5R8VD8BOabhb2mx9DkjtSrSSBwVbbkNO+T9jsOIaLq5dYlVU+l05geNzfioLKsPWNs7nSj
oRySOmCQjaF7hOSaAXLGPTPyI4dUR+xpZNGPvgqPFQKR41eqNHrofTc8FUOYpzJ8BoYCVTPH8zBE
oWb8W+p0Lb9Ytk6TVSD+rqUpaqis48fdAjoQ0bDZBhJO/O/29/c8PAB1v/dZ962MW+TBW7/JmpZR
P0XfEoDW0/ByyfqS7P9ONIDA4D2BiB/iBHXN998GSDob7c2y7EQGcPwZLg+JyNnl5aOU8RtQ9Hcn
lk4A8weVTXU5eXteXspu/swFHAEkZ70nBCgol2K7X0TeIgk3X9z+tH/QGvJ9XPgxxhhjeDog90rV
Lyjkz65ZCoHjTd84Bq0inFzF/4GHoycr0ARXUtQc142woQcbKIxfK1/xw7RYigDPw0dF6nzCy1gG
TwI5A2acpDVlQbqku3SENvpH/gxUs4P083nG8ZPvikfoWnxOPjN7tvPVxOkOxFwc0HqkikC5tWhf
SEognMhn9r85LY/SG6es6TlWbuYIkzmjXqOn9nkK5bOOVwLFzAzNl5qJJI7CsmTIyie9Ms8n6XgF
70dmEqgZtxwIpFHf7KXayqRkeJQKD93sEzDHVsewn0wqXbMFDeIFZsfkTmEmlNJXqx9iLL78bh6g
L3zOXCdaC8K19ORgfzxigdvke2acYDfodNExIbClrMdPNtIRa1NzAdd3h2dQUQ67uZX0h5Uoedmc
NP2aQRiUy3WtLyIQvG09EDJmVChhMabqanZU+KxxmoDuPysruxTEFDKIvHpkBu197cRD5VkuN4e3
e+rpJWsQ3SjF4IVu9W1xNAHV22Q0WiOcFz54uuXkAFqVWrpG2J8e3HM1Z1fGrlCfl80UL9ozNqRa
1ZMCXYOMDfd2j2LYmsbV/Gsc3pFU5PYA/+w1B6hWVqyfV16EeNd3viD3MmMuLtKyK8a3qYQjIhsQ
g7BCnTZPAlI3xNcHj56WeciNtKTdTaXJ5Lir91kD9FJZFZgzKddfB/LK7ECO2o+/NbAnjLLrOM2P
kiUItSDav252V5u4lURPlm7KSxPsdIo4ykZuGZQ5lytT++CU0ajsKI2vYOMD55gPNiZQyxWCPkab
L4OyCt3EJTWDOVv3a7Nr6cgWr1MdDYTYGuPksz3XyhH/mtFWUM/g/SYReJTU4Iv5QUFf2H0nao2k
QJ3fHWlBHPUqNNyoLOTV4qWTHqcR1XhG6jPDaSQ1tVhopt608lwG8KpJiGoNXXEY+wuaNY/cax6W
CirYq+sfy2+WYnlduA5QqkSxR1cMCOJqAnG0drHYR51aUKkV0dkbnwptn5rqy53lKR6hS1IKbC0f
JNoZTHwJUK9d4MXEwqMvCkD7kVGes4BEgyi3SR/7Jac8KYioO4/u74+7MicSv44N5dA3+/Bd72bK
SrNLat1bZ8JInhSwYp3ttlTWZvo0Yw82d8IYJQW5M5tQO2EMpy0HVwQmY05M3JpYTFWaEe0nwLIU
XJzI1pN2wPPS+jsfRPsgf06LF1kACf8bvnpAylhjCRqMqDsy+2dz4Vgkf9+NKTIcq0p+ihmasIAE
HErmAAmHtJa43xUHSqxqyZPChv1TPUbBC1POXIwrRsCkvXJ5KnbP5T7atjEBikWJ1aLoLvFiTNXU
eFOsS3v78Yw3Yobl5IeEPDAXD0g5WC9L32AouWtAr5gTeNFd3RXndcoh8QAx2hMN2z1CNMdEAXiV
MzmaTnZqfQ6z6Iw/UseSl68v/6x7m8g+DB6YwuU4gvRaJLaRS+FBPMCWjN67uX1qgJOCnG8G41B2
2yaYP4DI0cm1/dgDlzVTD+vzSQD74sDKOUCOeXW7qJkOPyrm3/deUQi6XjUx4pa163GMw1i0OjzW
Rgg4qsJcrTKKMeRhGkI1DK9h/QIPcZbPATreId0/fNclp0RDOlAKnQnzwofgYm7bsxiuIDeo8k/F
i5hV99vJPC4ghERkjrl/jo3gBYeEmvuKwh84Jpiy4xhdJoqv+0Eb0Tnbey0cg4GOAqrXypr0vQJi
Fb4AQ6WNGjj28tOYe5A+lzzDvk/d7ruo5zUHWI+43xHncrr+ICGQZeEBzbId4gu/Ar4lJc4+eLhx
Yk8iEKaJvy0SeR1BBgwadIMTHB1HBnRj83lrVnVT+bf/LftNmIcBzsXJCJ+oeRdzF1lDFoE7pkqQ
ZsAsN3KvZDbPSRXmcavx3ccmcko10n0c9SDchSDFb/YgQCw0UoE0U+tdriSuz6gA5IWHTLX5M0k7
wl5sxZdArR0+fIKUCRE7NZDB288K8mrUoxu4KsTx3qY+PaHwJa3dALj+nOQ0rWb9B5QNeL0Hx9xw
6Dp64ElhIx2pKxM13g19Dy5xx5xLkeLAavvMzUQW+CBL4LZxLsoLYiVwYPAJWViUaYlc10K+GsVP
26y4yMk3QMHx2OUzBuYDS8AWTpx5Y4FmmcM6qagm63XgqmVg+2/+4SAFn5QHU99GZ9hcEW+BcCoX
R0vBxq7v55EsHX28P0VoiNjfABk56TcMsYf1z4xZm/Emcym7DWevNkNSLDqNirVstQcT1s2oJ/U1
/AeyugDd0gDJdmgU482H27RKYQ5LiVXEoqawQSrSQB+9HoOB0AX0LElSF+U/E2mTjRYzC5bb0b5S
9QpGgEzWkotBNga8fkcodCcEOGbOzgvzioxJk6oOL/dmm0+MEHBmsygivyghAhVPasjxL4xvjML2
ZY8MlolTifAsabweXz6BEriXOtDa1vaxhAMI0hiU6ujgnb01HtP5U/cnFp77oRT38t2rAOlAXKj7
njp0T4pgIGbhzKqUSrHWOTBEwYqS19+0Fb+oq1Mv2dj7OdLhDuH3omrQBshBG68jZT5fdJwtfDRp
vG5aDBzD0Q2qb7BvQ7W/jQvMxg9zKexTghm2wA61KCPa3LxCZ3h2gXbPodUjiTLmhVRtV6jikeyN
mrkqBx27yfTlBgw5KQNqeQ0LYBN2mEh+2ScB2efmc1oLjYoTlhAq8Uz2xDoLuFFeQuIFQL6EVmkd
T+0zM+uRbBq9DFJc/Cq9NLQP9er81QuUlAIjT+RFmT7gd77WlD0tjXUO1rDrUbS+d1iNmsSgcyEZ
UOjzwdlEym7NCAR5IrX6cVDka5bnQsXlDZZWmyzk0F3o1fPVVV1lgdckBdN2ynXQEQlu+X85hLQS
m1FP4bT8yIWaa7TV1AaWXI5AH/yw0tADYoiw2jNK9De/litsWaLToaalrrqWHI4LoKmSOQFAdUnJ
UF2Lt7nv8DFCT7c4iUP9iAS+rczQp15i/eFHyqpYUVlQ5EKl7JJB6LOZ2dSaMl39vbwKd1dZeeP1
IaLdsilolWIcO3Phpupg0J07nOi1c8nBCDg5CNSmAoDfxdzZR/tibmhRDVQ1W/zQTO5SMSdMUWND
KEyY3c2jQm4Rl270YiBiRTEbI2VTNVZO7Q/9fswVzK69a6EDWLdYoWOLNbSJP/o3wR/eq9L6vUom
4omYjtUwx2p++EhRC1PzbuGE9U2rgwVftZ1S7j/kyKgGnIN4HEAqzobKLf95lCDLRLVHSWE5WxX8
wgqombBgXVRMJ9tuKDiV/5ELUYuk6XMkdkFVrVB1W3D6Py6wHz3B7EBy+KrhL0v9bAtEmK6u8tPa
GMacHGW0hxlo/xSo8G0rpNPpYIehwwBRm65ZXyHSZT+Tiv1JD/Qa0PWjVGXxcmaIYOR7dsmEO/6V
kTnlcoSC5Fl/wIFbNx/MDV7RRxygDID9YLG1ELwhMB79/j1hyy/AJFirE6DyMXSISAEeRBOLQMCw
804th5/IwCiORlznQ+SefcSXBkRreKZ3SkRMqxFu/SxD3xf1kBpPVPJ35piCAX2G8SjsxHxBmOxE
4QiTO+vu7qg4aBOz3RRsNcoVv3MFNW+ESHVl97eIr95VG+XPKZ+6yjlkZf0yF1Mpft4ad0es4+h9
XQqR8pOmQ7N19UTwq2AnfEPGU5tOmLeGIj0DWJ89qv2rhi6u8fYDcOK3NtQaY39fXZtu1wVsdezo
mvHaZ/ohyvNPcCiFwITCc0sZX60om8ad/CCvYBye1oKQxnc1qZvo6YqfyAysDLNCcIP4cOeQ47ea
pD5w7HZ8Yb3UU34jogrfwhkl4xFzeGbJ/sVazt42C7NNl0Mxz2R50UKst+mNIzDwUkFCbjqGAycd
y78gmMGeWQgQ3VVjzWtIAiqcLzxWDmBpvVIXwT2ucZVhwN/PnDnydcj7tfZiA8N8stghmOilrDrS
dbv0IBubnjxFkgGPPkBlcEORII4Q+Ndc0gH53lxnbHae19LFUZSLkQM83Eg0wavFT+DlAIBqJ/Qq
spT6resgnRTrYmQtCsq5BnhIkO65rgaQP6dbTHn35toEjPrzw6naG+vG78NANsqN91Nzsjlxbf6k
0Q6HlqQqNHB4qEwy7yRzE4XcBKgXlBgL8Y297Sja86t87d26iETWeYnfFIm4E1cknIBxB8Gj2uCf
HCyzI4D8C7AJZ1GhQZgr764On2Qlur/ReM1uHY8/kg420fLCS05CWfNqDdL4wfXc7pRuP/NjJrAR
Qs4YB/DnpeHhjoQNfwOWsmbIhVyY6k+9BcyfSOIFnaBpYfU4Widve3GOf/uuBa+e7JOrPi/4pjC9
PN5SMLVTT1g0BYhKJrSN7JwhofCU6jp9l3jdWeokF3hy5/2lXETQLKy7OOa4UYDPG4zfMcQoXRri
oXZqYK3+9sAEHLUsU3x4+cDKGciBIBI95oHYvLGx/a0KQKn1F+df6g04uLi0BM8H8jk+gaYIEurT
Qp5/RoYtKH0Otazo9kOpor016a7RGORLmNCr2ZVN98CAmDIlzM+w+0kX3rfS1ot2z2tczzC68v2v
ZkzbMG/zceGVIujj/tGRIPA0coFegz7+vwB1avjCdQdfYzzlMp45JWG50uanKccIApvqxN/W+s53
nzEFHPthcWHmgcZycbyhgknOkATm0uV0sq3R+q83TXcPNSCya9HuBEzacyOCwauDHqERe1lVQDHP
1RrRU87aZUZNCat+1htw4Hd87xDJD68NhY6GvclO2O9m6Go+7Go6dGBeRheOd+MGCJNvEnwEYQqU
3VftyrUrqZ2ahcusknI7MGsMMph2jaAcy3y636MtJuKWLsNEnOuaZBG/EGFIX1r2dOG6a4cNSZBR
jqjfaRqGAgdddW7dPnBgGtbRgBN9MuYLZh0dMMidHMwt+o1rx4jI3MZk1uaURznjzfAckMyP1T2J
01y4lP3jjXLRmxVGNbxdYaNqO9wKdwevvLIZlO+c8MGgzI+nUmfpkgTWxmlFfe2iaakeAExptZx/
OhrwNvYCwE4zChJDQeFwBeeG0akRqkSZO/m5stEFQa3zIGaei2sdHRfDOtNZ0P7SPJ0OXpIvMXfi
EHkwee6Y25rzDiTYnFy9OXM1Fcy09sxMoMLu3YqNjT0DZuBpQLACLAJkprE3Yi6orSlnFubFx1rA
X1Rm/ADODq+cMNYXjcfBZcaDlqqroKEoM270+RLQoQe6usIYi1fJZp6DSNDgoWXRZVXV4h7lzZ+8
tiG2+532zB4sfS3ZYkwXhzBvMWavpQJv9YlPHHRt+7Sfu+r8dv0cOJSBIT2hxZmA0xEIwKJ7OlcV
2rcxG8pR5ane8YwIIECF6MQ6kufEr2dSqlC06rApWGyYt/dyY1dvfUzp/XEOtC7zYx2y/xyR9Q+3
c1jDRW9t1slBx6PGcjIgpmhylydynTYx/153fffRkWjwkiTIftpf/hjJkK++xsEuQiUTryEBNjlw
dppbqX9EtsFaFxrUdVKwXeKitfEplaB+XzgDTiIyrWAZJLAealZJ3JQBf+cmkh6ncYZP8vl/gk+s
phJUcBNcMrc/JUFxsNhXLGxoim35BB5MFlNc5l+qMjh5IzHWKj39CEtGkA0BofoCRmhJPmfzO81a
zoGoyl3YX9un9kofZA5/w2n+7dOCHjabpCqzTwRT3Pzc7WBTRjpPjDrXH01RP62MLjlFb/80PZ/Y
Gz0QgQ2swwqkkFRg6dAVrJ3mrKowtN+a/+9azTtTst2OWUC076TdI57oWBBFPPHtECbsa5fCRf2I
Y//UgNW2UyR4niJ0Fvzv15ISMkpJCF8hEPN3YL0YnWq28EvPZOdWnK/dIZ86e7FpdukPrJ2aclQN
59LwDgGE5Wq7kCnhzciN4j6tqKCZPYaLSDA4dJtJ/P12Oq5AhA///fEkzbeR6U9jzBvsWkWed5FV
DOf3Khz+U+8p9rHT4plI4+MbxaxvsjQ0IwDCfq3Y1tQULoXJQz8IAgolPkLNo4cXpdDVyb3iT5M2
KyWV0ZEhpsJSeG6aStqS7XIXcKP2ilIKjX9wK1bsDM2JfLdvOlDuscjwzSEasgW4zFYwQVDPjfnw
CTWKhf2J4SkMoGoSRxLxzD5f03mp8PaWgROJhpuxxHV+DKpgzIzkBO0FpaKLfIcra2U9FOCT3ZKI
MiSVRrTMokctiUvv02n2ISx9R747bA0cf7lNGCjeEi8rE6WtqzyxtdI984wvJfxgrmmbhetQy2fh
Uhi/9NnPC55tkocZhRpEDKTLx2WV73iipfB8nsNI2RThwGChvK1vKFTVEFswV0G0wjs0KCx0FIKY
q1yn9c9gKded57oS/Ll+IxpsIR6fHU4vZ+x5sfAzDQQpDvX/zrurwekADgS4l3IksLpEuICLCchJ
iNz3yZAEPR+cn/LQTesmz6MefkkguNyK4x43AhpV1Ik6QYVdbqmBeM5rqx2981quqB5AmBqfhPgW
k4s0VrtX8hvceyAfidh4idyHB3LIh2o1LIraPIOuc9mSAVGrzAocg+ocO2xxIWx4GhNB1ds4sBNz
Aphu7Gq8MCFwQzjB3zucThSntFMZn1+l+6hzwLP/7Tto/olWlpnLrG7gMXwcD1EZbt2+vebfzpQU
FbiuN6wSk8RIvzuTOtMYjLDOBnVUiL222QdF444EAhpTFpzUXbx6IfuVaHjGqefTqQ9eyEzENfVt
Ls65UL461fzUydk4M+TlMY4+f/GtbgjzHnJuP4Vqju2RumyMQiB97j3Pus0CthhyjzewT950ldU1
os26EtPfNV6NgRJKCNE/Y6H01wQUerQiCXAod2LO6JIkYMGYS/AjjQZKXzo75oydw43m9PUWFNV1
MsRBgvo8MWrmmwaQ/GwsmnWMZX3XB1kojUQp/CvlTT0KJP6cpMouMHoyLi+8CZT08mpuGoCShFbf
6MbIR4A+nfwWbLxMn/9AwJzB8EuFhB/WONw7cBYfniw3/62hho3fHyfQpUNAnq/nTVHZ7/iLLjfl
Dc7/fsJMLwJc6GVWy1lNC3GYpsI2mgHIN1G2CZCcPd6+U++aw/3R3liIrw5P1CdmlSDPD60bIq3u
kNs63vIIWmcwb0u2pEu9FS91GmaCb/9sAZ5NuxAN69WzvufXy0pBvJUid79YZ0AAUkBBkCqQyfw6
mf8HqqWb5ZoqtYKCyeOimW7NhNVrYu5mz+cJXPTzceTn49njhWnazu71d7izoFsI8GTRikuuwzyT
dmj5myN7tPi/ZVMuanZi/HQVrxiF2p7Xza4mORs2UXLwzrEnu06Mj9V8Jj17ixCsz9CHMsHEoaeO
re9PpGSQpZie+czth+RfAAg7a4hheweuU8533+nVisA9fbaG9cQAV2mLCgWR+aPoinw5dmHKTmYK
uAz3AuVbCdRqfg5W5J4Wlv//224fBCMnVezeWE7gCA97Yg9dg6JHu96RnikgOEKTiCdwCkirjOvi
S1zKY/pgvLy8/2DdOB0THc4Gl5XT44i+bMoTirhYAr0q7BUMmJsCrYQv8mo5iJ3/8baaY6GsK8/4
Vqm37FgBpIQqBdT3JD21e9Ai+06/mqnebGNJ2tBRuIGnasn2WNkeFEKZIQMoIqNVhcQUjhp3eJGa
b/hx8zpK5HSKYX5ThVCnUaUcPAOJXmadpAX+ExD67yY+YEou3Kj9Ln+l5YsYgQM+qG8+KQeJy6l9
usmxGLYHT2uaUQa9dhsk8DArC+OKdxJq135se6v+jlgWqJ3M/48oienSpiXJgZ0f9szbeslyaiuR
NkgS7yw/xNZLZzdqA6LmlMgddoo0fvSDDH6Gm6mC8eRRkMY29kGBwigxuiasuHh8GEAr7Th6om9N
D4eSzS59WbL7vE5XgL4mficQXAmU0mXevET47bHEo/hGhgAeazBVyTD/dVWt/drDn10lzUHbOEk4
wdyo+FdDzKEidH/mrO8jXb1JbVlWlN+aTz8gKBRkw8RtaUWVvLTYv4pzOvfwo2MdG5pEVd1REkb6
U2HZZrDUzqkTNJNUJpFh3lmfeq1uD1Idot3N0SH98UhNksoT3IkKG/Y1QVMz3L++lDxl2RCSbK8c
onOYokStL/mQpnZtTdg3SwRrDKCk3u9bcHBaTefvmi2cc8nFtNZncRW9IO8+uXZJoI+wN1kPsV+n
kCmZnJWZiw/KmqQAnxFnYG+HmC+ki6qaO0cErXj1tefXTiFneyHo9TR/wdmYQ6W3YcJ7UIOD+7tK
FmYFjAxe9cIu/+53eRltcwx+KaPrzcpZlt0tVHipgjvT93QJv/czzzGGMHQ3ajEtaMozhekUkulQ
bpj81dfxL2S94MFNyp91rfW4OK1RpshDxgraUMUnTCndqw7wbRu/n8QKt2ErBIeRiCBJcjSU06TM
ZphV35/K5tOLMVe6uJtTeNrAwz/rvFORzoUFBf+0OddABEhk0SlIycpGToYhF2aJE+4+AYEUr9UR
QDvTp/Z/+e40l4jfSJD4DWM/Buo7b0ZbhuBycyN/878DFH7mxaty7XWi1tJ5IyKJhyUujxmSGJFP
ZjaMdV4WKat8PNMkC3dQnK0W9zpJkqmnimx4UNMx/7w9Z3U/UQOVjfRuycYb00lFZD4l6v5L9CJy
jQi2XgOyDQfcGG47CiVhlES9mI7sf5m/qFlhN690SOE555UCiMiirXF0EUOVwwDd14DNFRxsDpy5
3dPum1mknDhEByDM0z5RzwawrIZC/k7tghcC4v1Zjh8wbqXvZ+6rogLb1LsPEmklLhglOJgEIHfX
Ou5DveWhk5DhVUGa3LQ5eoK/waWvMGR9jp172z/fz9ZvT/iL0DbNc9j7AOtitYtwHfvndCzAQbd+
dgWyMCEteNAS4br8BlnzloY4xNYvl3JWxnXbTFpX2GxSUBuowBNNdux2VnJIG+C4jxnVo29V27Ia
AdC+xItxVtPyszBUPwn43pm9z+taMf0+BHXCZiUao3b12tH/44C05Z6/7K3ChVNCYz0ymOzDto+x
ZPh8HrNhs8ds6REXCVAFvRBJDcudGsNV09hDhw1teggm8SdQ4PH6moDFXML6vnZYKJsRSHPKOxHl
3MjAuK7rbjQfWm4Ew9E3H1fBFDBohu9HwlRHw6fSdsTqK/fC4wbUccFd+P/XTQ087t+lob6PfCXl
fmrAk0HSqvrhK6xaX4xRWE7XC5ImF8dDOJfxHa4TagobKBWm9Nx35aocYa9NsdY5OGcdfkDIIXes
1eIHA9Or8RynXRPGy4qMiP/56TSd660Auk01qhxKpfGVBfcB0aR7zuUok4edGSYaPQP7W91vKS4L
2qRDOCCxb9gerbaxKsCnglhKnJ5LrW/XoUCkkFzXH0ml2j8y/bZAndBa6vFICVaRCJaLq3vnkhk1
bIwqrTWE28UXMR/devsvfRMKbQyZdi2zH48LomFNV0LAqyYipNaNJ0al11zygo03n9kNOtSNPaj3
z0chur88wywLZzstaXhPuO6b+qFaqq8wTTQwSEADOgBJfw0/SxoGDxu7iE0FpHDaUCMb4sjqs7v7
wu6spOmx4uLqrTptA2tQ7/YwJYzbvu8rOuGfWi7KqvDuDZwDgZbVwvqqHLttjhteJjJ/ZFsS2ySK
kj94BP9D3Vzn2tgICnvNOO4upG+h7fmqQNnFSxhEquX6GXg7cAvz2B31swWQwyWP0HAsGvT/OmfR
mfJ6iNugi+v3UH+cv6L8pzSkCfxKZb6Egr5PgJtikMIWqNWA278mrGX78L5D1VqRuZVM50W0qaER
Nm7wXkb8cNaF/72IEeYQkky9GtDb4mh6EJHKciwD3JkxGs2C3BW6zQHaNgUnVqWUHICnx79E0m+e
Y1jeDZIsigWSkdhc49rlnkhJvYU8i9omIcqgUIcB55DXK7Ufq5BPuHEb4TCVJ2iHKyN05DLgB0ks
Umaqod9L2YSaLAQUdX6uS56VDWtKqqWM/TVX3GD8oA1TSXr2C8/cqZtL63ZytgFClNG88Y13NkNS
niLZNIbdrpR5/umPLsblH3CXn+VtHHj+bGjWfiexlZ6yWtUXI1OjTSpshyILGYVtNRFiqt/S0691
Xazx/B0hYS7bOZLhSp1R4QPjhuBRT1UGQw3PBvNiw5EApmDrv1+Pd5J7ygjeMN9ikL74D8YJjBrh
ZqpfbPbMBZa2Fb8hiQpUzLwLfun3KzuPtLt8Q3+59yIe2tkV2HLKAjj9ZnvOLbmNslxcZMUg5T23
R3g2mnAoevwCVCrT2vFwLRtnnp2RcUaIjurXiO7XlKoM+aVmxGkiC87nxXJ18VtFJ+maVwNzpotO
tvOQHvI2KhZSl8igmNFnSzjJ7++DN8lFMRu/0qU2lSCPngBq2K9WjCsUjySMScAJS3S+GGSz2Cce
ARL4EYFuJuCzfPExlsx/zqak+tnll7LxTSfPXnCTRanFlM/UpQ1YP/aMjEx5u04TUxj1r0NGfKp9
kZ3hkcykhbGmoQUOaywwqXIlv2jaeLvJMxOfH73czb0jQl89MDxYNJoQA+tuP3isVzdzkUX/cw8T
ez6SSaw3NeQcGqCvEVR+Gy1ofQgGjk0RxQDCFgaqTmMmg6FwWjHcAhPCV2Ovyl/qTymd8+35xTcW
VUphsH4qf7nuF7Zhm6uM6u40cQRRTJWSyJZ5Wl0PhOTgZZq49HW3JDXxRBumqRsEYgw1oevjUZlj
nVk2CaiySTULLL2HRsXGt3e3wg6HeJ47jcRHTmMAT3oa35sOb3/qe2VATvQYagVk1dDEXsV8ZG6Q
9duGntCeOHBP3XEudKytzYXXLbypdr4FKzEeyPs0IGOn7nboWD1QTBBAHMpIdpML3sX2l9ETgBSe
/2dxTLNFn9ZWqKFSwWeNFmAUHLW5WNLArMy9uXASmB48nEXIbA/VPC3ZzJgEA8HHsnZum/U8UZdm
RaLRRddvsuCzxzo4piaflob+gFfx1XpFWjosm5kknV5aZYZoCcmvups5p5W97OHx9AxA6BebemL0
UCNjAv8SSOD3iLBf5QTAYkHBwHHQi5WTq+Vo6qysE2ymkWBNAKYFqOsyyKBaSB+i/KXufTb8+ftE
Fg9mRJZc08gHO75Yysbx03+cCt778x0X5J3MDHRDVXr898ggG5BPLO0UtQ5l4yPyRCw4Mty+j0Qy
ZrQI8pEAVmar4w8O8Hvm5iidNgCIjd5LgW5bhvHxeOqiMqSkYUP9WHCeJDBeCHO2HgM+VcmhNKCL
jC6A8xsK2KQHdgUgDoQOlRlE5G+A/ObECQyjm3Hd+6ObDi85AnoAGNIcCj2b8QU6Z2A+Mv7mZmU0
LYa15+zvVkJY83XHLOVQOTeTuvUQAooySmWfJr9QcrOVpps+HD8Pvidhyp9HPRiyE4GcSSGVVaik
djavoNRN8qYoGHoYBruxXelaKTnykBpislzpW8x5330tEVbPKcMxuXuVf2tJKyGpIB9bhkHB+yzd
hy3OUs/38XQMCWuPomJ/ecPx+KhHWiW28boKiBUHhbFt8bnSu+ra5QnP0NyF1cmmlT/uN3vOnVQf
jRTa09ivna6gieuCUxmHZt9bjABvzxZ2Fig74sSY3U3Ygr9kxUhYoghrc2qgez6WuknHMdQ/5AKq
ijWh6GoP46Z6o3eI8yhaU1nzXiXrp7EuDilB+FNXqIAQ/T9pAJqgQava7KIJXiqlkbk86VpGKDoB
sV5FAakkfTGCAomsUHg3t4BWnznE2gHwlChY1XUls94OSmCWMoAlIwTbZRq87MzeiePLwC7cfAZD
v3wK7vNGYB28v2FTjxRi5aI4YW/eCY6tTY/g8FprL+V6aglAVBWwwEniwpYLCrcbJwW81ugEaTOP
RCok7Nle5+sf3Artyqn7aZXkciLXACaZiFTsNgDuzUgjTQ+lVLIWdMN0n//WS+d/r29qCYPGBFvW
qSboJ5KiKhJoi6bLSa2DJla/kW1C5tg+ExRbHWzOnrb1agnE/MORQupQ5IwSaA+D4wJI8M8rp8hD
whOZEY4WMAJ2EmIl6mvGCa9LeRgyLzqxrnUuv+egxqvFYs/zRKK35iyqIRFNCx27hAgHPVeYt3MO
FqRpY3Lx6+kJ33hqXKvSOnlay30iYnYxsoH8O+2fKhhYYoEctCmpLU/t+TTbNe87TINVzmifQTcA
XZfuSmrFpjnuOzeAfobeWIOf5KWrSTJMw/yurGoG+OVcPj00X1g1rqw5qwywKjm2FW24pGVsVAas
e8JMbj3Y5grQylqQ9xSYduG4NRwjLbDnwSFi1WgWxQG5WEMQY9FcIuTrnVJx4oZkufQzqdRJdIat
/SmRmHKWlaSG1amx0u/3txm7c+aewSGFrGhKnZrjD3FVgjGWdzv4efGA2H/ueKZBS5aB5DzZ4gg0
tz7HKMIX27uQc55JVVysqoAHN5q0fTh13HODHCd6abXb4J/0uAFG5Q5H01br61S3udBvCdk3Z/PG
qspKbcVK1aOR6U7rPEmbBVsUedfFITYLYJiOikNxd8iM6B7V3rzgDzbRfNUTVc00A9ETa6Rzzot2
pTgYnrQ7J0pR6tb23YXuT3dVEaYA/q4I1fZFMDRacU3Z5ox13vd6wtCYAYLSFwMaHmNNatkGi8t9
5SdKETt47ZSdNfIlmJMJPrBpdtcPRwroboh0RDMbvuS59TG7sNj/mn2C9ZmoEhraXSmlqCNJ6yfa
DrWbY8T5o6Pnu+tRilycQ52pG0NeNekjLKSTktPWFdjDbcTixqQ1rTZh7ddDWkDF/Pm+9FSXfSKo
CmuKwKsI9MsjOAVt7Mm9zmRdFJCkO0xBF9//enAWmoIKI7ASWhjhE7X/7L42f3FG7CZwH1YQWLLd
fn0SbmjM6XeZvldWPVP/Tl3fglKBDbKu0eIPO7O5wJFz7odyKY2uVlLcsPkQ18c9Y+bCU5WvHqvc
OQuvw4GnayJ9y5iQwQmoXu/icVTiUJP068Wxy/67NqMZi7XIm3AsEGdaadm3U1XLY8uWxhxsCdFr
tdJvq2u7UVvFisWUYs98C4PLCzdAISAdhMkmR/ahGsr4wRHiWivcCUKz7SqUBORuz7g6kEmpLmvo
BV8Wv9HhS+SlacHkb4UCXZlUSw+K6u7T10KD0fdWrvpz9KHQ/HpsmaPBDANDPtLavU1mN3FFa5Q0
eqXDML/XFlswaGPhwv97qaoZWsM/rTxT7T5FPkpzaUtTsq3FK9YpNxoEjNnma5pxTzFb0eTxgmN0
/2fKUrnBRT3frQVh6l6YNKbe2+vcjw0p57sx1uh2dwAJQImWmHvhYf4M77P67AdE9gaTo17hcyz7
hQTIvYdpSw6Had98h8NNHhQhkH05j7iWnN19N2eYZg6XcnkY29B+9S0aUpSZ0xuvvfjmY80kpcqc
5pPq95q0qh+1UfbZY5TS6ZzoLEaWPhBrqkZ7gr3A8QGiBYiOJyMlg1vM2TtETko/NRVeD/JuTFTw
HsUH0nd2sB4udsBItYMfp3ZIrvZiVowmqE2gg2qiJaSL5HuqzK3FFmuCIUhlQDUMuC2oCEDYcHza
GGwn9PGg+wJUNrh3KwoDlBWgZwWHoxpUVKfqRfKzgxDVXnYGDjBXO9yFgMZYJBDydc3XaHMDLnjc
6ZrdERo9sOlngkB5xCqra7CvQdkUAkOJpY0oTo0owsNeYSJ/MQtKKTraB8bcZKkpUsVXAYiRpFej
0GQG83mXVtBSHpt5LG7GIYb1wDdDWh8clVzq2/TpwEjbXySton4VOQ8l9JeUrZA1mU+u29ACoVrM
jUceb2plDObBatyUPW6QPVo3PvOcqTFI2iyPZ/bsxeykljrpMisPzUsnhPPHoe9meJDJT7LPxwuq
GBghAXrfnb5BpQpHEJ3PIL6J2WXVZbL5L3Pa763ILB/8Ne5/eRoiO5ANUspjR/Gork0FQQLnFzs5
l7UrKyzZLAdqx2o6I/68gpoSIojcDPKtHrTqLmxY2hp3iHQdQJqXkSnjwAC+xTjGmpINKlwU3sYI
0IuGVH4l6TN/BPFbvXdHUz+9CLCtJCLfnTcaZkoOzbXiqRJW3FSQOunlL4UwtPhU3n5sjDv7Ykr1
FIT/HWpCHouAW1DI7LG2zjsMW+jU8EXlDp66GvZEiaw2+gnzd6iLDJ3gmYTmMDdokZFc65xn1vxJ
dsa/yNMSsVv7d1sH36pq35VRCFJd8TLR2YsVyjvQU0ztuYQJhEug++75mcqnynEKRGzlvB3mubk/
Z5gBKPMDHq4ZJ/fIP07AoLI/rMRthbj13Wltb4TdughOeD3XjeUkmgmPuvkWz4zNKBRYhFNvPxg3
M4mWJJvS3dU4pJ3N4womAOGVU44b097kGj38O7x3ZWZEu0McCmqrBhQwq5TAlBTFoUFHOYUEccOr
wqw4/LwnBjdR1mELvrdmXf8WX8vRHooa4WQQnRkXwDDFBHhBJL1/6tFcQHe5OW5EzeBQFWWHYYPn
RbMftBUXP+LLs7Si8AvBp/8Q14Cl4DhYQnyswJA0jrGJFivFnmgA3O4rzD25cps3+wyfLFSMyVoX
J9OvHf31Yqq0p/BCJVt+gvqiizMTzOtKSyyyMhlMjvh8lF/9qUvjx90p15UQQSDkqxeQmlmSULX6
smSyCymNi4qaMAes3ZYbjDl4X/YmAgJR99blzGLU68zu7RO+JQTG5nzQGkMB+0/8bSJ0LtWs4Shr
FzIhBZKgzRDH/CHLdfk/V85JBSURBGgjJFWL1eoJTH8c6y3cMIY1PrdOXsrkoQCRngevOFv2zDLh
T746ZQpc2PPMXQLkj/fhBxnymQ37xIu9hL4HobUhoIuH61g9URh4Ymjz1E3GlRK1oWHe++H2BLMq
E0BJ7ULwD/JyuSUcQ/Yvb07BXEQ5tX1DmL4T4Gha27idMepF86Pt5Qac0XMpZ4Ct7Rpi8VUyailt
fc5sx5OH3NnZdRR4s/8abOHc3NvNcvAgoZp3milqRT3VvZvS9FO2d9bUTx3vbmG6mZ64s7wEGnc6
yk1O/ODvZl8DnGkNHh/t6Lnq0Dgxyi/lxYsnFVV8LLFogBiZETQe31ekTFXACIfJQDRdXll9eJD4
KQGqMijF0uLeh7frRZAEKsdZsqotWHTIsDD+ikjxkzmGmqZZdY7/5QH6gQnLZQhcp7gLJNTSxbG6
hz7Mro1dqNunolkeQGOIj2LcgtRJtd9pJfXGKzPWFcGjCNy4AXOZ1ttj88bR58WjZWvlwJItbL2J
LfB63DOB4IBj3TQTtjuKiKIWsACERNRjNW5bEHZLaXGV3Ny3TG6jkkWHtu4NxVee/AL3HCpM3Ahm
t/96hbdSCXQE/QP6do7RVVbP2VB2/edUnDqn6vkzQNZ5Ppk0urjL6Q17/rNYeKb5YRQSKK6WhL7n
En9Ols5Nr/DIzCHoqmLMb/+yMy4Gas15vbpp1rrbDLtGavUcFHfGVFED+cfbrqCniAg+UqqogM5/
93CUBxtIKG7qThxAi7qOLHjqGfcmm86sqVRkT2RliT0wP6aNOQR//mcXZb530IDqSBQD3FG+CkEq
7sEz2uHj90BnBe1dARl0+iusIPLLktwLctAA1IGn3FfUfpfhxFSJBruMNRKBsaRePjDJxKvD95wM
HqLUNKBggn2TYMD77DZMoOinpM9PqzPjplJu002H6EeKI9SRSRbXiZmbnKuD+MbpW90XtXIz9jAo
5YfHaZBR9tW+WBBe0hgAV44TJ5C7f1rpJ+L//oZSvuQEjrucjorUPm9/5mkbKNcXsKk8EvNlk4Lh
KyQ85AkzikDO+YKRCexk3WD9llLFMZSP970JqVrIQrSjFp68hRj2M0z2IjN3SaNorpPL6bjEBgwl
RWweMfhPpxMOauNVUVgt0jofWgviyiq47sl2PhIAEJGlcGlW6AptwFng5sgalfWPePvJzWdqqQee
tL9NXU8L4t7GKclZxdOnfpmarYTEkpNz9koR3QNvjDgwuKpm+U9JpZKsNQv3uFFeE6OC9GZ4ZXDt
Y7gnys6wKsDBFd45Jf35UhgW3En51Orovf3QkBVzeHbE0GYI2R49K4NoB/sJ/S6Be3bh7VDxnsU6
ku3tqzoQGHlhRURAYkof5s3MSw12Lua1bWpR6HoXvc/jC9Jy5YH4vfK5s+FdcyMgBDY6uaM7Gkwv
67V2gVax7JJePYtt77AUXZAzOykYWiSRovRqulQsE39EoF9vmpSyZ1RLO732n5mRcgbBZy9sCJHD
43f63h13nz/2sq/2yjeU4CKTeaa+OwkA9TTCmRb6uzUTD77dsmAcbVqGqDY+w6VixIuYYA8tpNSY
cUAMRo8EtYJ2TUMrcj4Lieuv4LXstWOIZmRWXlRme6VmZ3udfhL7+S72fdy75M1LK7hY6BF9icKu
+Ep5HtdPx4nb76LcONX4xp4erzxEjfwG/+aA4Us6m/+pT68SkUntDZykHU95uxiZ2bu3knNVtrx2
KLUwfMTkvjvjLfDxeFTMU6hStxJXfqdj5RJUJfldk9yKP/o+V12VFsVXK+lKOV0rwLRVgDroWbZe
179PwAXy9fNvSjmMiBZJJyxrat6W5ho9fo/l2wKED8E0AyK7aRrHV5FnJgEA863sK38P42WYTg2x
xoqn1H7Re5XNoFRCgLEPdFXqM4yJjT4CmSHg3RtlDwyRAxJEH0TsvbZT23CcFPO/ULo6iAFjES4M
tuRf+ZTZikD+JPtGv+Wb8//czECc8pyKk115Vp51lHtAP0C6obd0q1ORWNVhzwhKV6IrhjAr6Md8
6Zab3HzuIdhWcCNvbdRq9OnCtzxQn6RAplxLTI54jBiBK2dHPBdLsve8r45mIutMG3rm+ydhGZEi
jMWAfAp5vKxiR+vqOds4/h7BBv0wLNH6jPF0YAcyrJ4riiep5ZKNzJUoj2yJZxZdwjumxrYbBhm8
qrqsvra7ynblf1bqe4vr8/IbCj5zw4vORH3eC5AmtGiNCht9UeqsUVZ1pqKA7SudjlMZbSnc5bqs
TYsqW3MJuEbmKO+89IWra6Eh1m0Vy/1HKmclF9mK6HwqyNOCPCipyktmfawax9nWsS+62ZjNtxB9
X8cHz0y46169XiQqILSOeq2c8Wkfr2KzHCzop6r2djNjDQa3gXNhKXuFCSPLpaGhEEB0fyu0rfw6
PNx9b/EWGly6IvaKIqVjP7D0TwMPT7O8FI0/b+u5ryTyPcBMw8Sx/Ur+Kq1mkIG5anyryJj9yiYB
JVDXP7w44uPfbouLkzCeBmcnLqYcQVLSW40BegTm+izyD7BfSjGdwJZTiaFJH9U756z1JaoX/oHD
966zyp5UKLSncZpZtfeDj7nAjjqzE7hsmcOQQ6h5DeJCDFehi8qz4sKAfkeVT6cH8jaLmVALErii
NrIZL5VuIQNLKqrQOtXZ+Jo/wKdPJldF40zfxnwQhbuZQ8Q7je/NR1i3gnqtYtWTGTkAK9vZS56O
6srfxfIU2QP0ojN0Ogj2DJjisA0NFsE/eqi8js3b/UvdqCpFSC1EAJWd4pPtanY7MqMO8dAu2kJd
Qz30ub3xJHLMqZRStzo1mO9LblB0uy/F6zf30GUlIQEL9xkyF8JvQfjuTnNWlxiDbcPsK15b9B75
sBq6tXqVg5Di+Fm2bf3iYENbejTJPwft6AYx1Hmxva7UawfFedfAWETj8Yfd81JdfnARsra38Pxk
+Pq7aTs3UmYUQEo8L0SdB+6xUsOVRM8qmEu4ewfpu4oKq8yPduPnHdPrjZTJ9m8BdB0vz/xmYZIu
8/pncNQ8TLtMPFufo0l/FJrIFuCLr2Tuy+RlTxZ9ENB76POkad1HDn7RxPODGO+xzEncyixP1Xpo
B48L3XB49wKiQKYiSTk93C3wSV00H/HzlWGo22aYNHowlkuYyI2o9ktqBR9woF0RssfqQ6ZEfdXs
41dGa8pA2vqusWa2FsVTL97rEiV2+5pehnemfCAHzkxNYlxUFh98axb55PDBxGfKYlvLcsr6MZ8+
4sItHdESgw6GJp9mAMdqzKVb2Q7msnt976cG4ae48/mGO23MRLCYxP7pcX+M7rdRbfMiOw6qqsvH
ezYOTSAKeG4DRIJ1ssIhuQq7ETk5WicDl8iA2/xBMgj9HHYkYCmxGLZlwCAkcPxUGdbKdHTGCQPC
wAnMv7WzawWYim5n0lbY+snEgHr+IlKW9Xw9GTwNzhwOctyRSFqdyXcF/R2x/lrYt1nKZ6h6ELZs
qTh/ryMBV1iXXSPV04EehSZVQfzb2etz5VCNBZupNrrEiR6zWTlxcy0LnOoa2rpFRz3afpkkm78v
zYw4c7IOQcbsSTHyhwmJGAvZpmlJc4VS+ezLeQd2K1uB6KFLMjUAUwQ2sZ8AVcM165qrBFVCz4NF
7k/r+8J/QzKfUWNNxXxPYGzaJPwLPyspul5WIzTArCSyarsws2nDUNRbw6vKvptni4TT6HU0Ry83
KR9WKTlvuWuw4o+uASGbt2UnQoxvqHSPAmym7NeE1UeyVV/6G/IQyjc0JopZMYI9cbP4er1exwgE
lCWY384Sro1+mG6aMTwzqw6ertKMCessobMLwGH+2pLgXonSo+ZpQtPhjY4LfT5yhUjv1YoI29kG
T/R5mKbkmaF067mSSHMUzL/H9lnJYMH/tpejaJ5zZ88t6ZHn/N/UMqiUpbhVf2+QRajoXKIirjij
Mi3ZSNHHBET447t6WFAEHPHfw2VfaAhiy3S6XTTPD+XmgSS82EKbh2yrsKYTBxvU+m2rqJ3bo2vO
FRzvrp8gXSWkTRAk2B7GSjgvTIYTkdzEPI17Bzjur7VZVWTZY2sIlWJicB1ZoPRf/mGqFTs+jMOx
TYOASUtjjZCri1AaiFx9yQyDBu7asYr6vX0HvSvru4FlYGoY4QecxUJGPLiYmBkRUG9xi8y4EKbs
uKfFmbXW1/FZz9XjqYglo9SMkgscNKqwBgLsi12vhzKy5T2EK54eBY9ZkTBT9IO5vzX95GmKVCl3
Vxnj8dRPbEuDn3F+gzlqGiUyfj0MK4d6VjnoldQD6AMTEMqso/+Laudj95jU61bwQDPnFJl1wH5n
y4t3kjkCleR1vWrgobesuL8Euld1e9bLHA+ViChnNpZp8PbsWw0AY7JROgNde9tUhpFcrhpK6fZ6
Ow/zq4Z5pMz6B9kOzh4ME+2RyCyADxHoE+8GDJBAHUwFX66/qQ3TZbhjuszb79YNYXa4RmGB0yWb
qDNsP3tmK94NH+Fi74a23R6q2a2uWc+u+IHA6ESslIDL9BDNQu0UKFS5xsZ91WL4SAOwQvu43ThF
AyjCkcGvS24W/UeLmkLjNXGBPgUSiZmnJSu9/mng6myyahmVGSVgG62dCtBYBypARfi5AEcY8YTL
3zwKTZzJyYS7TXzUACwob+yKevFOpuaxtGgeYwMlk+ftDh0x+d5JKrBIB7gPTRG0hMYe3yI29+f1
RbwUTUBr4khGRc3gofDpeOpvBiLnCzJJhc50yA06lhp68AFDUBfEgQq4mBznm38QUfrPdkEL1duO
G5oizGRhekL/zajfqaV4soowzyEG2lkPaf9Y6X3FBQqKkAV0O0etr+0OKWjTtdANnNpXwkEkeEtk
LfNOXoR6r2DerAbwYq5atbH1iyAY86Af3hSDMocaI7bwhLvWZm7n4g7MBhXqrJ38M47JAvxMq0NB
XVaPFz+UDD4foxx3AjSf9Sx5dhf9EWviKNRMOpWadgqEpbd32mSKgEdNcrPUxeMEsfvYSvsneeJV
CcBUqLzr/jW8G1loJ/lpdkjO+vqkly+M8OdzZp3q81LtIA9nOEIXEzJIc4oeFZCq23czQM/87Vtl
Kd/McCihGV5LMOTBKIG3J+hMRjKdn/zV9wvvQch+qApPgYYeQG0JYa5gQLb9/Pvcu8IptizZbgP4
+c5+xhEqiFvrc38ZSmJSAitzRZeAl9yslzS/exJhyDqfYfX8sGscFqKEGLlsTLS8ypi/GTyAbuqt
9jQ4gnFHv4TpZoDSIVqJJ2NSON6tnrTSS8D1Y31v+Wh9SuRECwqOCWv8+YSP1LycaSbBH1ePfnSg
ZwfPKMLRT+1jNfcq1o6oDrxe+i+b8g5YxBQxJmG6Z3Kvze0mi9QQiVsmx7ZhnlUlLAqWGEK8oHAI
66HQITWNbi58pZxziXnu7xqLed0IySluI4qZh3OCXCkZ9a7hixQX6z5BZI78Ch4ZJbvQz/oXSrJC
N1qaPHBu9IWCIymXX1BGhfojGA+fJZNJ9PmCV+YvV0u47Zqf/gZljnMq9Qc4OlGo1Rn+VNUrZhGG
PeBPQn8eT43CCWxptPY+wlRiNe5e+58056qFfjX4FfB/ZEYvIGBAh837nwoJ6jn7yS1RNG09fZI3
P/ldonH0hab6a9JI6aRORkWqjwxggvwrVaHMWy0t1psQHCGmd23by2aJ7FBmPd38dZlXSh4Qwb7v
IQRMvp/kRg2Ze3IcHCdVdAtTI49VZc9UEEb6o0nUAjW1rxh9rGTu1wE9W4d07CoP93dNBjXv/1hF
aiKjkGnnMsE4zdYWcQNfBt1Xiy9vV+9yXMH+Dd18eRJslD+CI85g6hFQ30/JJ/ypEbCBKr/V0e71
d8bsLP+sCr25qojELTP337OpLxwYYXbnQ/n9B8X/KrS0bSYBuonDSPX+tAqG2WlvS70ZGu2R2w57
hPfxRIr7r4bzQV5DiBjyG/mATzeaRQtA3cRxohsqGLjVYloqMw+2cKGyNx4wk7r18bvAJG7wBEaI
Qorp38Gi9cymKNILSGtkCMaL/mQokyEIHarUtZD++BQrNy5yyvAuftVjCY9RiIDes7zNrNpiTceO
tuMqW5smDlhwPnYJmCnIAMMp1t0P+i6vcfnkER9nqsMcOV2wfOZVHLQMTufrZ+u+l1km1UPQMx7Z
G6v0xSDb7u8F112tQzimUxmLdeywPPJhZdt2Ai96zAnf8jawfx2EHpeI/tnelPYZMPY+EQmxICFl
zsLpxdFq63s0R7oHo6xwc7u66vDSL/SidyPpdkLVcjChHCn/eMZQ/MiBIBd1eBgW5kuEkZoarikF
3Om1Yu5QkuJtTYB9eiu9+nv5q2O6G/ZU5XmZ6kVun36ia423z3XrRx0OKQXwLhTtMIm1sidHEyC5
drtOh/r/oJxfSwiTY+Y3dhPYwpZRAXZbas2uGCYMzsmhV+SaBsHKdr4SWRoibNODzjetshSLdkt+
urxHBKlwCNRK0Yin/2lUCfEyG69dSXTRNkuG1DV+gRzI+MI9j6gfaoUbKxyflZYlqmTNUm+a/xJu
N6/iBrlvLAcljC98qOVeHEETukddcfqXN5NgTuXpvSbo5TD7j0txBC+UjGnWvMsAbYxynKRoN8ZE
KPhQomd/bOjMHyVYC8MCM6S8Q0QBGTTKXCCQMiKvQmcqANQcl+viyiBpgcgBWMwe8YyRMHJOaH2/
D2u/bsA7ZY/xT5Cm6V/6rfhRTkMRHJObnj866jewSL4m0vdqlL2+bzWMOVqtnwkc1A/MzQnq5uTQ
HlbebgylQjxFsNc66Cl6nquBcL7x16/t5eEuAVTln/npGAaS8TdkQdYGuA08X5DqFCRRqoYAcjGH
izPDw92IRnelAlhRB9BYDOQcSueAXzFuXhYRG+ySHfnr3WI4LcQtBEjFym4326O5Ke5sXdI98M5p
As8q9h75yl6WhOjL3AgCMmZ44KTGG28N8nBFelcbcRrDjaE2fnivfkLRoiglQdxWBqozZnZHLAkJ
ILpS6v63LTh0JTN5FV+wM6GfzQ+m6zp7PO36hu7L8fy1xxpbopkWrchH4UkDMrodzwIR+XfUVm69
ehR+zqMBBCYTKAApzfjH7HEcJzQ1VazRhSKllXJOMFLhjHn5FUXd4o9dxzkV0DaLrSucQFVtAMvl
9e3WtxgtTyGK57HiUBoKzCr5yAJz0DNgCAmZiAX0gK57t40DT32vC5sdcP4UNodVu7FvINGGn6Tr
g79RqKjj9PKRc4FwMSgKEWFH4tHxurgVyU35x9i8VInkl3VHP0M6KDI1lwxXhSvURYT+dnC6Fi6X
PDk+GBNEVlOsBsou5O2nRrx5CyVeMe5FAEBuJqibrR6NLfpFSfDTk2be9ckJGWG3mvXy5i31hPmH
dkcWn5LgkwyXpx0DmP45RxZaDTT4Zh8dfivzsAMBlKrDspFHoHUPEe/obyU+qzWK0iQ046IKsMwG
eiRs2lB/d3iPxGKNQ1LAOj/bCVcJbhheqfnaSuYHt+VhNnkUK9sQM/DyCOAjJ2R47ISvBjIypuuA
JW9pXdweEXd0N0PLQWj6XQe1L0vYUfl4uxo4MEQetsfATl1KrVo30SXc1pqAJKttkDtjCDnxioPE
y8yv1uK74OQr0Us/+tBrAGW3eddwu256tf1oMpWGuLTEvQCtC28c16VuilIfF2XwmJQOYP/3XSRu
FhCKfyk/8NlEQ+n2IoK6a+tWepKLjFjdYeXhBuody1fchSD09tx7iIfUu9D06b/ygDwXDakv3V+E
8SVcFa5oSMKxyslF0ylIg9wdxt3k9Q6Sj39cEloNMAXm3l3KxsQ8yh60C5GFhX20LPWWM/hPB3r4
+anTGonohOlt0AbaRQMR5cJmDKQf7UK/bJ+x7QCXWaCf69Fqq0DN6PHwvvbfgoxO+4JKBIS/d+L7
MNr3YVDnLcHVGpBqTPGF7W8PoWuXDoKyINphyVzX5PGJk3NPCjNPo4/u5XbdcdTtO1ktD9dDH8Xz
zQFUnlTZGQTnCsaDQXPIJ52NxNfnlmHo8OCWvK4mLp1Jwk/Ad4UoxdtV5+YWZ1WqHNy0JzVGtzCY
MeDMDCj9N2mOw2IFTAzO6+CenuylqyYoKiZxY4vhzhEU2gG8otCUt4jBToJDEzV/NbE6Lld+jK3X
BaSJ/DB4hi/b8EDZKCktPYy+O6BdmVAjEkqjHpFvBkcmQxs80zHuuIoG3eTBltfycPARll8vXG8m
c3VazWwyyHv6UYZDXSpDz/DknjRI986k3n5NUsCUFR1TZ1O9wHRK+u7JIQZFYxfhhbejPOvtBI8H
xwJv1/iu0zHEK4IdeMkyiVG8BoEnAOUdSPk5IsCKv35kxO10J99aliYf2+xEcCJ+GpExKFvf2USj
qYcf10mNjNMFO7g7p6EfO4LbGwXbF6BPFq+LpkSzCPSeRrKLjPHcur9b4NhdamHDB5yIlGKtwD9s
/Hz4zxbdL1W7O+krCBbOfb87UrecBhfQQAXVc82PvYFE9h4p+pRI+sW/J+81GOrknl0sTTuJOars
9dC2PQIHSGo8oTPVB20WDmeTEzX1fUb++BWT9b3z4FqRI6V55FjRg+lVsZx8LfHsOSIgpqU6DbEs
cBjSOifB4nau/OVs9ckfeTVzC/eWB23ahph/vyPF3MLvrre2XNdqd16msEsbeAdJiZb7Tj64slCx
3AuTjXnnT2ejmBNMwdsLo2K0tLGUtKhbucDPm7nIHN9nIeqo1dbWN+S55Rw3I/cer2XMVCUjJWDm
yq8XDxeHT6ixqO48ELaJ26jQHisUZqoxkJs7aKCQdtbS2UDHbCY4dnUjnmc5q+dixhpezkoHq4ic
ezlZMVwRh5853t0y+ujHWnDxNeQU1K+MQTpOXjB15ydLD81gAV7GHbaNoA0NCIDn1WAS2DPhqQuq
dU106opDEwmbXPPhc6P0Orq12tUE+WimqNlysHWNAsO4DLf0VL2nXh+xK95ge8YMYnIxNnBtMB3T
vggkM2VBPtg5s1wfSM0y2nA2yYByIlIat4FnsW4ATXLyasfqDAes4vT8O1f7O5abGmIG+ckV91mY
Pvfhci+MEMmhSLHNeGuExh2CxUy90dU0UdKhS7a+RVBq6TkveXTlVBuoOx0kmhPOkApMfh4KVeOK
ms+v6qpXoNbrwQRL5RlNa+/4NEU8flP4+an+G4nbZ70Y6vYurjVGosXfl8JIYyl7QVl921S/BxBF
oxCz1/P0B3oL9cAjSaVj8CPS4OUtYDgxQ6tvFs8BPhzLhHZsHU0RBnqFx4GsSM0ZMuj5eYfLKmN8
ZsCN43Kqo0f1HyMiHI3t5zXlLPFV5gPqfHRKvgkkfY4jF1PiYRYeZzApQMh0mqp7kLI87fRctz/b
yAV+g84X8GMvGC2L+cxAJxg6y10ndnrUD+qM5ateF+QzwYzrG0DrJ2N/gv7mh8e1DmByC0siu7a3
1SawxoASjYYLoMIu8cyhj/oztpIFxE7k881NVOLptFro3I0j9wVrAcMs2Sh4kIYE3F6vgJ+R6Bxr
9gxjizkQzgghWabz1WkzOej5VqjhZK4HW742djtys+qHaPo9cXhuw/eVzD+SdTHZRRpgbcZq+TGU
1pmTQvmpvWnkZX0B9Ocv4Z9Sc3I5PjeVSE2ex3iX/ks5PQY5C/IqSdKkZLmMMlsrhufquvbYuHI8
RJ9BgoZpzJZ2EW5GQq9FnNQQANgifS1nRzWRRGHyqCUzZpLuNYGVs3lDoHg/582dz05DGY5dmxtZ
BZNdoAFStflWagkRP3+PgxdCpk8q5ha3410F0r1MuXGvkjIQ2ZSLXPWY4ty3rBOLqK1C48PX/agw
p3w99D0tBpWoVR8vqGaB0HnyPULTRpV9gZELAV6LeHBUu2UM/lHzEL2z9di/ig/ny56ki0WjEtnM
j6vIGxVFf4Uisv2iMVoaZFyefizmu5x8FXxu94c3BtL0i45Y4+b4E0w2TaeQUaUHjVwZKQSj+zUB
KL9E3bsgqaCb+/WFLgxKPi5OqkNcnd7tXlOFb/Cr34WS5PiX4i1Q3M9BuDxixqFqHpIH1fQCDP7I
MPznk6vwhqic7wsD2LcZqwmE4CjnfAP+gv/ra2+uFrLa59plaN27+jbFleDvVmWnD2FaJFSM6V+V
GXA5oZ9IUP8XIhaHFlbGb6LZ1/BcAmVpLi8x76kzeR4o81P17hWRJtTijWZC0al9GWU7dYC8syWj
02o4kdIFFKaHyqRObRQnzLtdg/sNW+QyE11JXGVKi9YbS0KG9eeavylIyVdpt322WTlI5i10DcsT
DjdY5acTkaBYNumAd2nv8g70NsONjV1n36bpEgnTQoW3WNldVibZAR+FkA1zM/VyTzVOYR585Yhk
Z1BBFtkAhu0wVrjrHGTQ2OM+3IdwOGzWWQlBD5X4AQo8OUmrMCgX+st2/i1t4hSBDxcOTbp0VtSZ
BrJYQyNh98+BgeUWg3qcmFRfpRnQLaX230A+sDN29spBAczcyvip3+m44m+zKj1i4PMCNevjXVKi
sCmPNnvtZ3/fEzIH8vWK1uagWRIVyiYJpinvxPWhz+ymPuXWy1juNL7McKc9jTuAy+wgqnurFS/e
lqUKFW3PsA6uBlmHYuVZEuxugFX9p5izbFav5z6nxRSfb6KFzrfeQ/Uhx4jJrnF++XmSuh7lwupR
8plEexPci09A87Qd0t2jhuyIWYGfJ8TWtBfzt576PcS7nWGDPGKIlAmIVPOwaTXHRW9cbqB3fL6K
RwumLnQ9DsKpddDOVJVzmPkgraQm0V2cQHzV2ok9dWzvGsav6vmnfB7xhEUrv9GBFIUjokMudotP
xMr4z6HtEELy51crhH8Ns55kQVsa0YZIHMHm09e6hXA2GNLhngokJn3F86GXWNUjT44qp//jsym3
OBRjE6nNweBU2V8Pd3hkG5KU5LJC3iai5yXelG6d4HEHFgpBeL4NGM3lcteLma5GJttSpYzqwX6y
PF+FopixSYX3jvN/udjTzMpT6ViyED3eULEHWNfkhPwsD+kL9CES+40TpIEaBtNV16cphoUFJKKS
qIbOZeuytn/gUQB4qLsU8RizkKsvQPRie3P/OazLYaKwPujw4E2mqakBz5KcGj9jyfxvHhLTWXKP
gKNaIprV5iKUU/cXNlGAZDzJ2vqipJVvz3UNc525iR+zN0xPA9Yz4cX5/aGrI+VTqvZ4LWzksrAO
HL87CKrsN8EmG8qw9PoQUX3nGf476YPqbMiqdjunntDdfgTwI0ZzPbeyFCa+XmtQeOitdCNp81Ll
4UQ0GMICYLS1k3AD6ZIo+lLp71zRGzISIUgKAeh8PHLnyBeafp+BvLhvBukH7WkEADmVjgcWeQZY
/+Z2yw7/8yA41ANOqY7bDtAz+IS4GHeGGOaq0VPAG3srKEdl+wIP84yEvxo+jkKTgTTlKF5/YFkH
TN/wQ3GmwlJkLM6BZsfG7R2+NzaMTGoCExepr4I45+OTESRQlzS44Ip2P4vLPtvfYuoYWj0hT1C0
O7HIYAquQc6pvMophDRad6xHEkkcv+rg56YKu42rjjbmN9HUzcwZiD3P0CEkm+Mf9pRnEuiGZb97
IedGktekoxnneLI1hQec90EAVe1ElMjUAz4jv5Xvx6HNuPSvNOIu+CF79RUDLqvxXFa5R0vIGjH6
47K+ZynfS7cjEtk90qg5RFpyzoIb+zumFNGjufPlRKvNqBqhhhboV1Q1UcjEkJZ/sYzuDEQwg8ro
E7TMk1M3FXMBpdbTUJSjeef+d7zRjL7qmpDGzxG8Vjmf/43nGXoj3G5x2LjQ9gL2cql38wUQodK2
YaLi8jRw+k1asacha7trXd2gu90ogntOW+m8cWExMPH1xdeMbK63bN0OPfvrk64oRRiuj4MaBCu+
7Jt1+gDBcIviKeOpCoTXpjOvBo+6hOjzl4YBwmLVL+2PUwKG97/TXoFT0jlbdonEZaz1J9zgBNsx
lI/Nl/6aq5ErsUdxFFDgBUYp8WBeTIsfhlACKGSriQ/7yGAbrcTj0hqur8zW6jQmb8Etpe7IMSTc
4+hRVEYSSprIi5kZKTpaXnvPb9ExQ8VUhqw2rGLaevJClyw8XGR7w1Uwfox2R8jQp9y42GsW97O0
wd92fL1QHeUAA2hy3m1IyLn5zJ409GhXuc4ARXPcTmVnhPsqMzi1AndYECMGJAZIeSh9oGumCW12
IKPovjiqkd9xfGCnGoqbQngNIt4q6b8La8fmdjnoUwL4jhr/knIA7x7b3sPBoRLk7jZnjOeDTIHH
dXPOWitx1psU0oKdCnYeiHySjvMPc87RMeZGN86wIdNdUMvMvACPHHBAECWccprGiENiQTHhDmTm
zO5ZjAn9aIAjoZRtGM3l9nRR2CE8fWipGg1Ra6fGJlcMoVfFcuHGheHk6TDCAzLB1zgN9YDNiib7
KrJrjthMydYAtEb+gbW3OzfbRK0q9HrEHFwDostA2StbtIkdeOstkthBl0w/0V55t8H2UT+OQ9kO
7F4WFOa2YNA4b8p2nkDAPTyJkAePm8Pj58fl4x8t7QNeyz9mOIGNKHZBomK7Pp2sPE6y5VpWoj95
aA/rGJ5b8wxlsri5bAlaAKFv5djUFtpcGVCBeNTrh/t7HLWdzEJq2nN7rwfy4aEgKHfPr0ukOya7
5aD69WBkhph/86zkdAXSgDaX52KTObALJuhtq+b17NNTHcJfUzcqQc/xOqU8bmWyeNvvZ5FvNYc8
9qqH+YVcoOw18InwxwouVJbKpZbmJsxtVigSVvG1FeXi+oocVC2HUt1FvfAplsN7jA8URzPJpOAj
aNGWnjUKDMZ5PL/aZ2q0Fschl7H1W7+dTIt0Q/U5NWslkVuRqJG4mQsLuHACTm3sza+TELWm43Xf
9txYQFrb0wGkiZaPyi1gfPmrD6WYq7TtxLP3xgWc7AXzPkrPL6AH28dp46gGxUaWV/V/yVg3+beC
Jgs6RnSKwNj6NFLWHLDE8vEaHsmstM1Izt07JqruXhCc4gHvSEsjotgXCw8y0lWX1ZUq+PrY7n0i
89tnIQcVYFik6/CxOjVuPsWC7rCoPRsaF4rz8tq9O8qwnq7EvQTMFmcQ/vCZxpBo4vCnR420gkTh
ab1v+ccq2uaMmfBznwa/1lT3xOhiRCdSl2l2WI+AEhybXTN9/lRGZaEs+e6TIPfBoEBqY53uO8HB
GmBmLgrhr4Mblshgl/60UY1zttvDAja39OUtl/xCfw7Cg7F0M/YvIaoyZfIlKHHLi3R3Jw6FhSSq
VP+11bD0jWXXNESakRHieqG0UiQr6gPvKIHQ5UpNHVjs8gga+bNnRJrHmezmvwcpdtxOcmSm5wXF
kIizlZz8vg1661Rj2AZmvGmrCrJM3lLacBbcfmxZxIuQCKcHVJ1Cd2/EIXjskXEhTpQxizQp6spv
lA//BFPGshfNK+1aynVvDlg3PNcPr0U7tF64098tGeHpimYvc/lZnoXr0UgQx93uj6M2nW4lSL2H
qowN0m2FGLB9X7+WwVht4CfUntoT+4xnwxvomq65jACk1B8mkhbeOgLHxF8xfIfAhBKKqifMAqAE
au40cmD9nJS0EgIwJ3TLxDLZyZ+6dO9LWcwz7TXZw3/50/Tfy38sLzNO3vuwyFeuZiFSrFy8SYb5
6mM0P8OG1ZAn+iOFFjj8movfBJm7ZWKx38oMe8VW6Kz7HhXlG17kjGBeb0AyTdY6EXRlr2Jk0WGl
ig+vtz50FS/I7wfQSXmtyGtE8FjkdG9ymOSNkgBW3gwyXqhdx6NtRJlbwMCsYn87C5B63+DDnkrd
TQu+rz9eBB6BGDTytLnOExwyTXLUDlo99gQwD084ol+e6qwYLAFRakXOTjuViupU1czTErNvcmTO
z07GLYVbZRg46FkIZ6PJz561jW1MdneED9vxNwiog09/0gzyjUiC0JaydTxfuUb/7XonzG0yt8Iu
VpyL2V9+TYnM8sew088eqp1gPUZPByo41lCv5BUQCVRo73KHXt5SmEkyiUZPN7BWj4xygdMI5lwP
iHzLeXcSjlbQMyMI1V7qAmGWhs9Hf9jWp7nUArOjODg70A1sclm5EJunMrO4RUfPRzKEpH93Nauh
VzffUIXAZNIlKJ7ZrlGTA50dTFIB0mfl5c9IoYICxGaboj8GhNcHKUYsfJoRA79sYaWn5X7chB4v
kS5HKXhwZE9T43+xfH9eeoRTkfe2hn32Fl3uWng7MfeWqLaOuFZVzhRscv6UyOLj3O1Yh/r+XU7z
O57erG/aOZxOBVrfWJG7Ik9tEMSOu/1GO6EJyH4p4DkmIRfXYjiOya5Ly6Xg6oOTkUVKHG4Z5zp8
QDoka9H2YNO1Y8qikcCLepzGKFXn4UKb10epfVhMaxRumiolvfjp2WmR/A1hdaE/mYn0/pqrU56T
A+XXtRVBaG9knrcn4Sqr9GcgzeNCMVbU7EOIIH5TrXYs3yNREBEesQ54sMIrNeWRjBy/dsxd15HR
KI2idTPlElaxtAaM4E9Bzf3XFbKITmEchEzf+wiE7cxb0wygGXFIFKZOLzQKB4LveevXgdiofsYK
9cqr9WYfIt/BIqoTLVUBYNtKEA3rR5G46wKf7Yk7so7yymWOwtTxM1KLbm+2tDbz5YtYObV4HG0l
UH9pJh6Xen46HcDp4p0wmvmZsTNehv7DMa//kPaUTw/76AxIR8pPhdn6+vL2zT/lq/pNFcfi7eNa
1z9UuAFdpFaagyLuUBo8fFaA9gpQFg9442bly2z1dH6cOVBUnAp8szVJUvHJL8ZLeDySSYEaCvcP
ZqBUfXBMG0cdIuVg+Mt7D/YX42JuRYv5+TOOnLwQJFO50wNXiPrN0IbceHrebuGrDnEw/BnTp5dO
KEvv1JESp2H8fltEvfI0le+qUAzs49YnmxV0gboJJCpypVDiJVbMuLlPtBKh8utoSqYlXjSjv8kj
eWjWnVk1HtWa+DxGTKPUmZQLHGA2omiQEd6UIbOxm3foTkUQMyVjNqxkOROAxUntRiQli6LY+lR9
TsentbPMbrDF+TnvqFuut7zD5+DS+1UPW1/alzB1DOaIdrD8VQO2+M3WJYIEaPMjxEu1rz0y5VSd
svLzzPpDVhJxcMloUc4oV2LJBgEkjM64F4/RK1L8G8MuTWAPJTf4zVegSpbLmSoOBimNBKeciR7M
VvGGKZZSOP0hcxvsMK67DjjxH08acf3cSwpKG+9nfCyy/+mE3esBby+RLidT1/MmmGE5UcTvkFzK
ESNw0FplncO0Ms6rxgpBywenrMoB/QORE1HWV4ACkr9TZMWzkRZryrzEmAo9SptSyAn3cMYgM0Em
F9zXlm7xZCxnBd8rSIfiBx60Jl2qkNTn00IswBZgOgF0A/X7dHR2qvw6saR7z9URRZnoswDoQYop
y4YyXOtomo+ym+R62xRe1qEQRqCbIkF4YerUvZc+bCeUwi2mrTG4x347Z1jXJsLPGil4QNZcoNaK
HbbZDkhHSI3+rp18Sb47rO5Ppf6HkJ3UWEqqwA6jgY7Av9gSBxEP7KuSbb6YMMOe2DcpbWnMt8WP
sgKLKSCfud66iXOS6sWzydVIclU46Q+zkhQkFiEXL/n7Pr0r/JShX2wpDpocmo/u9r/b5x5O5HLL
DTmlI41K74oYwDyNx1oOnr9w+doPlNLqDDyhqM2YhCHEg6xjwR6SqGC03LpeP02w3JjUeyK3VBaG
NagAZE0ExqYgsgmB+N2STclna1G+zB2RgRfy63eYwa5ajy2TzViP/ug+5Xt948r3MhcfmSv44F7p
GBG4PwV/HPwOhaxePaqDiPRKaqNYUvV0psoXRXefG3l7Tb8IjHIzVor2MYIbw3NAMzZAKltlkdQn
R9+q7EzzV2Ad40YWGh3/Fb5LbnOj7yFzIx9lTxSpYZrGid9AX9JVmJQb8x2forlcKGz0MIdoDV00
TLHDPOaUGokzKYzw04TE7Hdb/KNY0DwXTOf1l1k74EC0yVunbbGznLD9nhFZOW6mwXVJ92GzFP8V
fNHbP/iqGzcviF02byTG2zeSSVdNz78wBhlY6m8rEnrADH3B/hqwOruaEbmtjI30UQvp9m9AWgy/
5foYkbMcM5vxKi763X4FSg0qIb3Rio1csf1qFAAf4sa5HkLM6k+am3dxabTmYDevopc8sPmlNH7q
XC9ebb2NzPfqKkTKX1VkTeLnXB0z8cgjZW7sqxLcAJpjyebOxgQ4P+fziOsJaj5EO5/ro7MfRd/v
sabi/ngr9FBxcuyxKoQ+FNwAj61yr5sOBBAqJaOSBDz1d6jszytFnovceaVeMRw7SiQ6qgwRR0/j
YWQcdSOqiumtpcYHwKLr+nDYyw3JmuH7pC3Jgs4Eb7sHRH7+9Ud9lyMkfqFYxGuYIBdrT+TritNG
gAfPEA7IvyrHh6fwO1F+aJUWDbQYCZoZ03q+4zmBaqcxWsWyWWaAOBoTHYNugTpK8afBZ0bwpP4L
w08PLQusrSEGQ22mzgljPqcZHB3rNjF8vZIPeOKlBAU4L9pN4QO7RjS4npYXUfDfc8jWfVQ2jOql
c0NC/qfjY9Q2YNE05G8kwd5QKS+pAAnvK7rIGcHAqSrDecCZvIASP7kIqSlhlw31uepxAnwKwSIn
BpqZImxRwaeQQaYEe4SoZBZxedS3T7x4URTfXUWyUqGuBpd7gVX+zu+Itoy4QO5nBgy6ACrvO1Zq
HOLFy7MmRbH5kQJEbqhZiz0wrUkzDZ40mWCjttjighfJYRIk1G42e612m/ay6KxFnGgTKmclQHx4
WmEN1uJncfYSMfGZw1rRjNvjO4cM/yzgU0IOa0JEZAeU+jTeWd3Y2jfz4SiP3wU6W80D+aDWmRwm
I6+jbJQ0TbS643MIhPLdxnQ4wz43kjqR2nup4Yd77yXFFPSqerj+IzTDJMFNhrgS87flbA1nqmcD
1iN3SttT65AHVO+b5kaSXI02FNaQJ7zdUwru6bAooeaFQmb4LjEbOEZ+HO0R9UEnXY8H/Nm4JQhJ
uDM8wus47IfeLdUjOeiVXGZjPExvLY4eWvnwvuIz7NN8Vl2hk2UgkF2p2w4oB3zRF+JD+sQTABTm
9wK8AN5RkdDz6Gb2zPTFistz9c8JOqK7uEMAYvtwLCMj+XVhVUP0InjWUmR14bdKBDcovZXkmYBx
lciOyf9hxOOFc6GcCUyq1ArW18x/wDGO3Lj0OovKegviOIK8QxaqNZnbTue7oCtdu3x42D4kdSOf
8k5+HpYyXzZ4HCR8tH7tweEZ4bkCLvuztEh4u4Qhr3K109iF4RnjTSCJiFQXyvqJu404UTYS9ft9
xzWU+lXOLacDEo9oFPoG1wq4G4HUG+U3heni2HZFv1ecUovCGsmi3+YH2PaVKKqbIApmmYJ8X3PN
g2/FWNiMXcWnScYYFz5EEkrDbdOkEPUOh7aEDlG40nS+qj9SaqOOpIzuOavSZoDTTt1ZilYdZzul
8UzQSwK+k5/cFMsnYPKtybk5fsld3xIfu/Vp4OaqlZtfwRsOGJioiy/QwUk+9cLnM1LW43SqhTa+
TlAQ9jhSvqvB3uYoLKdH8TQ5CZLSTOTFGNyM8Pv2NwGVS2UCNla1NdPt6vUoYgOIh5gTCTfUxTfU
2UlhkDYvf/jeNdZt7c/sr43HTcbIdw9tI60MS/foMyW+sebjw9BpzBUbQkkaRvSsEwN3R98fg/WZ
1wDkSa3JLHw86vbqRNaNEUY1YodRsEC4RRfJVHKDyevSF7/WIKPuOoNowKS/JxBnxvnsMCFo/TP3
+bxaEin881vjVNeGBWsDZThfZWjK1FyqB8GEzyYgOu5yjmWphRFQHDlgxlP+Aj5vKAu1S7zvQAuy
KuycCarqWsS8s+rYMt3asL/KRa6dHB7i2xP443otCh4LqshktSDGORl5dSOJTx3/aHwjl2te8XH2
NwvrPMYTLSUa2X+1wEw21OCCqhbqw/O6FQ+mRh6GGLgFntq/wW6srxFmECznSoWZTaduCbElXJwP
q5oX/IOl4DKkz5g8gGRjXP7vxj4owZ3lKbxUBRiv2bHWWd034hMGa0y7BEkTwuDJ0QhW8/QlqWsJ
bySgv1APc73NCZO9+jdoXZUC4qNp3xPcHLpmjXlCoxEwm/jSyUUXPxsAHSz4/82Kaa4d7cw5ARNm
3lU5E49R0iqPxuE1QC/KNSbhe7rPioInPluAjYFFh9qnqwVazsvwn5MRABNTVNkIEMUZxoSY/OdV
JA/SrfCl0oE5Q82202xI3cXWXG0ItlsYSboKfBCaGhqMR3xPRseNuylohm/Bj1Wb3HcafwTtoavC
8Cuw6A8mwOHte+fwSsPk19LeTNsMZacgcwe/7q4gUx90VLbGn9mwJnlxl9I/2UkEHC8pQVgefFTJ
fXIA2c3j3gQH+/F2fZeVU/vgEnkMpSKGqH151SJWGIWXDf/gQeypVIl2sQgT7OkwJpu7axaIWhne
LsVX9PvxVonaT0xVes9ZXBv8g+5CddKi5ygutCATb1nbvhoW5nor4YSM1zxUrah431SLbSDXIriG
CNbVPo9Pgbkthkk6dk/gULegAqOBI5ra79ftvIOt6pqWOaL+lM637KKl37LNTqeGbcH5LtQkIgy2
IwVluoiTWrcJje3uJJ/zBBSmkxJkRGZPWVS7OoQOZlu4QFDduVu3y1pgeO8CCcd+ATUJhlWZvKjs
oPJb7F0nPoeQ/Pc0be/iXpJuYMSI3iWM201Q2+4ygx6zd7EIDhwQBJrqgX1rHd3LVxYDTRzIJH+8
7iOOm1knc1FIFRJdgEsT/+vOPItb9ZKHTC0hsYyXcrH5C/zeUnFPFOyI0Uk1920/og/hAyY7sE3h
Ysz8xX+ixG8HPKAl+UCOh4pgtCUoOdy3hmqD7OCnD9euj6sIU7V3p53RJMH0DnK8p6F8GcO8WRaq
ATHgJMr1hrGv5tVSVBuesHqsT7z9GR/1YAO94oT6Tt1DVw/yNhQroEk7zDq+wa9UxWOwIKnK+RTK
WUO5aFVhy9pkn5znuew4zL6bVpTK9YbniArjfV9VmpeWVPs13cyb7mQfxHg2FdEuFVBgFxyegCC9
JL2HoeOQcYA9tkJfmaKoQNXa23nW3Iq1EvJD+T2OwoZdRROVQEOIT8LH1nJP0EVOFg4tdVGhj/V1
Gbq/gf2FBVTMcgez1Qp4Uwh6rCGK4TMVFo6rEvpT6Adxl+LGyjIrlEWHKqPlLk1d7au72rvbDtg4
BOurhpZcVThn/d+7ZfXXoRH5DlEcn1lRg7lXGKY9NoG5vKJRBHa9dh+wdh1Sy+sNIdpqZ7IMiOXQ
nod7uq8zN6GhBfr6OHJtuyYoj5kZBgXC5bR0E3bHAX7nlgkhdYnCxQEj4Fo1IGjk4T0jxopjHgkn
e6OIVAiBuWaRD3X4u6qPgDs39tyy8ZurJPuBb7ZvO0QgD6tiO59JasJ3B+ZE7Iav67pX4ZzGY08b
UIxmYHxU63NrgYqzOwStz+RuFkP0c46xRVPNw5jf+NgMHrdz+mlhyAudtT28/Bsyy58vRRfruEKm
5rDv1UTSeluDbBmbD/0R3eRLICr/5G4Cqa/HaipIpsslT33/UoFm5t5Ecv3GJ3RYZdCxuRQ1gn9Y
lI8RJ5odOpgL39e+KTmgUg6Kw45U466rYl5suEWaN31Fa+PVyhi/aKFSjXRzRzHlsAUfgrE7W9dQ
tf0e9vnxgIg5YHZxfFcTT/gb8ncvzbi+ra50TYiFmZ7lmIGou2dByrQZEG109OPdmH4BFSBUB/O/
zBx3aPxZqbpcwZEL055HzXoFDGdmShcLxE/t/fCcJwrVtpMX5FDzxJ7yIGaLgDjJOMc9EZaIGfrl
wmbWoCyMfMPpYMy0b5Fl3mweKJjx/gFYqRDCIxAwtE88bzBk0F6AS7UYGKWTI52BuRdB+ahg8pKG
Io+rSeXphBw7186Dxjz7uhxlHb/CpsN+ZWPDmT+iym6Xsp6x/PNT3W9/lu04Cr4kwq3k4Oo8Wev7
bsmyVLGmm2OJQcobkkqfxo7nYEwVftHnlTJkC3En6MW0u+gUnv0DO337gd97MGbN9HlP5YFdENba
6q4hBvJyDR/aGLI76ZdQPiFHnqTWkwlA0yc+AU42jim5MviwsGk7W62N7TXYi5sQd8xCN75ILSs3
vrsKCpQuN11imNa5vdomcDDAbXtVQ7h6AGG4a0dtw9/eLPBI+ZsyOXcC/XeW0Ug/8u9GrR+XDGU7
Bb7spSarUHh3lN/yaamVNq0j0QMJV2g3Oa8qBlgVPW1x9GvB9EdKDmhhzI4zxmLNSYGL/Kbxn1cP
yLpRjfNlKsbnTae+twIxHP1L0rzBdz49zxItmMsIoHTLnTomIaE+UoImuL4duSoRSzOTeiLf6dVs
VyWnJzRfXUEinsFoq3OMwMc1btrHN85NpSKX0WK/ieZyVbU6DYyt4QzeWai//31EIORdp8ROPNkk
WRvfEFYXCUzE1Cwy/mGb0YDAEjoIcvaiSztV2tjqQNCjQwiXNiPWdo5o9IoNEf/f08b1XTMBzG4K
B0W4LuF0/C0dkMK90bXd5Za959BSN8TU0UkXvlWxZGDVLTq6t9poEqJf1dIYDQjME8+wpt19UO0r
diRTkacdpxrrCYuz2xGWPR5+onuhgyBgTYej0BQLj2GM0AHbNZeSvRpDe3pZsqXf82wzeAMMJQ9H
2f7CSxiPMdHkm9s3HsAUVt1NA6aHC+Ht920yH8GopkUgW27S/LHYzxDadtWwqB/fDnaKnFnkjbGi
hTGbOvhdfDHQbLXVf6AU/O7Ac8sA0WdkPWfO5Bpv2dTMtXZ99xOntew7ok3duiaG0COdrpkRVdSj
2dGEevgh8rpzM+tCc/ONiySCf5YTcTFzkOfjnjM1hv3AUaIeknnZdC8ZJmHXf06G8Z9tvR5bZ7yP
ZXy1RvqwnIzRx3D5D1rBtIUL3cs2JynKU4HWmuXnsf1HcKpUEglO9QdVVpkB3alcsLcXu+tTb4Qu
FirpJX7FoKi3hgMvrXKVPnYwItWNxb5YTHXRrcQGBHRzvB4yN4rpYSJ4+f5Y0+oK2WgbqEBM6wif
Xxm3sCHq4exYF9QxOUJpcEdaCjdJgVnf+Jvi5TSTu/SuNd31zSkbzhKoIZr9pfefef1CbqYi5xan
SJdj1c917gAXoERIM0X6AzQE+asU3tebf6CGy4EH6OgwYCNpL0A6orqr5s3qlN8n6rwrnv48uvQr
7+Z8o+VfFm3Vx++hJff2mIQREGMcpLFdyjtBZnMDkQhxqDuefCrgePFZRIxWULfKY/Npdd9daFXm
zgEQYO7HdIj/m3d2SlNrzadfkaO9n4faojhfRUqtliYHdHptJAynMImQDzdTbo8zgLMrs/2JPV+J
3IA8mwo13OFX4uZw21s9mbusczjCvVGyFFG/kBnWbjoqg1q+gqR2rdKw7le1MXRD6zHgKFUHIyHd
4JBeKoF+Qwv6DkDWg57o8ykmTpfE7s1a68C+0RZL7wge1lyEnndtRP9mg+/e7goBmc2+e+Lsk2RX
85VC2F8WgnQhALs0Tq44JAhNVFKJnGKwNize8KLW1zz+9tlBt+hlmhfULcWzy2xfNP5HqWtPWwxU
RF1lzTU7f8CJUqXWDQmipw/5BNNr+7lZT3jFi/9K8iEBzn2iyhak/Q4CzV+YKdpaVNrRRzPr98Xk
0eLNd+JKT1iMdRt2KwTSZBJlfqVaFWdUfnE5gpoTuBv0rWaF7BFiQ99bz/P8GGBqE09J6wnZ34zu
UkEdga/+y++ZnQAEg4/5L9+wHXmDufDfRrN/Lyqz/kvkI2JO9R641VisoYYfChUEkV8ZitW9NVPf
QhDbZxZCX5gLkVP1iPk/OH4BF2J6HMXOF03MLKvG+t9e5Slfna4zrRFVKhVwcYsAgEVrJBMeARxw
j4MEyYd8U+8XxZw4s9DvU3GhVykiMV2BuJ6xjk9dP6Bm6+ImGePjWzKMfFMxywoDG4WjRXDESWpE
W9H35sHXBkZmfkd+DwQBUph0wbqU1bFVO4N/5NToNRzBmhIxmBPoBJaZp+9r1u9Q90eJWc8LHUvl
0Fvxx1QTJTcs3diVUwvSSLdbimjlFkbpgv+xJj55Wdr++p58YXSoffUuKxI9qxbyZ5zi66JEyHyw
9ir2hRCHm7jWgeUk7Jo99zDSE7AlOCfER9vDtdzCDonNrfTgndX7UlYmBcNk3hnOwUOfvNzzD2v0
2j4mB0gEiNCM7z/BKAd8lD0iItbGgYLVJRfyvhFwYirfZ5Nn+YtdFlVYffoEPx1lJNWfg4kncZaq
ZlHuF/amD0Io+Roa4XgxgsZHJVj0S14LSl0Pxn6ecVn4L88Crsf/te74JBvi4++nRGGglF00H+0O
w0j3IuDppUMpjmgsgo5377CW6ESFebBZL2YV4u55r7L307wuvOTEw8z9UKlIOMEfqSRcON6Go0Rr
Y1nDHNIkv43Ej4TVUYCo2fs6LpnS85V5m02AYWRxL3phP777700exYl5rt9HcuybdGrH2UsyFk+J
NSqQp/U3uwlCD57FSIa2lRgirLlZNVnyEVXBC27uhwZG1bGDZP9d/gvy3vuYFvJAmFUy+KLofcxs
0982AiWBakn0svgQGgbYRt+KC01BS7opxmT4Ozld6ZHGu0Ek5PSBmx6rnmZ8XxI8SrIjLz9EOosL
JaFnMX4TL2mYI+NxXGdxV26/Zhzo7TVMhWzMLpiFOQX77tkqRDMrqGu8CSChMi1HCKe0b96CsApY
VD436zFKoi2Bgly37Jy6q3Ztyhw/nZbso9sRA0e+Hh12RwyQKax0TgFawYQJ5O5X1NLkchhGOMkp
ZWj7ADrY7hjZQHncKCoTNGbukARhOXJ0muHxh4/gO2NVrBH1AWVJ4AdMKGrD/F0fmKR6wF+mbelr
WD+K898dfcbCG5zSc4/ijIbXrggT9wiqXu3UHyoj/0rYVtbh4U2it+g1vC1/2irJWZSPnjE3Cj/T
7yyMJ/vXNlJeg8EoI55k/31nT3dFQaeFpyNkve4FnjGh9LTsZvl1fm95dUb8gFGg/f/uswMsSDMN
4QuHU7ObeyJvZ4YcSVNs5UnoE2FJKz5QEJz3F5tkHkYJd/5DaZlCZmX4zIf1P+FafrnFRlPELLQC
74pe4YmMiU69PKluOKD3rQHNVC/9z9HfZEZnydnRdIPZ07UZL8rG8ELuzCem+QLoeSkp99OK+PvN
QnUHMYTnrYkU1mWMYXoSa7Mx3OeRNomOqMDxVVn1FNtgYkptjTyBhuWm3tlNDepqByhO30NW83Sk
vkOCKdEqnmax1pPmUFo+EuhW0wJVn2iKIICoaZ7Y/CngXRcSYmXd37bhMzsK1moudiC/fF9v09iL
muf+9Tjr59skOxako9IqruHaAjS9mUiJJXERmDnZq3Yc+pax4+5WrE2H+t5Fc6Y2BwlWsbod4Y6B
5UjLraWDvXUodwz2Pvk8yNNLoYXJCvpQqT0ovny9izg5TARJAPrmQeRDF/+gSRHTca57Fr44U+pN
KIg0jfaoNMRfP2KmEVqHSvyj75kWWITdDY9tm5CRmn9aZQlOFC6YjrQ//lnFifrqILRS4QEm65n1
cuphHlE1Y63Hp8VNW3hYwXF+CH+rKStvqTPKmtrD0QE7Z1gUjFW5PW9/J/ZYM5GdCpSRcmD/c9J+
jJwMJ9y1C2ACTeQlUWL7x+c+qgLf18F8ConteoBohaTM/RMjFK/xyqcE5WWfnJBkiGSjQAfgKgVm
CVPoTA8k3igCzlfMruYp26B6PpjmgGrGiYnUHqxmmQSmiTJ+20Mha/OchE4fKJOWUVRZmM5wIEbh
iZHC1FPui3h5DU/26ZsOgEwOwXuoHTU2fpHzFl6qJ3WGTp8pFcAKSoJ0bEg7ZOnfqqtK5wZClKIL
rwysOlxCJH67LBWvDQCapRtqVlapc6cQzq1ZOsygXXM87P/CLtSXXcB2ZlGIrSsG2QQRrYwstDH9
NG7X05a8sDtpiLGNk7s/FbLNda5G3dZX4zvgmttuljgGtevr/nr/c+ZIRUbL1uoYvfQzQvOgtno3
m8pt8IY78qZt7ddO/wchM2SZkfpXnMGmADcbHvcdRfxL7DFP/Wt6NLHtrSKB0jwYVlH5orXq/LTi
6C7ohFtLDaXCxY+aPafcv0ARDd21xm/n3tIdBvlRm64lHRAEy3bEz/fqajaJUFJs4sGprzsaMo3a
XjW4p/sB/P9pk6x2rw+AV2itQ9e+UYaHGtoi176RzMYjkjqsaBObtnmQ/eobmNFz8iT9gZS4jvQt
4RkrRhD5x7Ow0cP2QUjX9g8b+oocBK992C7eECirrhlzS1ns1AHvxlN5kCy3kh2xQ8Yb1cGlIHa/
msc4CeS0lR1xKNQrkpicKcEaXKSSZnfmnnOs31Y+1ShImW2sVPcpRg5CARFM2i6bW1P3K1BVUD4n
kxfIuFmKa8Q4gwozNFEG5PK7Tbv9bcplkc4h0HX6OwbCzVSuGf0BFFlDgeGnKKY+o4XGCvIi4fbG
BFwLlvjjQX6V7szCfhDXZlsAQSNKKcwjbAGVFA73tHXo3BShE44CrFbz91b58z7kdQugUja5SbcZ
UpesoJ3hlYnQvstUkhRfdQD/D3xRpH7WijZyxKFyZdFJ03Gojtzm4uvpLCrsAOsRJF6nDGIV+Cxc
SuRAhqs4KSPaHcStP3iyu1bnyjnDEDwip2KpIGnR+lB30m1qO2QWNe1bZTJz7H8yAvw0xVQUdvrt
gsLLjBZMtMX7+a4Zkmfvb1Bcr6qNNMLBHhxLD+ss/zojjk8DZM7oOuVgAwSnlIf5uNLk5M7D/cGR
+4cgdqFb8gf87yODVT3mmr9I6G/p2kMl5pGRHBqO+RXF61lEYZGA5caDyMVVA8LtIbF8dkg/ZUlU
N5Tu7JhUX7UPeZlRdQzKBaW/qlb+TFUfmW3yiGsiyKy36QhAKvp6uvw699pOzL4ec0fQfxxSMmHv
PF3g2gnsdFZjA/sanPsmGjbFQnL36cnJnYcxHJvyMG3wMFnjPgymVdEC60zUOvgfu8VXkySpRxDi
C16CCWrWOyp2LI3hxV6R2qsvtXC6IWOPSQX4yqC4TAy0JWFpackGoBCfaHpsqfw5Y4aJI3pqKI0o
1jsOIsd+OJRqz0rMBesALfIVHfnYqnG+ccXNxjc0DP7feDAKF/vMggUBDHEg3W+oasR1lukUGNsx
FQhnum+hcTONMm/xtZ2jW/YgWvK5fqtGG7p6Q8v4QbGLitA9EwGcJxxOOSNdYsmBoB2SXIA92aDz
48U0fnhTEJgEUiD6yeU/uYWmBDtPu/t/4oDyId+FtnmeWSg7W8+0d+EfVhzXwhSZTiigF+kdmakz
fHG2w1XVaKJ4y9b70/1q9dfOERAdhBO5I9FgQDKIS/quoe/t/MAczIFzePUeVUxA/CQIOl6NYVnS
tAEqvL9p3Z07lhxXq96TFMEhrHC0eehmNG+LRi7nFMFawoaiLw+x/GmyIBpYbmm8qBjs24jESrhX
ypCwX1QLCSXaDp6bMwM4cZQmdMEqnDpvmejYsIgZhY5SkREsKLozDq6gTpR9bKRAtPKdV7PqXr+K
87MhI/ep2o6yBkhDfaXDY9ITUxT7YP1FIUt5A1U1LEzJaWEdoHqiua+Th+kEmY4A2oGFnVdopu9P
ziI15kh6p3l7n1mnFTWnMP9RvSn9hzz+7UAjLx+AYUkSJ9fvKWAflZGvMOrOpcnAhJlkSpZIgCOw
Yhg2LrmvuiWY9zYSdCLwg6Kfzs1B+HQBlC4I5IKHqeecsj9D/RsGbdxvxSEj4EoXNokq2j4qBfko
RlUS3L9ROcK3LMKI8P/wK0VgkeWGF6E2zPGH5zvj4GjjOe9atJzf3r25kp5A184DPTVYI6ZLgEIr
lOM0gJzWe1tc9hh66sf+g5PDZidJgDw4U2lVWwvk4AID80AsxHvFP5gD0xvjoaeIIdSLKFu8z+YI
OyETirWbgLfZbrn/g1yAqrxiMmUIog/jxTl7eaTUQLZvnQ5Nil1ho16taDOzO/qfe7XYGUw06xnI
e91HoqeGhGbar+FV1G5iI3oR600WV+FXE0gX8k9Sb3SPjYhvumYj8F5mPvRKb5rylXze7cGTkAiA
Mq/dSBoJ804+tq70Tn/DSyDWBnAnVd8oAEVDPN5t7QhVYczPa4JR3hzOiwZcCR0aarIJcbzsU0cx
x6hEpFBkMnnQK1xRMyXk05ssAPGaR3K1G+xB4Ho5ePh/i4SINrWUDVWMHmtH0TEKfpPFV/J+SoE8
jUlb5/+dt1orh3zFT0JSjlNPWZN7oyQKfzifSJlm3Uq6QLf7mKg9/RsKFR5DblzUhk2u10l5EB+1
B525VMEeBOb/V491sJLTtXvaDZXVIqaaF6++uoxyjYxzs+SeXaqqbIpfGs6hC21TdV1vbE0E+g3u
7Tn0uVQC1VCKrObcT0Lt4s79MdutSs6ZZKfaGOGPqc1o9n3K07lHULgl/FGekhqJAwFh1jd0Q5p/
EdGH2bSC0dBUim1XuyZn4PhyiFYTk1Jogngq1di0uJ3RgWdwrAsbRazSeWde6qsuivdZF092JFhD
HOdSvBn6H+b7oKlj5+tm2pxWhQEFzliptYby3eTH4Okb/hWAAWy3TVp08wMFIU5j3uorpiPJpZUz
mFwCzqzw5i51VHknzG1poa7zop9PRlobDDukZd27KhNToqWMHPjPxv5GJTJNP5Ar9v3Q9ZkFOHKR
xnLN2patY5Kw1EKk1pjS+xZnvC4vD8am11M18PaNkiEhKPEtgcRIxDT4m0GWGi98lqFLcC3LNpel
H7OCrcd3oTMeBKmRQ8zxK2T/TU9o/1meon1OFXMNGchy3fi6U5t3EN5lkRc/YR6LTJw1clFaD6q4
MlKFXrnZHcvzbnp9300Cn65Y4Cnl+znstYHN5CC1ThV3ABowqz1ljNHmx2xrmgqPuOYmjMvUBfpB
25UyldmlUNTRNk/dJJiMgnpV3D6CQdzneL+c8N7I6TfHOtzuSIr3aLPNVRV/fvrgk6v5lO394DaY
cFVjQpt4tdf/O+hCWmtuJ2DslAJWH8o7tsf19JrlZI4zhh4pfLmGCu/YD/Fit+D/70dPn8Xni7ti
cIkHWWHYEdEzl+a5F8+54bSvRpwf8+R8xEXxuayF5jb3eAZOhbIM/cYqVWg2bPDqsMyTUERapZBl
wkzQkSW8eEo4elclPyzHGWksxAeIME+AljQRYd4UnYPIboEEjd2CQ+wvx4lk4ykFL6t65ynDKUzj
o5Y7gWCvCO/yAPk7L9CZRGryrt5IHDAh4FZdw+B/ddBXIJSmaYucwmk7JACciaSoD8WmhFiorWxs
jwDzblZnPRPalHx9S7KNQo4KGbCnSu7grI6iiTXXFFnoLz+HoVJBmUvQw7YxbDkT9q8GulC4Wbxt
6/SHN3fNIPMN9I4v7JKKhQ9ZNF0FXY0wPf5OoyYf7Hhey8gUHC2zrATX/xCvrhUKEXqrglRHqNnK
3KSOCYrlgvEZuD1veAS+CtSO0ZXspkpZmgfdV+njLKFXLv2vNVrXkVAxoqsm2iHQDp+Z62z6GCrY
890XSCUm3JKR2L6uJCUfuXmuCeURNaBHkRjPVHAEY0O2+ZAgPLpy65IyjVBbhCg+7J5LD1MG8arK
d8H4yzh1HASnexRtPl1vzSluNEM619rOYOABOq8r6deeA8OhpTZNShHFs+T0DCA+qzGh4Cxt/+2s
ed0cmo0GZtDBaOL4knX2PMAggX4v8jRDamAMp6s8jCf7DC/pGTGBX2oL8uPOwFylr1Kq8RNZtn16
sYDFVOS7NbDOJF03IXll6TdI+LwkjioJRdqt5Tk8aRsXg+eOtGUi+8LUBH9Mpno36VYktjdvQh16
Kbo9sY/LZg9BqHwvGtnfK41XTxmGnNLa65UEWGVdoQwgYfkXM31erGF2Tlk5zb1r4fnZYNh/jI4g
FWykjvptG3hQtx+sHefdnhzEn3FV5+rAJY40bSdth4GtGEgYy9tusjBlreM4rtbHdPFfO9YYPKUj
7vaDhz4z56CBWgIFxjcd0g6Pgd62RS4m1xy0Aik281rcxVhddNo0SFcsXBe8z6X9ilh87FtxdeFX
6K0hoD5tYvSL452Ai3yh5qnYASilr5lc+NbCDtoYwN1XoAmy2bwnpGstcxJF00OmNIbz6X1OaACE
1iewZWAHirPIug362ARs4e1AjQNY+zGPTUsi8emcdohHnGHr/s+I31tdYilJalCvP8XnhcNJwiag
I8mVO2IlGDyC278w9RffMyxm5oOUx/Q/PQDEBx3XcCzOXSHau4LQoN64qQBCJL/1/ZjOXJdZBB4r
kNl+WoQXMggPy5E63f/7vQuY70CRojRk1nRA0iRRhgS+XcHchq/Xi7I06ne7QEPQMZuE/EyPAavh
u4GV0PhghwSDJiFat5iiTqVIcvymGgJUOKZdv1ZJMcotrAgA+XEkUkqT5AT5n6HR/Kv882NeMXT1
X92u4BYGv1A5Zw9nkS+kLNufefSx5u+mk9+aKjOv/xnCXQRriQXtVm0QmuFkN9tfhAF4eqp7g+bD
HyDANPkur59nBqMDiJCIx08uaxZTz2pBLCITxKOhgW0llPP0XXZ/ZqWPh2KRLDkjCqFeM46B24AF
HYQcq5qIlonoopTokMqPzlWgGVy8+/P1daa9AYkeBGVYFCxkCPeftpCVPpvlrhY/Ve1wJBklUB7k
OlXrVki8gSiarxS7m4ZfCQx5uaS7B+UWqRz2cKfeN0YeQbfYOJjqLpFFq9tG3uGDjfoQ2k48SikA
q14kPR34kbeTOEKLbG9eKXXOfRyGPndNEvLY3IQUfEhHougsHQJ/bHItk8jeD1i2xe2LXkjClyNS
zMBo7hxCTrdtKpiiOlpRcgSxXm6mlypd9eObfMoe/U7odt4xwPRNmHF6fH5BLjl1orhupfI5yZCL
VpChfsif60JXEmKLXjuByLk2t+BBP4LIXf4cxIYPpGiKBoVUnqY7TwTLjUlIgFBJb+kmtOu/HJxm
0dGVLnWl/1cVK/dnfsWNe6Pvkcs+LuaLOekkgctcsyDBVhhuETlkf53H/SfOnRo2y+aceD+K02lr
O+Vru8DDmZlXmH4NF82USiBD2bQ6Wxupd0RwGSRU5UWx+r6o99kvK/TGRb3qRlAAy6oTwTQj1gsq
1F2nu9bF7j0Nd21bNogqaaSAsRkHZRB0Q4Nf50xs6fETGg4b0zjc0bYpC4BVZ1I5F924Ywlbz0Rv
hYrMJQ0ou1SqOSkOd0YtcI0yojAG/Emyo5XFxCCQSPnGlbug5xQ3sJyVzwWzo3avRPYOfTREUKYJ
dlbuXdpB59uEa4dsVo87B62YjXStnwkbvyse+98U8P5o20AgolwjATV+/w3KR/o135wSG1DhsHgr
LMILnKDkLD7kLsUVMwcxvmLcNTg7jd8z5GfWteyFsm7mBVcLK9NFkjukd9/AxWviPYmWoZzUJLWP
OvMh4/KRaYOYWc9ORw5cDpgERfpHMwdGxd0uWCkQEQ2eQjFJ+SlHXqkqK9ErKbmMIhOmzdXx2ILn
+Bf1a6C9x/Ab0YAIwnfWtiAoFN17ogrJ4o5VZB9gryp3WkGXmYMbsqShCiiHqcGqRUK5SfNa/bwF
8g/13mMimrJ9+Hx09gRflnwGsb6PgHB1DNDeQMrIrVYncD41F0oLusP/F70Oe/EHTaAGyC6CQ4/N
uqqYocLtYaw0e6QdptIeKC/3rssZVnKMLuFyEGSzt/P8LkmvhfVj7L+/zhQyUsnOCMWM0IDeAvp/
jDUT/yxQyi/YhKETIV65cVf4zwbIo1QzmDq5QL4PkSbHqN4b+3R7TumjKTgwAa+ntweG0MQDJ4Pa
qQmwYgRBaKWNgdgAU763WtU6+8AO2z8PoIcF5AFvvt+gTkXWR0XBITDSI9GRikzAuIY7k+RROv9k
KL2dSV5KYfPjqkvK0GIVikLj5/P3rWMs66ML7X0079YIgeUeEXg+WnhHkj2F8dgokUjXX4oHcowV
uZSwjmAtIKwFcJSzSZtK3Q3UZDoeM5hiNzKV/m3lYWyEDz9OftX5m8Sk5oPp+cIy+59wZiPFXnXr
9taHTOqCgtOvHQA7zKiXD4M5iEAE13UElD0n6Dyz55WpuRlqjZ+D2SM2FbHXVWkwTuj/n8lUyJsF
rs6k0OjClkUYawCL3zRpKmIITwizM9P+kEgv8A25U9+pMiDwPxxMKXaooWRETeANHIWDTP2EN83O
ZmA7P5J/+wqluLGy4M6k49OX6a5uHSLjM+Q+11Uy8w3D2Rivc2s5RrVlZEloKPnKZst0/hF3B/4/
FZUElInpsSe418s4ouvXN+Ihl8wHsTAvQwCswjLrZ5izLqkyqhK9ub82Ba/VAjTzSUNZGHr3TB0m
d8UxY4i938ayUom1M6E5P2UyJV00Kb95Lea1jBBmVoz/wSdR8kulw6ViuCU8Amo0hTW2zl5/G/tQ
YtPL7gxGIZc3ZdSvb4teXz4cXrJ+jyez/xoCSW/gauOeJqyMYVuoyGJsO7yj3jjhxRZLmfpdxnbO
NoA2DCxr6CubANBTh93f7HWtfMAaXphOLQFAFIy7roFehq+zpoREHkeZy4yGOggMh7ydVRhtNgKP
MFPJywG2bsKvIijnaRsTUM2b22a/NsWpBHSmaEiaoFH6QlVMNPWbMDub6oByHkd2NTszLHHLiw+1
dFSPMXN2CpTz99syvgmxv4fMQMFM3W2UpgKzPkgQ0tyEZZ1OZJNeIAf6EA2DQAfesyCLDp+3gCoU
ZC1cQaImfAPcjUSLTpflGB6qChB1XRYT8S6EmaJ8dM6QQvMUMsUi6oWcOcic+Mle9FSlVeEMyWNH
Az1aStbdAdlV1vqM+eYQFqvNI4WchjQJzwTFpzVDHEnayutzFi579HBARTYjxPhPalHyv/7TWAqv
Iuk3Ozdokjo34tdV6p+fVcRUTXr6JWzWN/v4kP1Bqyku7uK6ZF3vjAo8+ZTuBRYa/5bTj3FhsQ6a
s90upT78dsMayRkNIiliXH1mvpjgiZP9s6ZLyWhnI+w8+Eq2R//oqooCecxpl3oKRx/mzzaVBtAw
01jiJ0u4HRxTQjyFjYZ67Jwv8U57xRZ+EtwQ7a7xVQPOp9W5AVbwo6mv2Feah8MQWBDACawXqZpB
AfNqTPANnRtGep61PQiGUVxzaKlT8SVSyJMYxdLD5LngPJ9qf8RQY3Mjh3KY8GnDtYadx4bsebF4
sSD/JWP+tl40KycY5SANlUfiJ2kUJ66AbSUvVILmvV1mTZu+9c44Dxeonl9sHGNp+M48GpYKGUDA
wcvYa8OVTjTdINhPcOcE5gKaUMVKeqSFhgmEkBTswuEPBn4FSqoHOAZd0PR+ol4u716I8V1M0AuL
kCRT+b6giN8T7PbAGTZTJhatsk1zffr/vh+uD4JC0R1S2nsuRM5FRee28bS0Ajvd0aZFLPz9qLCl
CLkSt9G8G8Om0BZnmU2+QiDB1gPad/7/C4Ehst+5Cc+gbuxe2ZAAokMt1ieWxN9NnbxB2dRiieNv
/xGcX2DfVihYpqkj9SluBif5P7Qsr595o5rCXJA6monx4gaH+Nl9MO1nKdvDETeqM8fpeRaZ0QAO
Q3SowlbGbIMAy4yxeSNGnKmNg0AI1jMyVME+9PBtmX2mqIx5lHcnwFAhkhowLFYanWrcx1o0NI+U
i72Mjnd8cGz1gPWPM9Z9pePuHu+wpxkfWj6o0SbOnSzgTu2YavX58mlfCjqXCDrWqmUTTM6YRttQ
4kEZzboUX0Umfuf44xICAZXxHMMfsrQAbIDn229FXHO4NCXClSvuTlt/9KyqzX+BRExm58QooiMK
effn9jmuVhBFT878rUSC4KuHep+wZ7wjg4vw3Cyi+xBDbBojqkvM2e2blnDtfOp6cFAtiuQrusAu
RYcN0Zqlzpq44ft9MIr3RDRQpsj20ZNJvd9cmP+bI3kc7MT7Zz+M2zibBf/5bVsvfp9sdG+jBToe
NS5UrNjgKp2zVsIgIdgVDCxXzS/k4PDE+os1KhY9/HyYsarA2c/nRORIQafWUcBQkCbbXrYw1p/E
2iXaHQyymIk5EyQC+ptrwkOyHThgMsiDzJg1GYsXsGVqRmZth5Ev3Hy3pQJWU+U7feGe7tz3TGH4
cVgTAY36qmenEHL+0u8UypEKKwii/Mz0E17GIgbG3XrGzFBDU3UTqZRmYjZBpQiNOok7priBT4zr
SzSw/aOWMHX7Imccjz6xJ7b1H4Vh1sK5VbdeFaIwQGO4Bj8jhSkUcmNKKK9W8PNaePWYBnSWvYhG
mQn9nDHoTo9ER3fk9EKoDLtrsFTVycisQdtXpRRX049KznDb0MlLj9MvhKhKh8CvRjLeeNS9i54y
c7B/8wl89fMHfNbSS24WWp5sMRRIdtsgacZ7TYxwnE4Qp+PbQXnskMbYIv2Utc2Vst3rq/LJjSqh
KCu6Txj9iLOD7ONGcaIr1nw2jv147GrB22DCKyDwifaxmVhrlK2SO7I/G/5oFslnukHZp0XH+aba
IbZvNcFuZc9wlhadWKLlN4KwuOdgpH0XAT98A4SjcfyVrXKt6eww7TwAGkJbm9aDik406F6YYZKB
cnX77zcz0ppH5nfhcqgVd4N29JWZDyMKQ9IQOFcqDAKWOnYpe/eJkLEM0324+5M1cuvzoHPvLFl7
U1/DPHybTR/7aa/hkzVRrg/BhEJAUS1ZHJCVQlEB0dG4JnyF627wIOlgImPc5s1OvH/3SP72vb1J
O+nltwQvavrEoQ7pK6ff8AQH/Yiajx9Hgtkcq0dkon5vYKY6Imtps6hl7PMHr+U44Y885QQR9SVy
JNC+if5k/gxdeQFsaRznak414gALjySp0AmzHigtliXAJZp4h0UmN5vGsuH9ScB3qgCZDMQO9yip
3cbBkCuyvCuOz+ZqNfQBMmmmW+Q8ccVNa7HgtF+X5ZfuAterwPx21bQkBSmcqrrOt8ZHkb/CHBzN
R2O6KzltJoaV4LpG6gIglGzAHwh+NdePOLEAYUJzm8WkTNETBkBWV5p5hdnQOyDMWc0Pt3utRuBY
7zV/3tSfCQ/G+W8gqk4sn3d1JRfioIRqMrhlcVdRfU9RJk758ci72qyaGc6b8F9cjM7Qjtqgz1nc
SxsCs3VM9Vpv0qgzAeyAumRsBLWXsFAuMtI/L+34GJSOAY2ckY9jGNVFgcwhOz+fsb306aF0bf5p
Nu9QoBcA+DDAnhw3KxHKEA9P/MdV6lmyM1iD4dk4LxRY0Dv4WEYW5CguGepHQMbPjJxMpZb8/Yfn
9Lm3Mvbs60u6e3u8WuGdx605xrJdwRHxBBA08Nexj82hMaRfGx1BT7JeDcv2lJVME7oPi/CuFFH3
v7smH7KkQaWHr69tdMKkvo/1B0bHb0TogyjnMwyAEhUXf6cY/gzMEs0XY0pUKL+qslcXa7zL1avF
whc1olcYE2usNbr54orErfl4ZS69p4e35vr/vwGU63hqGtIDEdjGXRRnfKt8lAVzEsudMZo4pyhf
+Y22xVqNZpzxTnhNBnJBbfi3jJZp4a8voobSJN3mgnLfANs1Des5GA+tIaNBiGo2ZilVgpi4Z2qN
Thteg0HboAPrmm2ofbh4+LRAU9sPG8rBVah8HxJOOoLsLw/SnWmfwCKbEK/iYGoubefjthoYFdnq
VyxUQP2RCnNPKX3u9SSHWpM1tVRwu8CL0cPWAvxazviYFUlph9Wmztah6mT/epk1rGhVhHDoDiku
wOveGJ/ayN+lqopiZ0Za9pLv/Nk1GdIv21tcivuV5ImRhAvr1L27jppwljDqIcSXozzb3nCHXWjB
5k51qn9OncrFNVEuwCV40fIEJPlLFpl8JOdl+ycLPNqeSnSDtHdVpaB2Uutg3FoDs+TqoqZKa6A2
u0RKFAyO4i8Zon2ZxGCVJyX6SpOrXVTalNz1gqOWC5G9cZ9dBDlCqmgmFm3dTeUJzCnQ0HrrjD7u
CVVh9R6gPQhaIjYze7D1e0HKHCwb0m4qMmAS8rOmU7e8ztv1cTEEbcZu5FJfPCiOxHIgCTYYpNmw
SpkoPHELMNhDNXvME2Ov54F/83+TRJnEf2cy6c4u9m0VXKCtxGC1nC6S7vYJg1sLqYdOaUAGl4SD
3WQVxX9vyoEs6O91x/Dlgtc03Eu+V/DlLt2yZIRXgpeOZ+Y8DDqbN3KNus5bztq89/BgGufayeun
Orsw0JeY2jl0LJ4KvKcVUlpIEmaiStgjzhKg419X1ZAchn6xK34Ubqhx0oRRO5YttdqleuzUW5jB
47fyOnTNLJf5uv7Uv27QIEbh3IqCtkb+yjQ3LwkR6hbPZDmTPKGk9S+YbbaJAyoo+Xn5n4Wc2t+X
eSkKUdk1faJGR7ODzFD69FPg7y6FSQre//9g6oug4lfDXdKpt+2OaeKqwu22ac7IuEilDjYJ6w4g
mpxjIdfXasyUJ/9Ldr4mbKoVZcRoMwBskJ6LuAMBQ1DfeioWuty0oOhY0LtAJQWRh2ntGbLj07P8
RJcmeudP0oTzDo9EX00ommpQQVHE43SKlha19CyoDFDouCgao74qu5+7FcJBOXbbAlVAu0HcIfd+
Zp86QtfwHIqHzqzW679VDGOQemdcK1nyIxKNKdycKGQXI3mpN0O98KqcTKRWbMo0eSIFyA1wm5Tp
+hWwgXV8gWRvHiAy+CrUkTfoXrN1hShMqAQclWv2EjHHll00yp3/IfYJM8DsYqC6MSYHy0plNQVW
JFjpsNTDS4cBt6/teGWWPUJ0xXVnRIbCubh2nXWhUqltewdK6ZrDMNSrc/GpQFHQgnkai7MoC4Gc
DHXu1Ync4bdFVR5fxnyJZ4ksCGd/fa0xMP7z6YiSMopGhUgEpiBt57nHGImeV85/r0IaaCOLutkc
9M8p1lEi5vZWvtitOF+nq/LViVtGGEuuLpRS8rY1ham+Wc6zvkFBzzlr8WCDoNIPNUwoM+HaBcAU
ZpIK6TNc03/aYFW7RhDoHXamePiag474PoWlnaZxyVkbbsDySfMMwDyaVRlQxN6Z8Z4/IksNs/1t
ncbW86cNTsv19bI9rhs4Fba6fb6V+NYDYW1OR0ficdz/cCzQR7ZVKGN1HuvhgN49g7La/tTBS+PV
3O8ljxilH1zWfpLmy9Z0Fbqh6XZNd8osPNktamwuvNqasGJqZZNO6lAMvDiMOwcsafQYusHEkt4W
KSllX2IZ1L9OcrdoS/d1b8m3MyGXsaMBnpDd10aM71M/LAcc61VxnNnTsWn9HENI8a5UfBACs7Qw
3zOCg1O1KfDnF+mNJXsOuqe1BOZqMJgJ1uT0wvnDyatCZ3DSyeWTjupRQtNnkxzy7idXUMiYUI2P
ws/8qr3JPspld6Xqa+Ai1Ysk2BwX7AnGDotCTqmggVUz94T+0qxpld4+fUe4YD2wx4Evc8I45dfb
yDWaa8XXkf46gdQOGT1xbeSx+bGcT4DDqVFdji+m6V5n5KQAdX27ioEbPLyvBqve4NNS5mRUqbX4
sRJL/D+f3ocLGwyEaSbA8zYQ7vxCseqqrR940K0SsJlDeJfv63Z2yh2dhTlxA1R1yW7FkquZ7Rqz
voruyoY1kx2fQ+8avhZLSK4l9T9iwM0hCklVcF7j5VdxzuPq1ueOmFYBwH3E/D+3gBAaLEuTiU3X
cs3ZfEq5zOGpE231OUdZ1rdk/UxvkMWxPbX9YWYZzfNZHfqLrvhzm6HPY0zaEJl++6kel12yQTIu
yHfJx8y4lw+ym5g1Asxa4TSu9zCnb3duqk3RPxDv42ZLWx87JXrBwQM4DBALYiutqu2PTwZdjLu7
fc1lrUKM40QhLLQN/SiRjIxiKmdGVV3cK7b4DlBq/OSNMSs3lD90/+tnRrPq7lWLZznq76KO5HdG
7h2oQrMyZ7nqLqGwqNcT2aBVI+3zPMvHYoyH8rHCkNMem4F+TdkSvJF35c71TTTTminYBSKXKINh
YY2LDVIsD6lRB2hGwAGfA8DwCMumbiHDmbkC9hEcXG2k8QAsSr9e2/WCJcFsFCjKvEFH4HU5HGbL
octDEXv5bPNsKmluikEF2rh2pkJs7P5S8yjI8wLHZD8HPm5WQKHyvr55Rt7Gihq+uIAVbKnFNR8b
UoEewrUOyJj6tomEi6bBq2NMeiSv3dMHxopj7LW1OLrD5Orb3LnbqrmV9b4mZz4vPYc0+B0zMVA9
+rtefwNS0yKctJQ/+jbkEr+ZGhCBVnCriGx3vXsFs7uG0n+iR+WcXvXrs+WKXetjd/GVKyhpMxXt
xZzLZhhX6dOyXsv+SKWeK3mmuLFx1yX6Rin/8VvWMTRxoVT6JAkP/nCzclCqVc5hG0PWraWIe0qe
S+tRIFTgerdjDcYNcjHORKStL5yMQrzONXmar/fxGh3rSaeC6ebf9EGeo7R22NI7lXR4iGYOwRp/
3Jk73/FnzXfx0f0RBJDN6g0tVO5rPwqLcfXeKpHRaVWMu3S/XBTuHkqethDguuao2xNJXp1MXlQf
nJzEHVlGr17gczguMQBPpHusFzr6b+usrSkU9x1/cwpJLQtxk8oA6NYJ2ww3Opprbh6/zgW60rhc
jlqHuiF9uTlVQyAMIMPf3JvT2+9tlHPzGpG4/riU8pluAxl/gqX9FZ4luUx6KnQfYxNRYwOw44HA
20i6Tisu23wpy+iVtFoxgfODv6MwNHwtAIGkuIwXPgImKnqTNZLVsUD4yyIr9St30WUmZWkr8vWD
d1lcMHx8oN/kb5W+2N0enMSpD3mv5qvSG5gTPCYAmx8MeSd/80sY0mWHUysnY6YxAh3fn8IHsITP
a5dski9QVQzzX/rBHb/+Ciy3uYcFjvtVgI5PeHCm2YnB+WxDG7IhJyia1HV2RVihv1Jd7KgtGTk1
pR8Q/VCJbfWoEqXSIl2LZwcWRwdfA+fU8Pru5f7O3kY+ubWQZVqSXZBiSS0KBgHjSNgU7o3mrT/Q
pR5A/q46dsGlme08rL9fwR9ZQETsIkMBxlM3ni89oXr6Plmkq/E+M67babgW4o97VC1H7cgysfrD
ZPPtvJ2fCnEp2v9xIoTsF6vJpA0KQln37EJfJAkQx4BXnvRghq1+yWgd9rPD0vFrvqpqqid8y2Lq
AOahtTz/v2YYHnAnAuygjrhMR12kwz4OoI/GC6ZZNjBIxbw+4ViqN2q572npX0ey+HwDsj5N7t/4
d/V9vbuQ2L5Qql9iPeup+PRY66nwTtr98kfUukeylLAnO2a86oOcIwyP2mNLsHeuFfJ34Fw9EllE
rTbYh3O+zuM3o/Geb2BTAPnXEvMTxHPl5z470n40QE0aJGcOCdV9TOAxTtH2tPjON3lFURE/Rjxl
JV+kj26ESKy1Qdz7tM3a5HkHwsT6/PSTQNq0G0ewkuVsaIm0r6nJ+QFK875DsevtfOJXcxpuXkLr
TWtjWju2Q+CkSRkip2fqf5Plfq3hkuHmB/66CM2j0HHFgo9VtSvL+nEJ5qV9iqtj/QIEsvgRqO24
wdugtvzdZqpSPoKCVNK5fEdrcNuq/KnFbEVCrRIbx3xIMjPHb/9NFQJIhtLDnUW63AfOnMb7LKVD
miQ/484iLEqHIC47fMjO9dRMSSx83UWEmZHSzqfHG8BwDJ/rNiUfOwWY+vpV2cKznV0ECzieUZfz
kpQ3NvkQQJfPPd9aJsdibS3mDglgaD2JmDhB8yJEqIqeKtVgdkJ70U7DE1b5FzbTqeQ6e89Qx2VN
XrCfSgQNXygYIfRzSGMs6JKf90o9+Cgkd08G5NfWOYf6Z80LZgZluSBNLe7Gsra37tYS7N46Mijv
+ilTxv1SCS9eazkBqbAiPCKWEUWoXzj1dt8dAT06l6xBEfDQxFIuxqBxTclYeQsAw21QXb9moKsD
OGpyzSDubI0iI7sge/aJ9JnDR3Q00KQZBEJoO7gHTyHjZhhpcIyK5Y7qXj6HAw1//yMOwmR0CXJK
vbYvQkWFT+6+kQYNaE0Pkjatc2UYpJxmb/3xMcgonqnFBDD6RDIOLEJKzrN9y4bAvC40czKmnj2v
trwF14LjR97SWphwUPRnNmpMCOVgudX6ge5GXzrUoH4wFvA5ueyMPwDu/N0sXsPM49L45ml3IbQL
N6kVYsG1N7STBZPQ8nRzIvOEJocZOd63QAGEcNBPyDIbElnmPZ5qN67O1/5HLD+RXLrn4D5iMXGf
2bI/QVFNLQgCEFrvp9dW9z9DR8tJlQKaE6WNhFfX/Sxb6XeTwtzYlNim1i4nkeTVmdwyiR9r+gft
IvBqbjGRm2uVaB6YVOyYi4W0taBxlxmks33SiJZ8TeCSLSOySg1VvxzWER9pkDNlNkiWDAeKXLQV
NFjIqXXmDZZ09+FV0oqBfkkRR+nxnxRWUV6W3WS69Ny1I1Rrbmdo51iXypO/TZZQ5kVSAoJ+LHyu
FwYx1Yxxqd6qZXfQ+yWShWqVP8B2wX40UNSSwMpW4XvKeyOOT9k/uzmTQ4SY+KDOkghiOpxVkc84
dhjXQlBG/RuH8v7JL6L6I6n+qhfK24dYJPx7+hgykqEOp+c1GEOs6kFHp2XrBC/7ZQyMSFur+E0N
6S0zHFDwDHIk7NT0znFtLN/LBm1E21gcdmJL4W3SRu7B26chv9Su36mgDSqlXkyyp5OtlkhFNhzE
cXeaKJZLOjtCGps/jq0OLPbaHbL+s1LMbGhrTMATQAHOtzg/WjBsazkGxnBNz4Zl7Z1ltT3heCYc
gYLaIAohb0WCTg3sd5Onto3ganbfP8tRxXKnCIHdA9XLp6G+R+AtHlGh3zzIzEiCFXRwMwIpvD38
GsigySX+US5FLGhsfqfvZlZCjboN/GuBLd5sOnO2lRXwsyF/6LEe4Q7NzYyVlyVFhuMFPhXY81Nr
SwmLa0MNT0cj6F3e8PLdazdTp5ODPrUmo4tFO4KCywtDnsXgqonXvmS47YuV7sxrLW4qDH66PU4d
gHmg/SXY/WRnFY5aaYq3Eh8C77l2iq/2PKzwHNvToLFgvGTMSbdH1yG3ngmoEp9TnS+y1pC120jh
4co2QpxTT6NKLUlYU/FfK+yFyniCQXRTELHeAlweLNEsP3acFR6kEnK0nkPwjMHzWzXAsUo9VLE5
X1DVI6ti8xn/OUS3xbWZkjlTX/u2jrsjRjT3lVnXTTY0ElOwIWeU6jQLjxeDou448P2fyFmX3vTu
Awz9H9oIu56vwMwFGg9b3L5kdyk8/kup+WW+0FepmrQ72NTNmzOAGYSMbWooH96mWnPKLcDSpes1
LyEyvcpJbaSuQxWuhCJls4jp1NLNzFsCZsYv6/Aa5YHDlasMWl3xgqLH6WZXtESYBYlBJ99IN5Ms
9jpXDnjABS5MCTJQmz8fhj7i5vzA55U3Yt484olGj3EZ6YLHjG41Yzo6AfnPJNZiizgnCVDTUH6r
gS0V01u1pg9HAERGn71ITv09Jx/pLSmoFiIxBLED2sTsilDgSc4HahzsA92R2GUd06cErQPtnFug
jmWMMJqCkMPCd4DJN/ma+WXAdc45LiWbmvzqxJ+dFg0kJTXZ1wCTxEEvM274vn1wKDE05NoRYJBI
s+Tdp/aCBLyyaW8L1Hagb/QnXLN4N5+Hqj4KFZCwfAV3VpFf6YfNxm1Mg52pdaLncBYF/2wvwrKa
NAQ4YrVUkqrTg3146MNdpLC0JxW6JgJnbErLC2Jp/ELO26UkYhxkRgqJEaLbZOlHaxx/ZLeyK/tG
Jb0kaGZ9VwXYHUI0SY5a04ZHBtwaL4MkVFyH4DkIRGDAe4z0UFJ8PWb7tPCNsXgOf00shEvaQErA
uvZBXXX0F6F0sJDqY2BufffdKdrKHHJGI0tvE6VJCkqInP3XXMLnFEdNRSG4XhKCD8/Y5sL5Hwfp
oZWSaZ72dBJ3LbpAyvvg/qu03dbJRpU78bltJQYdXNSenPBSCKwX4wjDYlybE7fI+ByAUf7zxyHb
kTYSfUSze+0N837kD7/F6Evh0TpqDSuRCPIdghKTFo2OWEX0i5dolyrh81VHHAxyHofS+zNhWiTh
Z8es+bEmqUEH+FXQC52xbis7W8pUtHGUT0lUUGw2S8HbtSIPW+MMJ3jbV0o1KTYVhdtIO8L1d/Nk
qhcrRggTDEEtmjAj0mPj+AKgA+WZfQwnlJiqHGYZCrCtC3O2vVbvUG6gB0tUvaB82wDJ8qY3YeG5
2Eo+2+al8sLrDoI+qgpVS36yyU/u/6TjIWXVy+xGIfQmzqE/9gPd9r9N7zgZkF2nyZFOcROsSuFn
N8cufy8yxR20OgF3JmzYEEslueCUXAj+7jpBFotD58FvcrcGIe69alswm/B4GIuvAEoBhoFz5nV2
XTlnSHq16SQNGnY9bTKgehtau2JNNfWLZUS4JHctlxLx9Da3Fw0QKDxZPeUHCLGd+qpQ1dGG+9rT
2Jjaf/uujRGVOli4NtAx95CLL+KTJYhZ7U4aRp9yJZYxrUv39NOeKKbDeUN15/caV+DG1dnUNU6P
/NrNbDzUnwKnNIkKfERq82yN1lCmje2VYXJ1HumsIcXzqYGhDpnmbH0pC5JbZl6gzA9FApAiGPDO
LYkwdmVkBh2oI5pFhTtbnjXTEIs3Eo8N9RfleS3IZ6NotXSB6oHfHJfHCUpX7soWLzai5OtIBEvv
ygLQHLd3a6N5Gsre9rhzqdK8FBi9MOPoPubI3HpZYyGI8wFvaa8+vjyYcdfkCmqfWIBVsSmVms0K
wjeGiq36PYNbdLtDJWZJUba8XVKPahOSt+RnU5kc1c4t4jlRtH8qwMMv/2ST4mVy9CjXSvUv6EHX
S7jfg0YX7QHVbkDKK8xX2dPPrjCFAxVIMPgrKwO2H1vicWqBCtARFbhPiQgJE2SkIDB3LqiaeSi6
pRcWDBo+/2Kzkgpq1agS+mzhGTjHM0NR0Ev5KLxh2petKopQzBPydygcLxoJNIJvXwS++sv8yMdX
H74xVz1Y1zo2oE4jZ48kFxsx8Jfng28J9Zk2iJvSNWU9+8uFPh+Q04z8NNIhp3EiiLiaN9NQvsrx
d8ZRjJKyzLnjZ5IFFUdfz3rYkhtg0J59FvaAfEpeAWbkLO76A3sDt82nxKYVxnW3ZcEN1ByrYH/H
or7BKO0Tv3KBwnHZowB0Lup7FNwHomLVO5IMqZeXDAKNrS7ywrmClO4iT7yb594uAlYHztwXMxzC
wstQGhkM3R4MQ1P42Ppgz8SKJ948vyzvRUmFS+TajMI5DoKkvJ59E43fJyR9/eiMMEUul0gYWeiL
A9HPdbGTZE89yEsUGhXn7EtqNrj/utRVSI3XJEKyZ5RGrzoagQc69x0TIY30oCt2WMTiXLs425EA
p7cjnXcXkqRukAu+vMQjaaK4j4hvBHelc6jXRvVWaQ8EmFW2UHnotS+3eXdgTSaMe0nyDsZo7xiu
jywL5OxghtIzj8v97fkGUcOulTyUeHEaemBGveZSKivfxbSpQ44B3AaURNHj5Sr2PXn+7SNTyb6u
1umCPzOa1KO2X2XvsH5o5Q7im8+tOtmKqWho4ZMVBW+kApOUnCbRYAmhQPm9nISwhi80lIJiiqKf
6mEfRJJBNdHsal577XcDkSaamb9KCKl3tB1IywjolJWoMAU+U4ghG/VBDj4aZcqKwCJ0PnzcpsSQ
EDkZfcH32i3uL1B1JGYgZvB4PIDBbYioBo/qIDwuUsHTGQ3hguwVYKbdS7iC2qVIUVaBaseX98lh
abQW8QJ0r4ZQBxE41IS9e5UFmED2S2AMH3P/+0KM6M/nDks7A8iyGTb9LGVkfPIb5HkZTwSxO6aR
EiZmafyQfXWcer8tx4EkpQLggGbLZwliRbbCXSzfMYSNSxACpcC8OyTGeznwNJ8EKuiAWKHa1RMP
vTRVFRYnACQw+RFVNAdATrkYC+ew76ESLbcGJbCyk+x7l90aiKfG9euGNywAtKs1p+G8rrh3wCUu
UlWtzwJRqJ2WM85mrtczkaM3QlN2j3BnGf0xi4KcFGFmKFDQ8HL8tmqTFrNywJeE6MEHEBDF5LoV
hkRrW8Wb0jbD+xae9Z2RUo1CBjH/GMOclLRqXnTDoZbh7WFFGiM0UwZ6npy1hNp6GwWw7Wi1vwN0
1tKeqRGBIyVpC/Ff6dM7L7V4fCansESEZenEluk4WkyztD8ObUjoVO3B+l0kLuhZIx/WTwDaySQ+
TbphHaN8QoNKjlu3cc2aAjBMWGhFCVM8xGCJV5sjmHFQOFdamUpXLXqecdLP6GgxnHFArE1Qm4gp
k0FpcAfmNgTlIAiC8yq6wIQANCUY29+k88EjOBq9w9yd2wVvJBWD5cEL5kDTvsN4wxJnGfbbb1ag
vRjhDi15glfaf5Ehn3/lmqBXCG1Q6mUjApTp+HQ3Q6dVHtcs3LIsRUu0rbtvYHkcTxitvVdV6tnB
QPAdmOSWxgiPIdE7kSFwMWUyi1j60D+HdOei3qwUnB3wfQS9MaQwBvsidpsqCgRPmyulIwLfZ8AM
35kLkCokxIlUQGJ9ENswdXM92Ak+SC/WZ9x6lCcc/A6LKxhNXdyoczG3MISKH6YFf9U2p86RZCoW
XmJnIAVv944FVf/wCUz0r5GqkEr+B2+0gQLaN0bOfKrDiBxSB0u5fLak0KOTCbWE/fLRm2zwZouG
dEjHocakdQB8aJ/9ZBHChQduv61LOfYdw8Eq6D7rsi/IVBvIVw/t+rZGp37yM+IJOkh0SkEIz/9r
2fpbPVpqXo6GBVRI3rRjdiUOTvWfTaiJIbYID4DPp/41U2786URWNWMxiPf7Coy4p/cQT1MCoQ5s
C8HTmqvOgj370gJoo9c502ev02C2pgus2z4mSfvr1nzdeuQDsEKTAL+f16ZzOsAhdUtelxcJN3GJ
MFkxbBQ4b2+zVtIcFHf0O+z/MlphNECdxiThDNezxKDJlXY0VR1cD4L9ZXVaU7OluMhK0YEnTKMi
OZ9/GmsjIc/EUGZrCMo67Yh9Baw9uVsg2VNpCe8r/Wbk/V1pwvEYCjsDIwQ+caG/oiokreQZcHVo
k/LOoMTUh8DJC1M4O9hALocs3KqUYS8zr8yCWi470UBJ/65eAcPt5XcptxRhQ2H37hjUyjxCXZQ3
sFJthcklqke7B2YjGV85wMpRMBbWqozPpNW82py3jL697TWMbfjI8i6sNDIaJZ+dVCg/CgUv9BQM
egyoRa/+QfYYPWMF/p5ZrmrBwlPE964fSOO19SHmeJ1yNz29AuMA+fKjUDnZ1aa1QgOwqIIWSINV
sbdEwXejGYc5MqOOVbbQTSPwrlBcU64moXwp3EwSn8x9MOKsiEaanXUnHF6HrpKOQtqrFleKJsfV
z84ETgtlCSLqy6FooDu4CAfjuQfJZ3ktE0Aswf+PJxHKga33tBJwfNlNb37J7vPKHDNj2Om1/S7/
D3fr1alLNaHnOljYd/jIoPSDCWPYO9xBMuzoXAn7qdeRwsFdQ8c4Hx8jz7e53ywFR3IC208t7XoV
7pIdXE+o7uV1ZJEpVgfQ/kkjBK+tWWljsTbaLwpys1cBNZ2GMqlM/opk6nZSOX84hJdnOU2Rjyvl
oO1Uzjp42zYeOsdLCDIxmZ7MGxkkX0qbN4E3ANsbV3BQ1tMECitgO05bCvaDKSUJGeeYPfWno36M
LBwqXQw2WJGPbMtnuwpC8UqldY2O+YfYTvqwXMsudXdx5pFxF3K4o8HJnd6CDgLHQmVZ+7OkjWBy
v08r2NTkRuEkzmpA+oEc1Jn8FvjxvQaOD2hFiPZHM64beeJrJDhythM08GtzN5OdMA8vJq39nHjU
PCEGffXgiTlkyeOhYvss1Hiy+i/WtVosInBMP3rjdk5ybRfcadS+AMsks7BLCGvu0WuChMxiBkBl
TlKga4EajW7oxySAjYNdwlN3Zwzo1uOoEGUuPgJfkXl5OJ9/FNoLCDzoSHNjTHr+aMK9RfGN1m1X
uU147s9OZDcIpHXlRwQxIaDp1KtXPT50CrPtn9EGm1ZRLQ6rMoz/gXlqiwd3KCp3WPoaAxWvIKaT
deWJBn+sY/T4KP71sX3+Lq2vHWKHQ/USnYNu9IG7kZeGI3+ILUaYwHhHE3ANFzLJN4DeE2IIo3fZ
IgrFEQJgJNBR8zruuNyHu012i7fEmxEWb4UOP+MF+SbNiSGRm27qPQhHYKNE0UGFTcflomkFkEqD
IPFXgQUcC/u1PM2zPLr0d8AHez50VbASnrPxvBwpBvtap1plgUW8O7+/W7pTlquYs/ECL9bl3so5
u4W1EtDjy6RIt2vJRjKsLxyZcKt4lvEXYIhhgrVH3FpJ1Wi+emAnXXZKxINGzXHUpULhledjhlQ3
9NTdQRyay9qIloFsx9MQ7Pgq9KNMN3L/xyNeJuwOJ4W4miTbHQi+5No2NI/J5aQhwy2N2aN6Oeum
DvDgI0FonMJKqYRVlTVOVfM56DoyKcWh8dYoqOg9tnvkJQ32ceRmwmOWubarbNUIdXpkYUJcdC08
voSdoh4yyvc6NxtmlBbCi82cK7XR2EBunuKg5pcJl/HHn/U9+Vv2l0I1UP8j+Uo3n/+7s3CIn1bo
dukEtiVcnWkuuWtualiu4SleB5a8Lg7ngM4/uPYTfjwR6b8Y/9kFgBVIBonTmd1FPby6o2ihiKqi
dd9t/SiKP+acCVDJADzjcObj5whQ4rn/2MnDwsg+WTB3JylMHzM79/XNjeoD5+oSNueBeXy+FCpC
pDZJ7DrJ9g1yFLjNKvbtvmRzEU6ePq9jh+P2blER1J/NkPzWGT/6XVhBa70I8+Lh6GC1DangcVTm
PapucSFWXKbeHBy3IJzJ6wkaXauQUZE4Uu5vcl1GPmKg9kyxEkuU85lROMFoJnHTfrsmJpc+4iNU
hAXPn5kqManhE+4svHV/j3wkYcCDBV1XCG2fubVW4Wd1iWDYMgpBryDppqS47KoVLXIvobEyEnHa
JBcqyPoFEzrWhhtzFXyB2zAuk7cEjaWqj8T7fsouazKJD+VF4kgEq3xwaQ20Au3IKR6FG0TWe2YF
J8RY9IgSy2UC17QsilU/ZnkLt24E4K1irsujmUQ2tRHlsq+NxhpeuL0mpR0AmKIEiCZGoBCS+nko
e/WOx1bhss2l5gJz7xOhT44R/o+Lz4IF5wMCBGiPaeeYWzfSrksUkVcoq17DaWixNjLrFGxg48zE
6R/oXlEwoEd7PAOL2Uo1yult+inYKTLjVF7aroDtgTW3Pq2s5CTNc98jqxNlGIvITBI7r4MhX/tP
tGVSCmIKZm6CbPxGq7Sff3ippQAb+9DcTy1Fs1ZGj4arLEMpCAiEd+Zi4PLRozCKLsPqTHbAT8VD
MADNLcCazbAUPVEWj7W93z9ZzS1qROHDpKwtXNNiiMvr1hhzKAzsq3upwyMENwaEeknJ6wrXxGyr
Ea6tjp+0L060pZ+MeFBUZYeSazYUXwzpQGj2QjpThyk130HKPfW1iUtmSKDs6jY2/tIWCDmGCSBA
REo+nPcSgUa1M40k15ZXZe1+WY1ScT22LX9Yx0T//FXFIub7OyyQTz5IX69V4u4EdmkSmamklzbA
80aFEFPC25ykivPcLLefGDPtIYBJNx8ghv8UHaUW7D9/d/NENkefFz7Qh2rTNL9oQurhsXUAwS/5
mlOQj/vyr79oPXGa8GicsWw2DAiReNzYyapn7f4dTCK9Fxw8ZjS4tvLU4T0D9TqgbtQSbvcgkL7k
00l9meyuszQooWcuhSy6aYFRMPTqGgQLWUruK0QPFGLSNDFG4rp5tttHk0nRXd1jnfjNklH5gKeT
YPFZnWu0HiGzq1Urwnij5AkUTEAeQeFMZZfGxSymEbZQuss1XUryff4i3KBNVmUxC+CWEGasCOlx
oRO1kODqSP1XoaGOEWBWE5IvTivXpaPUzRjqMZmqnc8J+r+qQfc3DujSW2beWmpKNyjNjnNKC1BV
gBAbtELzAF9OktXC0Y3z8BltX+49SFzBegcOEJK9/45FoYjR38EX+Z2gQ4TqD2oJuPyf0D0uhs8u
fos0+m5bywqePKUAVIWBB2/THb0XJeZldIAlRv7m7qYY/OWg9H1g89CeuRln9VcpO9elNAwMSb7v
45Vw5qIGijPIt7J/2pU3YyLp+tV7qIS1X9DJLHSqm3iGhsucqyHlIcP+vi1uTm+Qf9XF1iMbKVg/
9dAaEGtKVsR/W6jeUbt1jnKM1b6F22yZdtogiS0/mvkGB3pxetUtNqYMVy5DEpU0/KRZN1ucDmCt
e+9KjByMJ/fFWbfK30niCRUg9+qoYEY++YAisGX85ugPB3QDhUojKSVPcdBhPazVZc7HB055F7kL
sdQDHKKFr/eQRjtgMhQMXduElXAN3+NgZhr8EUXzVdm8pf55Bumr+vpYR9JTnV6K+nu4h8jQnfKy
lZ9q6t7I6KPQ0Kg8iYJ9OX9HHz4VT2Jg0RpMjDj35VK5eTcZdciki8p0gxS1ZX52Rcvl8Qj3RjOK
9h10M5KPAEnK3ZWCv9zQjiSA1/rqp0w2nh4yQHtfmSFNe8yCMkCSRrsiTiLKB6VRbWN8ekC5W55b
pKwT0OfwcrUYxR8hiw+tO945vAA93q55wghhU6gqZzeu4HLMfJ6GnOqiHbTfF2hb5SXprLI3vtVU
Z4ZIFX+XSOyB3vQBgZ4KcmTm45BMpiKsj4qjhMhaxTT+Z+hLMyNF/JcMuHmwkGqhF3Tmwy/ilnDc
pN5j3LXvIkYCC83ifc9i9qcisD5Zle7Ix69RJLVs5yGsZJ1zEN/bj6RmkJDlnMG7lmdVLhZ9/Wki
TJUbvjyZHjYhWpUINqBlKWCHL0q7yb2VYWNLJ1gI2CjAV7SvYcTJHgOLUzt3D87FCPvIryaikC/4
Gu92a988ioFKyhL11uxEIyg0C+baNBHK61+YHJ73j2szoMDoZ9/ihnlOH3xSD1VoNWhT82by/n4W
yklYGyukrtOoRwuy1ivYgL0vWvp5bsRoNpZv3Czl6b1+hKX2mfdCjWgkd5HIA6gX3V5Y+BLKPzgs
prMFBGlK58pLY6MNQjWTX/tMBEdTqhCvyoSPWHywo8M4rFiGubqvKopztmGlzvw9mkqHPqg7qe+p
aFV/LPwaafbzuNlIJt1oojLf8AIOffOM7C6AvYertVbW7kA7P0vTTekqa40TM9wwifGWvBAtVqno
+0zX/74e43+KJPk2+KIrTLH4ZQxM5foJkr+PgM9ce0flX+WeUHf/cllwft5J5olVUE/EwMOYhdak
Ecvm5YMeP7UEzTNFJLtVic4efK4wLkk9MlwzRAaj0y3pEyMlHAjPMmMoSGgTMe0p1hNXctSVuBA9
T3lprBMmDjyZChrnl6CKo5gnGhJXNkZkpVUQE6oUYkQnCNxKtHuHGLOYwyHrd5HZw1ukWAp31oTj
MpG2Ms9nzLRohnfqChGr3Q3oXWW8oOfsx0gotkqGFjWvsBmQQFf8uo0/FDIvgm+B1x5erJfbRoX6
lf/d7uvbeC4KpK9RerCYjxRo1TKVuffJ10mqOyqFSD7PSgaexuSFFIbR8NEjz2ZLtDRE+gPWuc3k
ES86giIf8a7GqyR5z0zAm9B+HsGkz8t4FwFJTUsZnVuQWosvL/5w2GzF62PEAMdIr05I67yLZ45h
voOMV7+kIWTpbAcSjJ8NSkmYRIkLJeU/eyy57/2lLNEvaETZ5THItCKQIM8fF7JxLGcrGcGZejOV
FO16lOQEx/TaVzQscMufgm6msuIFFXuJazUavSLyxaeh+wLAOW9GhXUbFRjm1C+t/88/lF6nccgd
nErdd96FVrmlpzXl+H8UB+ZJZPJtxxn0GuV95Tek4U+tA6oFONjPDvcxfapTCKIOQk9aZ5xenV4e
yz7NKIK439XnkuliIvn8peI8o8WFiedI3mBl2pLw2+JMokpIH4ObGVgpshcv/eh7Zn7vfPzNawST
eVF0XFGZDDRxbD1RkDjkVfeqreWRGSIGZOV8kMllEnrqvFDM36N2iLh6jGPN1W769K7UWO38xa7a
nT1Rhe+LIUeIUl5eNMjynZpN3QCtjdyUtVlzQFttFQ7ro1PJfak3ChhtVLJu+70fHIMuL1rAGVVo
cDRGbSOv2TkLtXlSUn33g6bwllUzVw0nQNWj0bHx+gNO6a3wnjgWntdfHgJdTO5l1yLuxCsVJx2i
KhxUDlqbZGJVgiSGaO4hHCr6+pG3/x/cfc0gpdaBDV1U9GQ+Gdn05HiCzOCefh9Q1t6/3N0jJ17a
QVho8VqanDG3uIeFhnzWf8AKLpGUiHd2DH8PL8Yt6K+kNwSTJyaw9mDAq3uAGPEnFBQrAs4jKsWC
ELLkPH6kptXSBB6oeoo95EM0YwdkgUTkOIB3N2iUjZxswkPm8BODpTo9oHXcLCFQU9LmicJlSohz
V8bA8z6CgGdCbn6VlMXPwE5+5vnHgWCgGvEJcBgEsXD8MIeptv9+wfbd/naoEii4cnHC4cfr+9Zd
vtHDcJfJvuhH8V2HSmuKHI37sYLN+CwVbJezM0lr7UU3Q1TTfWAQTvvO1i5tMEAL8k1FJjR6LwwT
LDcsJxXIPmyYXk6+ESa8AovoNRmsoq7E2DFF+n2BGPpR3UEJtpHpBh7C+Y1NtGaiRtQd1bBrRPoY
JXjgZgPpFokkYqzvK2VC08ofiRPp0k0NjpDBAVNcMY4T87iK/Ew7p5vDXWPzT99bWlZxhs75ymhh
PorvpRxNX/z9hRgwn66jU+EhCThu1iypLzKGSl8nPwppqHhOJYQf1P9nhmzUD7T1Crp84dvGGJ1w
uR0mvxhKv+nxlZ5Nr24qIYGQBwt7OfFxp3cefWuYWvfmkybESgkbfkr0r4pDRvWDOzmp0g1AUoBE
+Lumhhn1E1PMGv8f7M9bikAKM/6QiavOF5xgOy8cAT8Muhm8PF+JjB4SeEwYqk3t4eJBoz1HbChB
mVAb7+xAf/ZGcZM8z7ZMflm8yO0Uz7/TN3LkXDKGLnMgT5Y6bzknFUaxbxJbFyn5yGCntN9wIrPe
iHwdlluB5YIrpnB1sP3QHXreV/Wp/7l7qo5Yx9F7UmDTieaN346qinv0l38eEbdPCEzgus4VMRQl
QpZX9m4Xc47470c0JpkQxFvjBzc639+5NC8lUjz6I6tCxc3BcvkhgwfOnsZPZShUNWIQoKOw1hpz
bkiCBCh6BNlNmfrucFR1jnmZ37KneXqTdO9Qm7I3t815VNk8Afv/Tc4uJEpF9fqR5PHI6OkxbJwp
am55h1TQgUt1ykbC+puprnF1LmjZgQEscv5Y9rw+M2irRpkwjLB5OC3dnIm8nWt1irxMPPiGgbfw
5fLcl+BVFSmH1A5MKhlG/8lwI4uJ2UZrzVEvmXd/nM7zOisKKyz1ibfuBoWI0ivqNggpbxR78AFq
Ho9GsJs6fdR03pyTP6+M8f5zfeNHXmrJbtoBBx0tzvl82yvJ9/U3I3ZKG251T0yh6jRknppTZLLj
Jz556IHhtk3ypAY4MnpiOlHPN7t2UonlLOWNMPzjYwkv5KGnj0XDE7Te4sfQ3mST7irOW5i/mv14
ZT40z8doCgCKxvx/fIJES3e5V16UQz93cj/st9JN53aIuGDzx6rKdxmqvQMci4Shg6TMh3Ugu7r/
pqCnn5jSwWmOEKIklVJdD3fJwPd2HetXu/wOjt8POJxBuXB6OkHTSvfmLgaR188Unag7sEfhOBP2
k9QwiadaTDdd4ISr5bsZ35YimpctJ9f+acbrJPT/iWWv5RSKZ/2ONM+vPZjwaAw4B3IcfgPKNdup
0mKWlblfEAWaLuy3LRuxkJLzmIc+wy1IfViSBWhp7KzEseP1eHCWt3xwzUp9BsHRWh8nUCI9kNbB
n5LHRCF/CBvD4XTSpoqb01fQSeV109ASGG2l8TrUJfeRhuz/i8tiaPJ6F2mUZjR58j3hnua0ooFE
JWne04dxBKCof18ZocVpJkKo1QM19d7q61I0Zrd8MB8YOMZn+AkuRejoTQTYh4cEiCjiKirIA/pA
V3B0IqMgwZNnnm0Rl+Dlqww1Tl3YOmduSL/RNzdah/qwe/+uuKaGi/U+idZbyyjMD40pCgRSLx6b
XRdjmMDVl/wMjxuI4dG/2Dl7yyGJlCJ6s6xC3eGVVWINq8P9pzc4nDSdDUbzaMd6B0tA8b42YUrZ
26F2bxPHIGZa4PSMxHzD4udCz5DEKEAXBI4rbi6KAEzQKcUEhL+BzA9BvODQpF9WSKV0UIMkSD0Y
M36RNXvtYbNZt/3ApPrPuoCVvCvft1AKUIVJpbkZWuYUV6GvCxwZaNnyRBAA01Y7E+stA6uPe92G
JnejBjUulelgMZ78+1eHAErjjvWx6Ic/tb9jsD0FsdusmuEpb54thrykqwqhdwkK+xi+f9reJaAm
Veo5kCPT+21eNwPaunR5RZBXKtVgDuLOI3TKAX/WH3Fb10N9fQpPeDGk1peXw/8Kw8OGFbFqyabb
3ZM9CoJ/RxZRfUCDnTnz9Tq5+EkBEIP7r0mNURlwHbOp3igJrAMxffDD17l2Ufkbxu+uPOrrfFvI
vmzZ7RZ3/7Rvgv3uwqrcoZXxCSjIu0gmSLMA9kp3Li0vMrbAi4hc/q2u52esNbw4K6Bb15jNirBh
r3Zn0MiWG9IH2F18xola2OBN3YQWhtUWHD0eLLuvIhP8LkSjEh7O0mpDh11P/eboFD3MAHM8HNeS
jHajscUL9kWfmovbbpR2rQohi0h0oPGEqzacNfyHWt9HcXKKj835V3yw8i+Sdd6wdAIKniwVNz5/
qHSdm5xav+zSrHhPJt9kQ++sHdyw/snTLmUdQEBm0ERWSPvlMO72zi8eqdcAS7cvtrhq78j16Ntx
uvOV2dTJLOk8dNOAvGahln0XCU8Eyha7R7eIqwMqPxeV6vhAjA2AE0MEJHkjnv5wd1TDemISQtgb
5pkhuBwSnC6c/I9wXn+wREMhwXG5wmcCyC1Q5uCGDUgN+Kb+AicvEqcsiRKvnpk4oAyGi/qQ2CID
nq4PaldUGYPha7qyYj6aKuP8O6vb04GM27dWhPEZXLRZdm2MycBIHiyaAMxtXno0Kr5saBAT56s9
z8jZZDhrXPdPP8ZIAaS4zSDUS7iq96kSOeJWcpJ9GmhUPnbJvZ9K36PLgMO3xJLxG64+BdN5wxD+
vEmdbWZFTGPsqIFpwJMITUiLlwtQHBA8TM5jZdLQh8jZycx+pG9SKTYkTtgkNIlZzEv2gUVXv/8i
ovhS7A4bfNCrTlUTfgGcSyghgbkwjTtt5wcw6Jy+kd6g+DxH7WJOyoDXxF8gnDFLAeQDLBvR/5t6
f2oJlO7cvaoighTEOFpkemdZqmbhGpl5dzM9UK+GmTQ0r//0ixF8nSsJYh+JgTLi950T1QN6y/F/
y1MKeRZr8ne107SREXphet46Wu1nPmexVRuJSUbv1is24ZIS9WGuKS8rwsnAS/QN9BBAh6wdHKy6
Id7oosAeDZBpBrCl7cY09p3+5LILY9b/6WINk+T4zixz7cght1Y8NTiAFpevLXS+22t2+HaLdxno
CYRiVxCl874KeHJJDLqygkce4aiEmi9gZjAnSqVb493ufkHlknmQFb7b/kXJEsAsIXRrfdng/b8i
qinGIeu5K60QvZ8POUQmY/VWTEvbChdkeFTvBs/xigEml9L8UcSFh7raZzKtzbaR4r4y1cDvnZtc
MysqXF1cK64Uv/OHMhp89NxkOFodCnmlPR6iWawipxHCaWf7kZDwiMe5FInD+ey6pHDRpPEkt5Jt
aaIZND5aD67w3K4nCRGlXtAekQ30hE2pK6wB2Oah2D4gxP7pf6ZTYkLGtxnzl1K6h5ikMlxLsQRm
PpFV/3LEq5H+BzGGCsUa0OJySYofM5W3k2Aju7Yz1EnP+GTBpyR7TFjBz6znaIH5Eh4Gp1aqYn+4
fOQL3l4gD8stP0vGmzknUpDwvVM9PZdrkTlP126/XApRBXjsTdmVm8ByZNev8M8nQ/cY4rE9pOVC
DnKd/hTKRlz4gus8XiGO0pnFy3r866oXUYLB5HmbeFIao3bD9CadefG+ivVwpaljvgEb1O1p+TmO
1azMmFASBaqs3Px2+9hagm9N6zIxQZYlWpDXoMpZdiBKdOLrRFRlOnOZvUqn7C2j1qLJUJ5djjQD
WolovUOfvurJKHtX/KpA6gQFWPF0Poz/sbWXiV0lqvj0mNgHSyLQNkPKAfLSxo1oPmboFNOv9ozR
0exZF2q1lYRs+3R0VdY7lt2Ssoki46Kde+yQ07wHxI/PRZ9/17c96OdoSn1v8EMZVJ7qoSKdjVdn
6B0C4qxBEuhFw15tEW3d6l0iWA4AEFjBEmoAd9OJM2jYnVRFZjRLHwbQQdM4kqvOQiVN0SUMQfkf
ZbTUz6/80GIv67x+h2btBcjkyvNMeC6zlb/bgQhtkFJqIGhg6mt39gZZupbJlxOdk0/tFUu2o1t2
TBgq65YQ9He6jiXVhUVui2TR1t7wUCJKexPJaOGkg7BHsrote/6qZR6ED9JbOC64J6wFaQoG98wL
7FHbZSGEaxN7a9HMnSjDpNbfMliO2Hyt8rk/u2f56Y3PM5Q/KxiuJ1tf+zmHua2Zi1mkpAx0IwfU
lsm8QNxCzlmvgKrM3uKErt+cpeIS0F00jAQ6xN6zFNdhxeWcZeRx/SvXYDDgO/1oV9k3dHgrYd0n
yIMJPSljUIUAoCnMTH91NhSE/QnVCQ/b0WNrADrOfk9Q2mW5j7Wi9NwWl7dsDkgMwD6JC1rc80Kq
iO9eufuxgerYk9MSIO1VzCvRUPWdAQH5uTAMAznSKVV1dxCz1LXpd0vVTkS6aw56mrLpgmTZcYcE
YypcrGce15CMbsp739GeQBRaGPIEuD7wcYdyrMGsWgHasN+5R2dPwyvFaa0fc2IdTUnPPJNWSBLR
cdGYl6d5Aq7FhljZHO4Vhv34RiM1R6YfRi29YpQ6WkdUTluVvyeTt5nxRv1n5xTahKm/tjnKmO/M
RdOzda5nQnnn7P8ZrdxGYrIqaNGdKSu3O/rtIdWKOxVkjmz036kaiH2rFZmhJRNvPRyfkmpBtx2J
uruTtvK2mxahJbWVbisEP3DzAVK2NGoAHemyqbGjmzzl4h9OJ61v6kE+sERd3wSxirWmkSKf2hjW
8AhPZzTuhQ8tIZlXKWjZE/EwvclZ0BkrhmYEyghy1z5TuaxRvjZ+IfxyvxUQ66VcR0SIRvhYhYtc
6A8GrXQWMnm+PPsdmKn/TroUD06KzM3xJBT1Djmwv44AviMPoZk+ieTbteA3xtUcbTXWNR/gG3p3
prbsSY6QhuHAC+zn4O9l8JI6iS2Rfo8bmNm5YMrW2u10ujQhG6+Hw28vfubvLNMpphxiE3T+p/nn
Qqjpe87mqH1mgk0xCM70zSzldvJ5WO3Z6nRnseZU+4N/ZeLKM3vSffyiM5Xopy4epCYO2SfSWC7U
QLube3xZJR5sCL7psZAMhMSJO3leBewlcrYw5xEBnwltLQ891VVK984X986hzL9ZaLchWMQ9ARfh
AxIBdEWva2cLc4SEAbSXEjfWiIupw/6sHDZpQmCH4L2Mg9JZjEn9r3qWzcld9W1PFQUPShf/htyb
yab/opRp4+D0e3UWNJGYmjzpy4WHBTxvuMdR9n7P1chZbZT8FjKF4Sxvy45kHYOfIkSET1psTC/M
UXc+suxUcQidikV+zFkAu9CK3uKWNBro8ZkMyPBwZLQ+61ehxt3yRutq+Nz8gBzr37ATRxLEcEio
TaPg0+6p6uJ9wvOv6ylubBzqKi2lBvdsXHGP9GzPI+2o1ZOC2mTIrxaORP25bbGfAXCRobI3umhs
qJZKOFwUgeXR5JlkArxn4+m8rvFhZSsBBzyeoU8qtw3akHVhfVkKf+QG6MjOx3XhTVrIXksp81c0
64yLKIiu4s9aai1NdeDHDMoS7oDQjjejjljdBbAeMUTQ137BBiDdGjTSaArf1EaSH7e3pjHKLifh
uDoV67xjnJacm5CmH9HWA0s0PvGAYnr5mVIuK//GgEFaQfBjd6LZ4TB/sWEKOZnqf/iLh76RRQPA
6RxpK48+uKl/9eg8FVSgMck2XHbW/36yGQCdIXWUsEarDQa8ao54c9M6eK4QUDWPHUSghORAsoB5
fgxYMz2FEeM+u12LqO8uwagqnWKP31/OGTGBYb04K8FV7vRc1Tb2QR7CkFNZm2cN13iTRl29ggh6
Emx2S/d6RCjQtKp/gv3NYtK5Q5fhth+Y+ie5cqNBolLyal3dwqQ2lMZosL22RlwWVwYTtDNnH9fS
8LyogdEAzUocyTC5+Tpn0dZNvT7zaCo8fXn+mbmbDK8Qmfn2DbL39NkstGOt5PFU7G2dVqs7+u1m
FBjbjn+H4+ZUoE30rW1+9iN0WAO9qr32sUjR6HdIj8cyoQc9aiR8XnwO3VRS7tccjlGZWumMM1vY
p2rdF1GCx0v4PSivmO9CqAP+f8XEify1UIsB2zEYI4+CibfiWxw3jh3HcrEAfTz7UHANEmic9LQz
m24U4WCp0dQdxxmAMDlRhUQ8hGYR0bqyARpXxfEVUig8q9S0HWnz8tEtvt/ZD7U72UAi3+yoyDQ5
K/yw3Swoq1aRQ8n/ELAHfJOiUwOfDYtaBr8WTBXNweyUHXJnSx9CHQKuJ/3LbW4+QVB8P71mZGvS
d6DNG1qiZmLs3w7srQpETdC/+j35hqM0iigJDSmBp+08+AbvM29XopgdyQRlLP1BxSMgHv5xxFRg
cdSgcMVjPXJDJqJrHEB6BNyBcZ8F19Ne7qBSDIqlfNL1E/J2iZyqLJthxN9gpQKUDrBpLxwb/IxR
8g3viVzKU7uQxZG0yf6iorSvoTgmWeljykpv6XLN8tEBYsKlOFM+ZtkYQjTyKclPmFQYW7hN8wJV
htp1H04tOboh7RvsvweRF39NeiiKC9u5yK4HrKDoANSw/cF7ftPFbXiZoc176VMm7n4zOGgtnkfI
SCYo6kBOdFykJLY4gAKt4oxsUwhYPXnaHTwBw4vihc41izH0VkOkW4uU6+bNIZqYwCYaN+MrijDH
cLlOlGu1ze5Wb+C2Vr3VQSW0U2FRVjeoVk/gtF+UmEZEQhE1pc0MFLtxERNUhCrXZw+gQJnQMa7f
5fkDY7RGmS0ZpPgDEpWTLwYv6tkZmiXIJmwbSnYKvBevvcrHglzsgfAqblNH8G1tpEr8YMkBaikh
+653w5Z/2o3+1pxSYM6JhAA48oJpsDCZU2eOj/Oqj7Z8zk9osLUS/0rLCrv2y1M+DoOP0MeAJt5T
HfUw5rMHjDDtzAGh4Txjf3ygAmd8xhzDVD9nSn4hfI+Hx/9mb3ses5ajrAXUAqmjX19QD+DzxI4K
GmsczX+DdF0eEGHA1Pgzy5mVfHsT3aMewobfI4HK33BDcr6iKt1mQr+K3cikaa6dVDO2/0wRunPb
y/gONDqsDhVDsQjHqiEsWtJn4MiMVG0fpKXSTeTzYCjnPY0rJNj01AT8Lwdxp05pKqyqnca1Nhu2
m8zi1AnW0ZuhStJfbDSlc3Xc67cOXpCbEGdd0KYmVqbOKD3CLH05P0xc3IKcH5/WUuUUvGxalsQa
7MoTs8ohLKm4vIeYwjfbMVVtqdpZpMsux6NUdv1a/y/UGgFIQRxd0vejA2j/ejkEm4ueVVI/KIL5
eItKQ+vZaMIbkdbtjQ6raSea4vntYQuRoJY2lpIvZ2XFD3tcIuw4ymshFCD/h6GZM/RsJMgZsKRK
lZu4NYS/Z9XPgHC1hwCk4nvuanMFN06E7IbBGtuA1D7AYiwb6QcIVZWJN8LL+7fGi6p3NDp6FhOR
xU8tQsBCBZ+AiFmP9vfx+BbhR40DndSo6OFUGn0UbAj23w0EsxmvD8kl73VbqHyAw5SSyMuL4ow6
D2gH94ACCHGRCuzaSid478xBWb5npWmWCNI5xLxqQ5H8FX2qAJDOtOl34zPKmMLYD4nUjluMkeSt
IZfiDZWb+olAQkrWd5z63VT+TPLk8IDutb+sSde6osN7v3RZ3Shfm+Bj7kddRP8uq2Nta+KbnToR
CIQBw2Ld6VcTNfhD4OvTL1BVx9tdG9t56OXm+UmBiEjWA4Vk3v1a4eXtVNnsBeSfpzSGMbHkzO5d
+l6/0gn1l606mxq9FLssKR0NCcjW4Nv34+WpOh+jSdKfkjVMr0BMmZBFfr7avOqRtxmRvRz5fgd3
a8zy5E5iTzYdz5RuOGbDfWbNU4BERZGZOnY9UFxG7RXN0YtdDyMjVdj49jnaKNLadiu0DdoD3Hhf
KGe+dH4PHaOr2Yowlw16AAM5dim+aYP40S51NsbToq28E97RyEGs5cxDDdj1B7+OU2ygWFTXr38c
GKoEvW5w3aCnMjW9CLSRpIySFU4AkJ2RIEC4jF02KnvVbV9ym0m3yJhakOgHl8b12GgxKG8k0xcr
gPYalsxwcGc0Q4hKmrxW99esa4JlvO33XHVab8U80f3oWs2eyEwnd+Wib0FoNhjzM5EiGkpc4s3U
IsPaib4KwSSHkN+9KcM05oNZ1qsGE8araOADshqdCu1R56DKFcR9Bvd5r9Fa8U943Qpp/AUap9WD
vp58oAW6oVtuo3VoLr36WXnwlVz73alu7zoj18KnEuM/FtvyCfofKFA2rwZhWjd3/2tTi64Svt/d
vgh0MMw/ydcIYYPKgYPhXqjY3Ye3ybk6YHVqooxvEvhMnh90NdMaY42dd/344shQ8D7sNxa1Ezjk
djZ/QAFjigy+8/REDko1IU0H4yDdtZM2cGYUGFGpg+CB0dUYY0OcvsEVWIBnkSRL3e742FDct0qp
Wsugv+DMvbnn84Rkl8QJOPv7TatRbq98l4COpp1Rsrx4sQ601nCV693Mzn3uQmkE2RimCdMYMAD0
3GVBtC8qyRVT+xYRYsrLajINJUKKnH6i/PtJPyz6JCVx4Sx2taFqDFyyTZ06n1ewpRUu3DKlPdpA
79EiJMHUuN0mfrDNEVTK2omcTLDNqrWf9pplSnB1B7JXrwdkC1O7rZCNTgx//78yM4dMhN7mpQ81
O0UYcie3p/6gGcYr29of04QaZ7LfeAhbxkSvqmqgcamJwRyVzCFlnlzto3rTCBjACU0MKYLyeEGF
FqGwgxKMM7iTBF1mgqoYQhMRbGn4xfWvuBiCVqne3tbdQYhPyVX8gkJKfY/8CP4dFvrmYOWFRtue
A87PgeUIVxsOka/X7RsJ4AYEWrI38tsAlSaaiVJ9AEkThEnQI2IpzB0PyD5IitVQwz8pz9VY6rDi
2LdcwyQMlgucjGtoim1soRgRMfzMn0pfSI6DA6Xwv1PDgcYU06++OzE+zVsBmoivkwlOZKhZVfOq
92HdJA1kfIQFXbQyeVYjoueCnuFUKhwZWQlYkB5lprOYWQcaskq53W/AHecrSEIHL3p+QBnogKWs
m7Sckc+rt1qhWxV9E9aKU8pqiMERbqSrmYX1Nf5XPfiqm/OZiMGx4Cn3Lc9sK839FyMjxL69tmgQ
dbiYMB3HrF3mQxJyd1M/YkA7qGApSlgZxn+BMcO42JM9mw8HLH5peK+ukANBA6094lgFyopRy5s4
BxqUwMzPIzs3LV/dwmyR1c9lqzMN2uHHoFu+RuSIxb0fX/WA879WEBeQN5yLM8gXXBrf8eVBy7pO
DLMMOu5RYbhsaagIPBZLDJGmYwy9OuUnKgZwjeWlcdEsdinHJEnigRp6otrcgMD4Uni339YLfofH
Zs6cdb5yBQ+R8UhgdZjMTKY+6GRkdHetAT4dDiyawUMSZoSTJ/3qHQgA5C0podShzFrwW4ChzCpX
vcCPJkyUt52RKbHFUV49hx+Gc9ZM+0fbW8EBSe7AkFXR5PQHfD1iPhPSg8rXkjsLu67YM9D+QIqj
SKu/LasioWA/wpk0Sw9UVf9YH6i0QxAB2RUzXUccyuSfcN2gpT78GbX2KJ/u3YjKBcLJC6Ykl3B3
dp+Egn9f8TL++dX7pYSzhGTfXzb0MrQFAO/tP4j/uOnHRvQyYScFWJ233vZDbIkbAohSeGLJmD/D
lIpmzrv+a3ULLM8HCl30BW6Ffepcr2VRvAHRBp1agx9VyB57fr4QPdMsa1meiAaGCRIIT0CTr9Ij
eBqT1k28MMOrX5A4XKOzEfOjHtsHofRYe3TrGeS5WtZA4NRkZwHhRJgWn/JqUJeXNajhEh7RMtsg
V5wkAQxo68fqCmbPn0aM7ayvpF3sO8xThkd20CuCK48hJolC4QxU3+WvLBo/aQbw+kSO9Mi2OaS8
I6xacjYyjZL7U8EqUfhnjbEYdeEWpM44NB5AnubKmlQx51JSuATG/c4Qx5kwtxNEmQinQu8bBc+J
WIoJBWpRcbcpNVd4Ugq7He0mpiWsykCa/KPjv2CueGi6kO8+HIBDhRnVZye4zNjo7eGUc1Wrk2jM
NGgwRCQdrCLWYtbJdzqmEXeFMjgzsAriFGjBrLfRN7OybDiHpwMryqPwfRVR+Ta0/4KI4MU7W715
9vdNJk45FhhZThv7sYg6cWgNZ/ZEiY3TAjg8xPWOQliIp3fvut/ViHNgAEbc5fPyuKOxvz6QXzSW
Is0KjbN5WRsLQl8Z2FNAvenp+tBFPNyiVZnErHavbIAXL3mkVX7jXidLjAMfMr6SPPzG/feg/1z3
Xd5LAqYoZVn7msGVgOQpCU3vkv/mtxzGL1SnuFrsEy3CNVzHIm/Rb4/6P6BXAKBi2WpagqQhAPkS
p2l90RQM6Q7yIY+F3+Gi4mk4p2KE99iPe9P4/+0numunKPGzm3dnGkYgbuxeIf9uDC1Bhb/CLcKE
dyDIoWx+Y38+JQerFDBREwThgBHvx+AbN4nUboRJAQzuK2+LfA2wjdBq7zvqH3lkwmWbw8g8+1im
K7fnDzZP8P1e4sNkDy9Q46LIEBqAWw5T3vlMFxEI9PJbW+Ex6aHXYjqkqSfVVeRX3o1C7y+CfZUD
zvVrlTYt+Sx6/tCUpZVEF+JJWbmC4gXDEfT2vdAfm1QcV7bieKDJOD/8+VIqrKXuhzn/CbLQuaFz
4VwpV5r2BmJ51sn+sEB9UtlzFnO+GXwmvWKQEhAmSiLo/FZ8s615UMiCLwQNsFy6uT2HG4gzsgOk
RCw9FdP2AI2uLBb5WkySLzw2J8WwG/KEuigvEnBxLGU/VHkGarsuu20iclVn1vkTVvZVat6qEnV5
YPxISszMpI08F+bTDN0AMbCVSW8pXJB51qdwfzhvHXwK1G6arTaBSTLORRO9bjKgwLtSnk5SOmBN
ekrebRzhD7rxn/Wemf3xC9Wv9WMi7NDcBiDsgWfN41Ii9nf2PedsYeoWX3t4NTTjCPE2T23A62jD
CuB0LZPfH92jzZg7+9CV41uxTw8rsgHLSefA1ZWvV8P5O6j1VZ1tTqsHVadlHR27Q8r+7wNNeOKs
/UMc2pWU2Kti4JzptyQGb+H1uid9YjZJfoz1hosle/C4mTdsCyW3e0MouS71QOXr2ECH0zg22Xny
E+U4il1bMb2TyHVlLZvj0vFQTMTjxwla14bT+VAQ2bBcX/cqVwDyBgdjU/Gjw2E2W7rcoLHwuN4/
FDl7fIrjaZ+H03j8DOpCdkZmf6clzK74Zu1gfRI9ioTcq1yuyabC45dwkLfvWBmTrBcdFN3ONH85
OstuNnKrwduionbhWljMN751E+qchFH22VE5IFSl1/Lsd1EQWUGquUoMTQlOgepd2kOZZMC0jZg3
60GmVbijgAwVr7YlmnFPW7XXMP72GGXkbOXClVRNJVVRQqNL6EPj4YwRiq8wTXzePcqaJJJ1aGE6
5RahvvjjZgBIc1XB6rtRzqs1koz5YTj84p8hr0qgbAuVSmbhqscu9stqqHeho3x4SHK9NrMqyy9T
fUG87IJWGUocr2IJA+5ZD1N6cxack9VemMgbC130iX9nFEc1N3QZ4ok1WVJwlh4HdfwJWEZcW03+
lV/8wRKacBtfrav6rc1l+R+Z1Tj+EBRoRwnUbHNF+FuQGUx9Dtd2oYTVHV6ENPVjgYVYO17OfOZk
vWRLZw+Mhaz8Te3eOnozPQsDjnNTN3rWhO+OQk0LrE78bmo2PlyLpf4Wz5y8wgut8QHx4fGTjUkv
xkq3XeFwHG+iCvqQqVzP8db2mfgNhP55lEUuENw8oyku3EjClAaMfG67KGge/kuxYG+siZgkoHqF
dAYc73FfolpQ/X9Mmw57yHrW7odQ5gjvTj5IcWWTpi8ya430T6x2At8g2sGFgy40s/SIHQhCSfGZ
k38npms2BVDvrUkhdnsNcLfGSEb8Yu+dLajWrxOxhQRfHVe58TDFTAk7op2PeIYTMuwguMAV7Qc3
z16xGN/loz1MqaOSZ2jzJ5JSEHFZrzhD3ORFOJKP2FeF2hNLcbXE5AIcxa8GuasSdrgQMayH+xLO
jozn+qYrmwsNnxacTvbTO2+Oo9he3dBn7m24IE85MUaEMCr6pgt7QLq52Q4gOIh1/hrSVfOK9SHJ
gibyhYTS6Rxj+uSXuAHA2oZEhlhlxNTPkjjX2wDilE+gx/h82wahD0iKrJsPimIr6Dut9CrTrNjZ
ckA/6XOCBjp1JHmcnWqlvFM9H37UvGEfhrHay4mKhRuPGuIYaSm20f/QCNC9iirH+YNBBYVZC0Tz
I0IOhYmzyQY6yQB7m/IdRGvYFu+/tRRsMKWx+bD/kEQJ+AWFQX2KP60FAWXGr093tPcMwvciAR4z
zfe+cPcTVhwZzSPFq5ugKufPRGWPB8P1pRRtIALXg1r0UwpDhj87ySl5rDDqlEw5paykdFCgnFYw
pCMphN6POQgBPhP4l5MqX/wLQdrV4TbmhngPxmtoQbYrjMirEj5O1ABTTPzueTYDRzWvW8CmwAO4
t19DMZLGOp2WiTIlMuXZDu67/G/wMlcR97MOWIFeQWimH5rFXyPOf6zuAEv+24fqUlwwjjCCimgR
3KnybA+FQeu3euYt0lA9FINF6Xqah/VPqNw9ne1OH6MoeiYl1ZjYHnbk5j28AdSUqKAR8JwsQN6u
r0sAI0f2ECArw8hs882mLVyyPymp3Jo3BYqQT3pkYH9Eo0xvz4h6UwN4P4fUOSJqTreP/92ebeuW
LeaLPE09C4rN1fGKjSSXRXQP54dlpZ4bkfpd6RPrzeR8FWyBvCcBkbB8tfEzF6mhAsjgLmJV7rXS
SGbhfOQfI1lafHN7PKqal3h5HXeA8kWmnDlnsdT8lhs52Kino43BHsWW2DIc7K0ybPNMkcw9p1fe
36EO/W3X9JzPm3g3iPgIGQ9UIVWjGj+Qw5keDjQgrXcTJjwPs3i1V/VbMEf8MOWgYDxdgjoYfS8f
hgfHLxE+Z48AjR40m11yoztS8o0mUJ4Tb/7Ivn4GLdOvMAyTf655GWqpTWR7Ht4gO6ujVI1x6H1f
rloE3lOLfJ+MjbADRFCQNvH7VNRhH2K06QcLQ2MO9CuexL2aM+nMKh5uv6cZdG72+VadqEoAUSpX
xb7Xl55Cg4ChSFI63lFVZ2SPecB1gT+gW3GoBZZ4OTIqxjNW9tOyZg1Nb08yeUoSOgSWKKgOks39
ZypTJBaUWHVQMowtSF0M50nPNl6eOOCJsDrZgZQlWFnxf6fIM8ZVKY0J1Vegvisb3ea4UFU8bKIN
Sp+d3QcDYjnixzg3HySBOp0WwDaCos1kC5GV1B53aG2s3ooeZcb8JLO2GDEvnUlt4pcCZsiuEyWX
qZUHC+2Yjo76tYTcJ2dy5oMps9moI7420+rLR15Cc3OnIjqXiC7ttF1FRetjZ0JIjt/LKj63u9NQ
h6Nka0nOVBFJevfdire5N+PINkE31RKtJe3L6ygQLyGMnap3VWLA9YMzRXygF7r2CrgOZmc1YZh+
4W2+yeF0UBCLqOELZOwEEuopBavYrpFoOS1/FZf36N2cFCAFkq44mOXOoOUEZFuMk2GW92LZYcAb
nqIW40CjIZMEifsaMomlXzS5QkaXd60AKW1lo0/lvwct3K+DFF7M/TAuu6PR9zY6mMr46X/uL7kt
DP5vCOh0MCjE5oR7oDXf8pss8RikrVMJ5feyWY9LIKuwy1YlTyvG7xEYmmgX5tjyeXffQaoz+vfM
YUMgyG5OKzrk+vE6CRdr7OgdEYlIoeJj4YTFwY+Oeh9rhWu9EVNt+3kMD2vku29T5y4gGr8vhR9g
Dmuj7EOivn+fjO5VnWPdoGBhhCh4OW9PyeW/RQwwDKQaeI1z1QhYjFKbEGK6Cxa6J2GnKI/Ncfuv
fCK61HELpvcyGjMg7nYd8HxIBI3rSr8/aqhWbbeFJkB6wUE6het1SpPogQnlCw1GKB7ENHVrRU7Y
VP0aUsCjP/xFu2crpCfS3xRyDtwb13VJP/wHeHmBpaCm6WIDTArC/XzfknkM6C4QxPGqetRADrIM
EWtA9QK7pZLzdUJo6y9VUKkDiuiYg09/GWEvYNq+JFCl2gGiezzqgG06A4vomC6ymRGWNHnIHcBu
WyaalqBn++RcFyOkgTJvwBU6g2/ab0cQKrlgrCUAZEuoNoVzY5w2ncj58WwHGRllk4Jb2Llpx1M0
j80ou96gaOgKVpZLlW2Tltd7kS9l8qjUnb4uvVUJqB/Qd8WHJmyHipI4fCdF1rD0b/SjqG+a6SAR
ZyjVivSMqshxB6jYoDpQmpiZcDdiw2ltJYcvfvUc05DFM9mBeynspaXOO9/lcPwEQIjET/6w0Mdm
U6fU35vTU/Pao/MVlgBUGOzhusBURPlgHdn/fIfYNnowhdHydjLfNAUak6pLapsTyVAX4SjUkQxD
JuEadJN7lqgL3u2uruFMi2LIPOeTKbrLVdtzGrLwkno1peZLphx27uhMT1efIjo4wiGie3gncOAX
Qg5BFIkmfFYc6bwBPQjxiSfZwANUZzLUkC6vSQBRtbH03oHxlrfg/EqcP3iH7mftcKWB7EP+XhdZ
57ySYkHF8zcDqf403szOMZJwbYjHAP94VQQV8o/fy3I0UnUUZVsoXq5C9AlE1CcF8Q3aaK6+CZqD
Hj41wcSRLffqgN0zMrYq18k0eFWGZhZYCShgd6vX+4t/lnuAqXUICGIBNaoOUL0A9zqX8d0QeDgZ
WDCTDw9Wzrp+LIGwQ5mUcbG1jCneXJFwLhbCmoejbDiqa5yFlPuMxXnsdCHNhKifYdL2i4PQPVMR
QM/tXZeEq2SqnbwljA37IBPUNLmGua4mO0RvCFJ9dpgw3QJrEcmq1lV4pXtgu/LGDrsTWRv9D0JW
g7z6l338JoP45daRotucirhacQTMKWz5tACAaqu5C3g2xA6cDQWcRFhonhMRXjJjt2VLjVpCUtFI
C4AC2cqvLMamlBlFuR5J3Tj3j1ibEIjVQWJpFX3hxBnl3MLCiZkNR+RJdb7uaqGfxToHI5i/iscf
N9HMHNSENYG/ZTbNB195liHzHh8Fz7HDfYWxldfqgFMj8Qr2klXzudzFKalXSW3+Bn/IHCuSRSVr
TPCIN2mhWEMIgIDmj0fwylm4/mXFxDghFwlQrfANXetjkcuuzMHd9MxUZ+bIdhD/BKW1+Jg5wx9N
wLRde6l3zTGBTlF7oOKNuojG0McLDvG4aD8mVkINZluBFeR+dw1YFc8mFTxFn850cQQgzhlYpvaB
MNK3Wa0JbBotXdV7v1HVhUt7UwXfaIsi700756AjMXm3W7QicE6pcO5r48W6lI9p5AcoaxOy37B4
7gwrSRgiwZxKXk5GFsAwU6NDWT+4ooBya5Z/6NWiIlgAjGSDTJt/lR5tgRbYZ4jcP/mfzniyQFQT
VKV7+B5BZOYA0HbT8qNzXiKhPL+yMlgEyMEaBDSp8H+FPtBYDeOa1oMO4P5Mdvmb72y7DdKTr3uU
5nsarc7uOKdMCBK1qZm6VnOTIrDuWUSLbdE8Or3pmDoKX1jh7CJPTcu6PpnslCIrp8Q4IF/NZGZV
Wxmf2C1tbQU3u0BhACxefcYdqtN5tcUgNNineOFzFavHYSu3oq9Hodfc4rGl7BzzFIwLjk5LuQlJ
YHf2d7tKOzeqUhTBFOxRGydmqYO+0yirJTGbd7Vzjo8RFi+9pQrSf6UBaGy8h2o0lvTtKFhzj9kb
BBCXVCqhQV1TS8NRoeojVUM86k2Bg7+C1bighnXDf6ROdQMsg8ILQyHdhbTB8CO0L5cHSYZ5PrFL
HWM+E0lKH3+jLWvwvVx7f/nA++XvoC6eZaBe2jVNir8bP5AI4h3+KgiJAao80VCb4yFPANfZjBLp
W6bPIl9GeEPxCzgWWb6sEjYSNywDwE4j1g4nxENHltmaNml2OTkuPL1vkekraE6sisiTWeqR6/TP
7fUBCMI4/jjaSt8eRKCVesKifm3T7XMbbdjI9PNmN4q9rs/SZzC4dkUlt/CDeA9nbtq7TLNxaotM
rI4TX0IFf2O52TBA6Dn8lSJTZm2oReacNiXBrN+zYP/b8pFPswZcj6HWOkWyeP1H1XnkYo94yDB7
VoSNJHx4vQOshCZYFG+gzp2yXFNA6mG0qAgEyPZyFDNcifJ7LaD8+g4BMBbRWfvdWe1O3a0isTzu
nJZAZ6uIAt7noxcmcSWqqvyLmdB2QsUv+OznkdCzCiustF5eK3kxWfLoRrlb+jGQ4kxv9jzUQAe7
gvIJ+Aqy8ydCnirN86ooiiiMqrP5TNkyg7nuF6/3T57INZO9zf/KN+Y+CoZfds9cf+HwJi54wSSn
dXk4B+PxowTcuHkcEaZUnF/3/DuSEi0aH/oAyIqUa8ACWKYHe5zaybH/ctuo4wJltikdxzSj+EeZ
lza7TAecTkYI98aBlJJgBefvEtiQxu4oMIls8MTdEg90B0tFx3KXEz29slyjqibhjRxkQArL7MOh
ATHhBt7RlG7uC89N8UG5l/2pkxYKgcU2NcFh9YPlLfq+U+Ux4r8xlLhcxaCGeHo5jXXf4/kO3WLw
/40tRY9B2sdxFGpVHYVRK/YlIUlBA+venHePunW/GVDU7zIbtw67opAGjGjDGih7BEfb6585qRof
FKk/4ivMMS8+0vDX6U0rcdxaP6DdTuKBUb/BH/sMEwZTYDTVk+2FU5SpfVAI4a95u2NAF0/hNMXD
TlPqTCMCtsS/NauosC35vD8Hf91M/R4NMMdWJxx+d9DYRfDGy8bsj9g2+FUNz6kytZ4jtfuTQxLB
oTEAdYVs1I0rZjENF93SDIAMl+AzWHjzIwphIfccDbGHDJ4YUj0Qq25uii53nx6bHC80q8Z73oVd
RqXX0FAsb03D5JuSxZymQV+1WnHdg1iUSf/cIS2FDvSECGBL3Huk7XPktKhmpPfXbtlme5kzyKB0
dktqnRjzOcDmTVhKVF7LrPvS5YGFN1u5vAnc0qFgLLfRQFCRsfJAmdAIYQkPm4otkeZ2rLFx1Ic1
FtI7y3egKAxMMKGgG1VLokJFw8+BEKcg3eKMxR9gi01xozOr3VISCu8Umf6mb/Z8h1jnb4Q/vreR
AZda2vvcWRGw1VKTGnzuW0/XkpUHFqQfpAPRQCsHbL2vfilzl+mmSlS0iM7PPsnb0jwjT7IRHCv8
DcCK5oHIQCDsTD/p6aOLZyejoHgShMPvPFvK8oMkiSfYhzq3AfDJQH0WegOxap0CTJgCMr4ynmb5
YNvdj86eRORHs4zo7gq6GkoMy5wIIV3dZWElIz7z4kfrTw6hPS6W8Ormy4WA/6cywia7qt2tllXB
KPTKzuvn0eqzAkhzNwBZ5KCv/1wk1GKWJzgM8Wv+NOIWMNb2Bor7V40pVhfWpLCTh3GSx6VCIPut
5BXJ4JqGmUcPK2c0wZq5UWF+qZLTT/6TWnQ02sKEybfawDKRZYZl3N5LpMAnCCwtrElHA5b4GNiS
rTlFOXWBmF/x+r9eVQsu8qvjlcVp3grzX1E8kO+bM36ttFgLin8/7f1FBe9fS1eNPcsyhnKYycMb
o0KQao1CzboXEJ3jx5uYWlxlvBz3PGCSLq5NTNfDLR7V4ENgomsd5MEz1RqmjkLtMZrlpBSZlqM0
GviZpjWj6riV4fAqtZ46Z5FA4bcKXmeG02dvhSmBJZ9jWggT6anxycibKQnVhVnLlV+unZTKfZJw
FO6epCiugvvAEcLbNEv2VwY/g2WPC8C4SCWIHfpf2XlOaY7dQqNICPmu2EiwFeYoLQMN/CCvCWpU
5SR+bNC56Rzs9rK4Mm1vo4igNswwdb6FysooE4Zl4WLZh4t4VgZcWJMIuC2UN1gJAk500nIa67/g
Ltvb9hHAhLhL1PW2itqxwqUaZ4jAARhpHPkjGFJLgFaTqN9bxwzq7gQVfJcikVbYsypjU1bqdg0g
0tZzTMhsJff9mQwWhlOOwX8/8V28ZTbc8YyQ+XY8FNYRZzUih4YUwQGFdb16coiyqTGCJaH0Wdoe
MXEE2VF987OqTWx7XBiv1RdneKdRaQFiPlRNgIdpSmRe8SXDabzdPFzGzYp68uDj9mHsqyWY3ETn
vivYP5RjlLlK9FO5YFSdqyWzlL+yWcMy3UdehpmVTbwx955RjftRjWEGX99XgPK8mCauI5IkmqyC
/8rZgF0oEdXVOkxSZoE9Z242Wb2UuDEnglLmJqJuTYmU962BMFa9KPW5gyS1Fnak0s+VaVwTkjS8
6AZy5Sz8DNNtqR5yuM25Hce4MxRS5Fjy84fBiHvVKFPNNGCKx+lQWV7vD0xnomqkjpL53vhT4aIf
GMmXVPSfB+VyFMLYbKaA5LrOkmUF3Ral6Rxj6ed0CJwkewDBOfXXTVFFYmIjqhO2XIjRPjNGQxeK
OqoHzROcS+W8sxoUrE44MFaJVeh1AhFTz/OS8qBAoDN96iRKPGao6h7mBCZMU7MU6TmunwYn8IKm
zLBs+tFdjvQvTVHqQSnIRWQesaN62zodcztC8GzdaorNoRXZ11JAQWe0mlTgfjzb/WXFtMeCbq53
Ic055gf//Ns62a4/WOvQMCkBMu4brbCrBz8wHAVDU+ecH1+cRebQAq8gqCE4I1uNi5m9vPH7HgIG
QidxMtoA/He5Gexi31oGfE4/in9TCmfufy7u8MOjxAdXmI0otwJo+J64Jw1o0tNYwhtNrVWRE+s+
eBeHYdG+67oGTrW9iob33rvfTQY6mJVTN87KKX/KHcxg6QD6eDp3WFNjJo+zafApw08s9TD+vLRA
u4BfZLVYSYqY8lC4+grUkbP4xkNwrI2nQLKqA8iNHVdeKdSB1T2Y0uaMF1l+wloPYCSd3iloNfSJ
1u0HirM9emvKIJ7Q2v/inWAelJPrN8Mra5mtUlWiJlmQuNqBLkBqzuDW87o/iPuAZv5ikS9rr7gF
bilbQjbhjHoOB61AAziWa0LT7IHFkd3HzN3YNnFEIAtLjQTgdyfRYTY/oMHHDZbXU3O/IPg50hbF
UNIvt+akAy2JtTcnGwqBxgnCGNP1f308WcKSbpUE0fpTLHU65m9+2VZoua5baX2GB//d3AdOYcbu
wkqFk7GlwU3Hf+OZ7iYf2KSkE2h39AsimsTPPqY3R2POGLO4nsIOToBSBhmoeFRGtWa3GPin9a3x
mSvtxZs+T2OIsVRjv1Mj5A0BwBNxK4dEGUHIjuT2DpHPOtNLaA2jHU0qpBiw9hGSsdaYbpydzu9o
l+b2qU0vKCaYnSWHdAu6lbGixD+RRE+18k4A+P5e/GwFi2WA2L19SHFZoRx5aDvowwhUe75eRdQj
jLm5uzeUFA7/Z7CErjS9fNKOyN2KjShG5ksx3aHUNU9j4TfiW9uT0d+qe2bkBnMffr6s/pQ7yxoU
2l9uRf+YFyR5knb+B0JHsvAxJ9t+91PZROV18UFgXfHunwHfihLzhh6h+u8rQuHd4sHLHD+MZCSC
mQ1qxL+6Gxb7dyC9AgttEtqpPbSidg3GtdmL3nV0CXx9A/aBZwzwqFYiNYnZkgkwXKNcyyWZSn1P
M4vdBkhOGNiBitIgdqz1lyEQDTgJs7qu4koQ6LfufMCdJqmGsDN+PTutgMowTxSBP6dPAnZFuHKV
ZaEZDV0wtI7TIas4YD0bCxK/9lLtAmYebOkyTt5QNXu7n/6ho3W79qJfcoCvhujGEQaKPeRSWHMl
iA54X7j7Ukd9/H1CrX90Fvu/Bgu6dj8EcvDGjhaFkUgf6MCeJH1tDpY9XXWAGJiIeubdJmxkZkcR
79rt5Ct22ng5nJl/Uuw3vi+fRQSxumAWyb8C+liaSg9HL+bM6cULcNmMHnBhFXK5pTKirUXvjwy9
XqmOOb8H0w6TXydwLSHyVhySYjm8lzLEIXwuT7NfTZPrbQzl0p1Je14UmGnnUIjFE2GUyDJKV0pI
Tel2KGNDCcpMdXVbJmP59HIicBfBL/8K8EhTfIVIk2POnXiODPAv+BE1tm2TqQqtIubejiknct8B
TQFJXw1f4OG72HSwq/qdCQbk2NHWn28sR0KvJeP4aTVz2K4aW7HBsWdGBhTlEiwRzqRouWwM8SQy
hAusmRVPvCsbqSthC36njIaVp4GNzi7qF0rcCba4BGf3vQgiCSqUovX/csinIAGa+hFB806xE2rD
cehEEfEfED/34f1oediyByBkFw4efMZmQWElRtqJrJQstMUzok7NC1cTPvbM88KIiUvRJc8LvR2T
FgVRk6ILlT6k7eFh5+hY7YyNtOlZfr3EIw30nY/RoPWqf/aMKeyUfVlvuWQsP1efCG/5oBWK7yyn
fzhnG4QF2dqu8ONP4fOs5JucQcsM7C3+pZ+q9S/tfXqNixEU/IJOkQRUaydSsByfzeEOpGd98nPE
tEsmunK8myJuSUPYdRfnR3I/spV1SDPIxAQkcfltU1mDon9uLBDiZ4ENMhNbCaLvgAMRd+bLApJa
x3qNYxLK2EUv/yHAd949iHHluiQyOt9VtEXZLR9dD+dj+qodVZKgA8VmkyjLLkfMhj0qaZbSF0FO
BiPVZ0jH+xGU4KTem+ovqm+r8nFrd4cyY2+65BWEnSG9dJIunES9I2d0B+8W9E5d2YG2Z9i8dDZd
mF6imcnC7fk1R99Ulw7vjpYynX/r49gm498FxHAk9B1qcFIqIz7MjqLO2PfLbIw0YjODgLP6gctQ
h9+K5yBeiYNgo4Btg9sS2xuR0CRklDhzjVQMiDqFapL6mFJeUsahmlo27CD2CD/th7Oao9NibUl9
RjyNe7tbSyyzNjXw/RxNQ9XekfqHrzlJPdhbHsJcZRTsNNm2C+HM8Dd2zR4qmbzpRm0ngIR+VWgG
2QgVYmQ99wOGiZ4fYq4LvQkt8rrTGtUVSb0i+odY/sRv93snxrlXogyuPRcwNeG7JaeNyiUjxGvX
B29aXMRHQuELRoOSU1ezpCK1H6B4evaR2lQHhgou3sdTk8iWkMj4WzF/MzVf68zs0tM9T+uL+xjz
Kd9NMnIaTlhK8TiuJDPmY/nghZLzrAJI+W6Pe4wiQ3Qmv+h2BITpDm9GW3za7X/DCbhtgv87mrs8
JxcP6IaYbQKWM3gsiHh3rn2CpaPBoouaa3MVrDDQnAMeZTO2YnF2PB6OwZ8NYB3hwUGufoAUF6gj
P2tPOn2uI6L7OUmUoeMD0l8hVNZRd7OeRENJa9rNbQJ9G4qNBJznoTeSJV/2TJdO1tNxICXHQz2X
NNONL3BTcSzJbS8tAIB4YwrIYBd3eK0gOM0CXZoNqtguYDxzOgYUiLmT0hPU+TAYh3rVE4Pr+oxB
v7MfTZ7PfDojgcumUEgwjSQKAZXcwBnLDeurPOgUzSR7lU038nN/AMk9FKHn64ynn/mNoROTp01z
bTqVN4F6QwkWNvDY6reCAd4WPj/ujRjcDuB9W4Q7AJq684UFNKXfSFt8wtBVNNl5nQ9ME6T9HpL8
cwShJRuvW7nPwrZwRFJ6keTHzF8l6tCG7buyfRYnn5Tnwzs7im/0uXRJJsCuGTsSy4G7CPo9gtTP
c+96tTpiVmpAQ+LJjqy54+sMqM1i5MCPkhQswrKO59Dnge0N8E9FMSdgYkDYk6nW8Pa3aKfL6K3L
YtbnMRlGhVqA4g05OXprKJ9YyWZQ/UQkC0ZYgRcu8NRAc6qQQ8023l/wzAkJag84bRAPuoZYMwWf
pX6TFQQGYn8yk1vIuFq426KwQ8SWO55mBeql+chp4ejREa/4BHnFzxsSh7HJrsRuGu84QmgxXT5T
jlO6RRAvkYix/l2yJzMxf4PDiapJw0m67HVJgDAE8+2Z4o2WLe1CKT2Mt4d9JwEUcQQeeA9Znpsv
dMJzo/y88FHAvtpuL2sdZiRkmO4xMX+LMTVScSYSp2ajKiJTbsmMJv0Dmz/6uhKHAOtb+W6qUzMV
dE/8IdQ7VTnhmxJ4eltxhDRk1LRpNTGbtTjcjExk6ryz8ejBSaXw82a8aCyBXytzzzO8I+wYyeZk
IHytJYTENYG05Srm4OtJlrNwe9ODN538iUSgOBekynIbaDIJALXftIBSgeo7lmzyGm+Ng6o1jAdb
XPl26oqyeN0iXa1+Nl7yZSjEKeyG77QHN9JaekekQ6yj9dhKjl2/8+L3P+ixEGaa6Bjs5vvCR8aW
s0vPNKO0/7qZhOe8Q3uPKphg4EooX0Ni1fKNKOfne/7bw0yUFxrYYlwmrDev5uOhWmgR9ZZIBZiQ
00sql33hm4+PsLR+pa5IoS77vEEpVQV5wkMBbmRbL3y6YIFYsZ1hf2aaWWIu9/Wmnd3oVgGhaYHP
Rvs0esuFy7MhuMoSsHWVpsZa8P4fkuRGhZFBmP2llnuQRoWnEhWSYej4PsKlFplQlxdCosCQCmIU
wPGs7ooqmt42ugqkOdGLxxALk71bqzd/u17WxYZcQat+ONhVKJd61/JkXRU7G6qRLgnqQS25WoT7
+TcauCFrFsMJ36q8VN3DbVLTZLGRwznZHSDYJGhvnfqNjSRqajn8+LQXTDhXsOUYUBiXTSmiefow
SMBtxQ8m9e79LUyV2TZSiTwYCkLPWf9ZQKBhBYvmZdTWKyax/P26lChgq7exn+tUjH9A5SEBjvfp
RZnADvEnRF0EMZDTmnqjYUapt7bZbW/KqlFxgnUJBbx4foD+nd6hfJk6a8gizwt4JckWZLE3RpWB
94RfXlnsFFQTnw64hzrwiFhIb9/XkNQ2v8dttSMroLtm/qxZN8ekl7XlVXFdydkzzQIO/0QAAshH
Hl77Qbed0mPvh8qdYcmd169LngvscznLm1M47J9Ynn2p3Jnqlubl+rSXyebJilKkUKjdDTJrYOl6
Ph9N6ccllmKNDrgEkYdZTQQKO2XVBjCOkdraThHPm0pf4C/N3alm95c7YZbMZWhOm09hSL9gv/vP
+ZHitX9aKmsMXJyqG7W+sFazOt6JL+G6HFWCP/IShadRKmtd/kohYfgqdtKiPAyP+EcMogQ0LdYJ
okWTqZarepgb3OpDXZAT3jqaLOdoMQuieFsNdJLBJXzDhDfl0V0QaOAIkGG5bbEsIatG1duzi478
eJEQGuS5vAiuBuUNVjP9R97GR2QhC+TU+Uuc67pnXoGKZaDT6UoMJloE6Rtza1BE3PU0MnQCVyFO
BD+JCiV6/4iveVSBU1MZab7YbFv8cRrtmTU8IDSdA3GeoNDlK1RGjqy5nVYuYJ7rTrfegjiSiESi
feJWGkif1CC2qWX7tYd5UoYXSKhNA2RqSSgYAqTfKNJvWtg3bU5gD5+UDzVY+BNULqsw1Tk8cR1X
kHzH6k79nzA2in2OwhbEopRSBleULhHp0Hr2nf0ha0whrkDABVh3hOEPp9y+dDXysok3UW51zihp
anEIRZIsMtsh7UH/iKVzjDH1MBttuaZew4PshLZvgKupnmu0NMU8qyvjQCNvPiVPQ38zFfVUUN/c
1s8iSjsH3TSnbVIl5szJ+Aak7j1e6QmHRSjR0HAVfXfshFRCKScVvBMjuSOihlwVU5O+TZFH334G
QBrh7YRg4I92WxSidxfTDsOptJhSLmqfELA5N/s1FPf/7gruv7ssrX+YhysUSMOuK9WCWWa4Avc8
8oXPp1djHbLo3fSd6drln/pQJbY4yPnUglhXNEPdOdTkEX+bvVkcAm5410plNxxkXOjFRU0b9Rv7
VoDwNZsbwwA3mOzin0Y3DLsodlEqbo0t7iNpXj7Stvn+fPwi8FTFV+Gy56oj1WGqMS9rhgW53166
8ek9i6nmDG6/s/fiGp+Bie3LtHBYibO76a9y8MVlo6mIIVCx4nzFoCH1zmQ+JLOwYunLamHkL2Fg
s3Sxt3jReF/W+WDJYIClzBv93qYSZeqeXWRUg6h8B/CSjrMIGoDq6XjCqM4p+5x3P789SEFkJx5z
vFt8Qj6pt9iuxqLvPhaiQ61Iiqffz9d+C8Sx10PPOWHvjLScq9YnH3H0rMcZd6DRcJeCPF6/N9ZM
BK5VV5/NBi7xunuy7OIz2d9CjlT783RqS5LGqzdneweNZA6HdaqPALE8bdJ1m4uBQ43OhADRmllq
Xx6VG2v7RK7pP00MO+i7m88V6oTBuTfEc0lrsPYCvZhGTLOU4xJnONVyVDdKhR3oRiJsBbdAShvq
KYHWH8dMnqI/GUCjw7TqSrBJ/9+ZVOx9wPdhBRXomX9tNo0xa9JNckaLXAWK+ocJI2bylLcGgyJy
+GvOScGLRbCsuq+Mga3Lvw+oH8uH9G4aY1oeottbnPqY9jOr0jxcXSn3WNySfHKtIB+LiDXf++gw
9DaNLy+c1Nh22ZnFeG9Sjs7aTnqZToTi2aKFubUPUVly/DGjoDgx5jCoV9gWpYWyg829pABfqUFY
F9MNIqFJFxru5vzbIIsC7ubn4u7rzWR4OSg3gt7r8L7c1wxaYzC3may+/slti8G4/+iOtt3Y2oIb
5HS9GsazpzDyUcQrMznkuZsczS/axuhcLARC6jc2GKEJBMmBVrI/bKFNXkHunY/lYZmWkvYroObA
y9pg5RdhXoXCsFxHmcWK4Feek7zHabSwgD/p2u9S+qpPWUXvwk1m4V096oYgSfp8kUINo0sTiE89
G1XSI5ChvNIXmhSusQBYEwQjglnoIQBP3IhxU+D8yZoao4nff5R3IUUo4Ro2SIRe5WkphW2uy1e6
XxZMsJaD8E+5+NOwGm0fhTExlLTNy1BYaVfiB9+XdnL/cgaerfGKmwr2UbJwYH0/evsCV+H7Z1AN
7mUdnZv4cf8phEIe0uUsOzMe2/qNBkjmemH0mSWWdu2woq6cm1V5wgJQd3Vws07Yl3n7F2LyOYvn
fHvJWdfKE+x78EhqZJCDIU6xXwsGSbMXJuYU8wAm5b/MqAp+2J5eWmTmB/33xmim6t+JVvLAhJcZ
cF5lQNCEug3+j6vvEbpCVhJSvmblmazUF+VCo8odYmILupGwdJmRZXoMEC0yec9lTM95MHbFqD1L
9mpSFxC8ZI+aJ5mDaj63Ljg/7Sq3bZ7zrAyQyHKgGfFKfsJjjrn5CsThJoBSaVR+UHpGfUIRiMoE
A9zL6PXEOUXY6/WY6EFzGTAqk8pUju98AWlRO2p3Edy5wswQjZI5zhReY8yyS0reo/SF8TIdqL6V
SOCSJeft7Iqrk2ZraaMbfFB2v2SGpQAlnGcLwnPCHywNqsBMKRrYkg0m7aa/bwq2TNo59WoHHf9Q
lLWuMOTEF3IO7LNvsjZqjx8YKsuGK+M5eRVwz1hvv80lxDD33PC9BNFweLMQ+0SjD4ItfZwIpkHC
xRRNK6DvegSeidJN2TtE0brZgbfJk5KUxF0oP5d4i+zlHtuzbUrIn+w+3xLF6qA9E5TBrvgdd1Zk
4wE6zF0zyWkCq0bYKU5QcKGtYnPe4KYnFVpb3OJ2yVrupcY+DoeDeUv3Oh/EWPUw0pzC4E++swhd
OIY/2s9gLSpp7nJ9wto6u7L4dbRT5m27jaT6doACICzwIZ/we1MqWynqJy9RLF7QxbOQ9SGyHN/f
4IUsPdFAcbygfPI1n7B7HHBb1ODhLQjsiEueZNqDmZmf4x3n27BAOrl46SMtlVXAEzrv2fb3+/nJ
HbDQVbxKGwBwz1xHO/waTSdpQewo32tpno8TmvlQx0JlrCu4hdSoPNm9hedA9vUCr1kK8Tlu/gNh
T+zRFVN26wX3RmVFX8ZcxRtJZzxMYiI+qH3pd9ROaW07bG7rw2vWMVDB2ZhSml6j7uPyZWMVDt/G
WyYbb8Vm6UGHHrWHgi2KhGP3u1qCbLfYXPEJeRLMQqg0fpA5zYEN8p6Gg1yG8ajF45oXU99Lf7Ep
AhRyrCM37NjbVx7BSytFRynqwh5bbjz2q1noSG/2n1HVcPJUweoGK+esnL+ECHgR/SGpIXVTyvyZ
eZD/QyT9kzmttHhDqjvt8srkKhxcylJjgWSHZE92TJW6ip2vtXfB5CuW+hEQvCNID6fbNKDr42qt
br0kGtmRFwV7iiRzvBfcT9WToa4Wuh+mO0RMIsEEt6vhFOz2QzyQ99nNKET1i6IIgJiiS3/qGUtC
BbDINEpk/1LzYap0cqvrbaj4JN8reKS7/pFioKs7DAV2ecbacZnpzq/Lxgz0Zq8gQae9L2wNtzNO
UJImdzyIc+K/mU42BJArBlaw11xzFDwY3RiQlhtDX7Upr6nbfiVnl6LFRbz+tUe4spq8YuyLNY0U
LjjVX4ydGUJRi061XDF+83V5SFumdbXzbBFcU7jme1LL9kB4iiKyFNnyYDMvTlfTY4tsEquIYxF0
CHDP+Ty6HpUfI1GyCa61ZDYSLQ5jDx5zxvnZn8DvjeLvzOV+7AV3IGSBi1TKxVPz7YCNkWX/BqPT
T3nEqDtAXQDG/WZ1HHLmbjXAhYjpa37spI92SLqfNBGFLa9JmojnW5iPp8/f/i9506OGSbkcgtjl
owznFkrsxxKTQasZdN4o7sxeZTFncbheObZT2LUQ7gpKAct2JgiH8eMOhMONeArJ8LSmorVPDiqW
srWq3SHzOkXlLrNypCrDA+uzH4JhoW8jLngAjELQfDOdQ1RMTccrVGupPpWp5T+BuXvcaX3LzGdb
dyQQGWO1ftQkhDOeoXUWloz9MZIx4SqSfqxj8030p4+SOf6MVrgtJc573UpMslr5cq3r4XkW0EVl
vYXkf+hAJXJtjaH61CH9jWy67oejJ/NT4Bz+Zo5PUsbFR8hd45es8bIvijQONj26BCuvDk2otUBb
iy4YZ1/ybUuJ+DbVXWZvjkbAPnHlODpu5UWZDD67p2xNnN6PCf7Qj0kS4IkVf44cWVpzRRT9E2PZ
7ZJfV0l9zUy/Ad2O6bGYw/JP2JwdFcYrS5TUdTvxL8GlC+2r8aSYBO17OXpEmlii7Nyg07XcfdZr
ZTxSFmbY+Fwz/jTdiUCRoslXSmQACP/wnxZqut3Jj5UpvzPAnqyXABT93lyOhumaulzD9X4DAmsF
ki/7LzYHapvzNDjHeD6hhX2GxNq6TSIPezfFuq4t8gBJEVVq7pisFzCuhWgD/KXK/krqWLGIt1z9
CwzpgwQIaCjudBqWXOyk/qzUcfdnhj9bgzsI4Fw+NIR06Zc6SkqTImCDtql0IS8lQFFSaGeflL5Y
qUPHiM3iHS4NPLxEYWWuIucNXlnv9d1gsYIBHLjmRyx6w1WD6DwQGq7RqnbvO50Yo7EIciXwMvBI
8xTNbNyRrTiwzrM7xrGXv72VSAifbyjF06JcBaeZy9V5y4c79y6Pi5oVDmB4RrSotMAsM3EPMCW2
clr/BoGhYwlaZf5W/v1w8L4sX2F4u18WjOcExSsHi/m6TMTavIQnRGIFqYB6sG/EvPz8tqgypAOJ
C8jGayfNiPyBHF1caqT+eip2zudnzChzdkheATVLq0bHBzcclMCmq7Mry5lwESRY/XEunTo8FC7A
/w5K5PUiavNnYkc4Z98cO6Ye6QBfudLS35Jdg/VHnRfzUVAJ1pmSc7gHV2N885ctS0Sme/IlFBID
8RWF69YqDXM3QzbuU5K/56FybpbZqdqW40lIqAqz9vVGZta4Q5TFGbW/ESWmEzgSoOH2ptsZtOEv
GUr4DvvFEyPYBZzOUwL6vCIG/lgjmm8JfLGe2K0uDdjRQGay4OehZ/bqfL7oW1s0ilOjPFA2m4SK
cK9ubb9dkziRF3YDq79jM4fnY/NQ2FGXcRmCPmeQtcwQoTxiyXKMy9crvfc0qD7DZp7OKCzLsmbl
l6zF/QNIXKZ+qh8TgiVSbosjL83AqWRuzbYj+Y6Vy8pS8YojlejeQkidIJ/O8sh/rU3hEHogFyAS
i9HGHL+XOqO1WfUFSmnxQVd21UvaoayZqkq0jqHXafpw5QQCx5nd2N1hbJUoKpKCbAk8BIO5HZnF
AVp2yzb0qHe/FgOShip5xr16YaZfrN+QwrGcsJrYp36cTGWAwmD4/3UldNmfip4p1RZJ8Tp0079H
eWQ1tIrY7oRbhbYhjGHOZZZSzOToQZF8LLTA95Q7mb4yoQhlUYME+EWFVgiQUK1gUFyBRHHQSGBY
kBICDZPM/IH4ZJJz7OfllCWWmNxr6abh4oKarYCWHbm8dGcduiyC+R6lSw9xcAnu0CedPB5ZxeTh
FvJfms1lzSzIDjecEMMaLjnzBsfFsyJlBDBYD4k0MS9C4aN0OSv8Tkvf0PFuH8TjLM1aZK0yZDK5
y6Z2SOJsVGGqCX04nEXUSy+VgimPRuJOcYUj8+PdOZMCfUTmlO7hkHla6iX5Pc7va1d95laCeJlm
T/fhn4wZwNQc2EOXP37md5zHUPqvXnf/KOgKmr5G1boMCmvKhZ0TilqGhyDAHo5CMPmtwk3O500D
BVm06HBZDVY3uG7nDWm2g8BG7DFlgyfJllruZPg5S0fLbyFR4zecyQIoFwBy1ZZWtXqPeZ7owbsb
DFgikubrZbSBrekpUHN63dql30s/lEISaLWcZ9TuVNKkm9fOo0ntfyBw60ttQfAGOcgtbVStNLt+
CdZOGgUrSwI0vlVH2iKJXyVf9gOBvRJSUdNb+Gnjdo4J8HYvqErL2BCO1773wJ1LDHWoV6/G8oXU
WS7xyonD2mT/kTTdICjEKY14SEbRoPeyR6UymusyI99Sg6vgC8UuUf3jjrLJYOWLcxaEIcp0qG9U
2+Pgh0HJR2a7pSTwZ9xtKq6A3P3TX0TVO2ZFUlxir6Nw69nuITJ+HraGHeZ8Lrb+pio5ayubArWu
+DQ3X/qxcgKYBup19rP+H9zmdpet1/CO0TsCgEBwcpkygJIauMDGfwDZYT9vbf/BjC2knm+lMcj0
1m1xPkUDLt4+Yf4BhS0vaZLFmhymzOFSkgmY5SwXSxAv4phVFNZ5AOUzqEVlfirroNCJi1gVpQ0h
RXhPBtNjk2YeeUk7tdWKgwOtv7QTuxpncp+xd4V55Hwukhv0zjf9c6hSNbo7CAxCyCYGFQK9WOf/
vZpIeFddMIH4I9vbK/auy790E4NbZ9ps7M+DHYfJiWzcGj+cY66NIABh5Orh5pyJKSQIZAetmp2P
wXqeSJhGdbPfMuRlyPwfjn7RKRp8RVdjHjQR/JBk1hLqnt9ETj6GvJe4TiiGWNKK8+4Hgwjxp86f
ZQlN3/RYwLTLjNUbPOMD7Oaz0x9F4NrN8GyvQLwsNZESv2DGOajpB1iup9Pcv4aKqGSZkRp/ruBd
DUjQ1+Jm0hQ91fGeOHK1xcYMJowynb9CKcvVObBoxMJrfliyumnlJsU5K7cTLGAjd49GpoQuiPNt
apE5n594FSfPiUonbK2HNiAIJwxEwze/oekhUG+ebwe+jN3UIHbJMg4cg+wMKYspqpXsuJoV0XIl
IqMdzj6pifE7UKhipAneoEO/iV+RlbjoJKXGUTCzMt/Y6/ZCOdX79EaVLqGLubeF28WQFxb19yZM
eT5S5fWnnRthE8xovh6UPXuNOR8/MiHKFxds1xmh+Wejnmw5sjAH5VtMSPweUjcZ33mVizvt/XSi
uXul8CG6bYr+sDObFCa2FAKWUMlP9ylQLkNsUZsVUaLM3GQIUOT/vt1E8t9K4k1g2MvL9v85wDsb
xVlhaXxxC8bjNRC2iMOVl8W7eaW6VEYLGAHJ/S5tT2LMN31mnoqhYSHTbYN2ycagRajs0lDa+Jfx
O8ErW0fv4956jYVB2XTgFDRxb2O3GfnhYy9PCIP8eu99/gRwa5zTEkvwLc7N62YoGA+LWcTcX7Oz
p/Ullmakk0FumrKFlOt7EV3agUq5Niy3aftEv5Wg83Wz9jskmFGZoJfmnTrBa4kd3oZC7J3aqJw5
tnuGGKTHqWINfH5av6n+MhC+Znw8B4wBpOJkaZKNu4CFj09KWZAhOmuez8Vwmf/h4v66Tj4oFOof
nGHzm8AylPWf4MsmfSbcnZ76P/+xdKvA4EdCc5oL+a8iIMS0mz0ybws/1hu+xl9N6EWMW1sPM9ot
CHViWnbCBM2b/BoAPAq70pEwdcwLiDPKshI5dkjHpiLUGnO+PYGO2m2TOAFhkAmunC4f4rbupgG6
oPEAo7i/NZOBMTsCyXYa+X+ULSlYS30yR8iQgBlaG5EVwL9KjtrViTFfla8VGUrUdklI413FCuAa
wEuvlaiwN2yHK5k3cHWEgw1W7iDbksugOmWV+wNc78N4NEzaVPbxlHAX31ybURNYIIi6yKNSyBBf
Be1q3B2RvJZTIINGml0wj8mqe+tOQOM9iUE1TXmQCzJBn4v0K/k1kzJHQ+Lngfrr5Kggc94U1Gh6
/xL9ZpVJ+X+iewlpxYEQCjt7KBa+dhxaVMlC+G64eghwFFX/DJiLJDLGavncJxWHG6F4Wy3nopSU
pGYI4eRF+brWBU1LvJljp/mQzam3ctq/P4d2xtQzpH6NTK54WbpvJ0r9+/ts+tf/afMzExFkBPoa
ygd/Pg1JB7kNGKRlcOuR08OAP7+pA57EKZc2WnyEIss488tKLmyC28yO66Q3u9SY/W3iCEC6c7xN
hde26BqPp4VctZB22Z2XZpTPJ/WCMHk5ogtGZJRqRgkQ4hUOuaWYt2EabFcHJ3nrq+B9jj31tUC3
BtZT8oX6q+alTVKH9EKbK6+clE7ocOF/wye4ZRCSyVkr2PUkiHZoiPX2HWOs/Kc8ZErwqKYSi+De
qX2ZS5W55UStPlXV+cENU5DTjlBF8/kbv25kqyuy6vx/jiE5V86VFApYqtugfBQMzPqmsdFan0LT
Op0NIWdMHsqZqP6X8+g7Se+jarb3n4rUCAjwJmCOUdXj1aC8TAPLmRAFxUwzoVOSxWV1kSlfbPv/
UwZGDi6F0nPzD9wTwGq8+acnzGKDZzRfn1Id2G54iFcyZuT2MAPoYKH2C+U3gPyWzNf6FlBmBTnc
CmVZcs2J8jJnIh51UN+oQ0+SYVKnUvnj9Julr/xa9EE7/J06RRa9CqRSaoiMqjOD5u0qS9V0Ry+d
oeyM2RYlgoKY6cRsCMMkCPE9rniZAJNNfhN58swD0sl2Vb1LPBqbZeJXYe88m+6Zl9AUXCYNElZy
n11En1EgcWkckMOoMsJynxCpgcSVG7dcDx+ZqfsEC6fQcIB52K4TCn0oFzO8ofPQxET1hSlFVqvl
YZ6caNyLlEi/sIR00GlzAvF7xPKkKPl5SjDIKtITuZf8PGZZ/YpGOE4SVHcYBauJ2sIUY9+nGcgb
UmkFtqq5w29xnOLA6uYVMS8sJ2PJMbtb3gzrmGDRzDzG35aS7dI++pevviVnNDvEk3AnJVHo/JWj
6HZTd/ezsxaBWkmHNddnZ9yIp3Oj49G37oHLarQdkII9SZrLdROnTybqWCjjewLE12XFrMvY/kb/
1q7dNp5w36w9bUnaGJXEthz4hdNspDPk+QyrnaP+bT+mOaR/l64wmemXqcYjbQQM+G9PaTzxJFgE
oNPw2EvCRcHh9cqN78PbanVTqFFDQ+vQxJYyRgCaVlvd/ZGyvQLijx9h6duTJH/XRi2Ou1y0mzXw
Lq2O7EJ5oRXf52twagoyjRiDA9N7shmQ59XBudU+hYVUZySuVydP1LmD1HrJWZmZqFGR/QBADUSG
X0wSCMEbgJm90xpSTdMuUMyRC1HbgKSnlOYKTnKxkqwpzAbMOsz9yVJbOs99dRfioOe7ApH8SB4D
R/F402N5aeMPBOuLX0AfXgyR+Y0iV91E6L8jKsSU++QDSlns8rW9ip+GV+Dxx72M+ybhjrNnOsXk
QjRn8M67eSemPbS7DpNCf5zrrOA/xosjl4/gGs5Jd6WF5q0vko6Be7GCWvq/oIdxGkJtrA+RZXnE
/SQOfmD1E3HNsvJJbllaKwOnMSmNSakvZWG4BEc5it4GiKJmPc/2mf5wM1ET/zFPjAVM+Zn8OsR+
7djlK21L9x9w+AOwpaLp3W8B74+rpy/645nt3wttZ00b3B0N2mYvF3pgHjAAjYw7PGjDne5OWEJn
kBS1TpAf7w1tTnZIsidx8Bja6ZfdkG6bky65hJJsSy1rFPtOq6uti/xioPpUmiLubhNw849MxK32
PJWdecqsLwTSvbsx5MpcCPEzIJ50/ySYkYDrQKj/lepMMi6JYjn6qcayJqIWSX2ycMDHykwpgetJ
fWdlXFmiB0XWulGtHETBhLCLuRuz2JwyZtKiASGDE3GrF3O7Ai+nZJL6Wdfm2VGCueM0vFIcPQP6
Ai6QbX9e4F3rgl1YvQOFTLtM2HPDTN5U5GBu1lRm/D76SkTm9q7AcbesF4a2DPcB8NLkaoYzPmJu
meuUrh0cmCwEyLTF6iCFhXO96+B6luDHlrcghcs9QUGFhoQorpjda+tjqQweAafmj/t5ay1Nw5Np
VwQa6PaTTsjZLGI44QPzpP493/HI7i8QCLOfK/wXUN9fWuXrwi4VrnEyqLwN5b/9S2O2D3Xm+54x
5Yq/d1xUBq3sczJAhpG6WGkVK5fNTJRDWhyIx0Q77T6c+DZEz3F8GDA10IsOJ+vby79d03aUGg0N
4xApCtzug3SHSSDjgAk7A8pZpH60gLJi2qdsYq8WcGlilCplP6bwSLRxlM+zGFfuLr1/frduZMZ9
kxerxfiiT6xTKBxm65mSedxIRbN51S2mkHWJhZTkhNKktc7S6A1DZ8kNdm+/FRB7m7w1fIGHWJSl
hI4tdV9LJj2nEoXBakAGwXQ0dOu59+5D43Xb/27Iy2Fgslir0Dhvw9Pt4MINo7jz2IDmq7wFivC6
piQ7id4oYKVLOqpHxIZSIlb+EEVtfJTsjkxebvpIDB9PId85GGSreylx1ytbETKhByosJ1y5Qesy
R1V1eFkUCpN7SznjK4GmYj+7379ecEg8uYoHuWiQnunKsb7DPIi99C2SQ027fIJkgaq4f3uOdVKX
/HVEWmVQJeortjzhvuEnut3x8zVJuTcQrcpW/FR8Ctq4t+QO9Fo/Ff6NPXfiFruC2uAzu7zgONk2
qSPVFn0U01VQkRzaACJDGfu3Q3Nss9+c5KSiQPom783+zgnAsnpwFa4WDfl8K4oipFRhnPVpuXYn
82U+phE+1vS2dz86PpumGMZVxqEdOaQqDDKrj/QPPTuMCcHqdvvqQ7i3TOUO0oGnF1xgpqd21j1B
2ILSNZqFQMIsq9j3q3ZvwwPsw4J0P2bJ+LjPDM6QGY7hzIx+3xVzTEh6ks2nqGJkQIUTAe4wuBFw
beSo+YaQNWDL7hte74IePu+A59eFjz0pow824nCy65wJP7WLdnvqhMgQn7H6vDqWg92Ar+duiFaf
Fmrc71mxSVJbKBVqz4UIXV8RC9amR338JLG7TS/aC3O5zuZD6z7Umn7YuJMuA7Em102bVjIC/97x
yrRO10iMzeoL1Pr2wAPusBo1TRT0mtdfe/LA7y8PrqRU7nsChI+YCWhUqmq3rVKHANsnfxn7o1os
4gOhafR8kHqZVXz0qQOyzrCv2kaH6+5uw8qH0elqyEFymMVL/pdkbvOP/EqP23gB8lzgEIxtqAbd
7RlEzGit5AkhSlOAMBylV7Oyzw0R7qAPTXbhu/0BZRGRfu0LkEL+1IAVjTZjul7dkMKwKB8W4yIo
u9To7FS8a9W+p7gEGgO1DZ2z0yW3c2YUbYZzFQ79VgLMH0B6d/jWt45Wr4k1bf+nw1ZjsfN7WRoi
mJ1XY9WD4ROmEau2Hvt4wbszQ8Df0HOFnEbYBw9QzQP1Aio2OfV3IjPNy2W/zuKQj6GtI17IE8P/
1dT4BPQ5cOkN+/xyHPYJ1vT4ldTXWwreW/+ceKn7WpC267u6misGtp4N6IuUfRdCdsE/apeoP+cd
Q76roOw9GGdJsNk4J/I6/WQEYt/9fZv0UO/IRMTdRY3yReayF/qviDL15+tZpYpA0EMI64W5SRes
3okPDJbvlp1l3flCGcd7J9awrai1Q7OGlKPstNo0FdBWx9MZPqLPvr5iniM3sPk7KvVAj59Po8+Z
Qlt49LjgEvIABGppnTBnSr+Pbhl8vh4U44yZePl6A6UD4X6WIkEfAt4TfGKcgVFVs0MZthk9sKzO
P+NrMbS/ojiRaKnqyr5fYyksw2aT+fBE+IZ9TIc28pIH8ZIR+BVD0/mTmKMXD59Dgt8ru4ueKmtL
8OhC+l/QwQicWu0oi/zQ7Dr7P2IzCIIXC6ZloPUw5zpzuVPDZYGvQjQcrnZsTY0u1P1NRGlbrwj4
7Sa+v02PAaQ0NAw+q5tCiVSmTe63/oyhACErK0ehw2pbCK6QMwiyzqYud0k2xW7IrVgNHDGmRKQX
irccYEWy+GNUrmQPvPI6wnSPPD8RkC3E9pugeBuFUeV5KE+K5ofoDfXwwtrkXH/0+Nf+0A6V7xLa
1bz9S4ELHav53q3CT2C12BRu+KRwRSkrPvSCDYTvNKsYug0DCnHdcebiez0mR26Pp857nkZd2A11
wfaEli0Un9L1c0g81vqTaYQ32xwBAY0bYwY2M1NuELqkECVFXr+rC1LhOWpH4ofEipzFENZ2OOLr
OTAcDE4VmLUdS5eO0Jjkf1yQDTlVBQ02h64bhgjgs2GM70ygD37FPgn6N/v0fGH1zsWUGp1BBvhW
RBo/G6eRYfjLIMR5L1D9h48vGcImb+4hrbXPvuTeYNgcmT4hkBXeyDJLMNtv/Vr+Z3iDJ0ofcSul
6bKULj1TBlQn4h7x0KhkN53H5pqOMacgg7uAHRP4RWQjadA+nFH75/oWUWe1/ElBHO1BPTaOS7Em
prKHz9PIaqO2vhM1rVQC36Q//UPVr1C/GfytNBsKsneicLVPWX2bGHYIYX59zxX2i2Ee1rMi6qc+
Sew3Gc0FLynf4ckOozC76ue4aIH9KL6CO7DCpnPxVJc/vQXNuEBK2kTgTuCEB8zYabbBpuYCE3QR
lqBL6EQj5P+s9eNLu6kI61v5uXLdyrERCUZMcMHxJL78yo6xNi5Ocg5ikLGLNrsqgs4EG+EciY/g
qbpeFKWhQ60YR//eXw0rXQxzZ++YM4BOcHIIavqQh/7fszIgAFkeGPasnwQIRAqKWV0LgFitQFqL
TNxsUsyUeG+mglfb/uIe8Jr5TDSw1se+noXkXXdN5F6h9NIjiWTpuPxnXDBpuG6LWP1D1qUVI0Ym
waekg/o1zgBrOdaed3sFNMpg6Y9EEX8LV+SL2gFT1afkfwc6h9WYijeLZNhtm23dGmqQzBzvG3YE
npburnzpGqJx2ayz24R1645kXh0eskhinHgxfpM5yM0JNUCDtWFtGVjJfcfEneW7aquzKiLQLvkI
AnieDzD1JByYqlLGWjkk84IPi20thwT03CZh4Zp7Ft5mxOVzmg1967nx1Wy2CGJ/0ThDdpGFDltV
OEZavmOKdPOrYkfbf685adgO3M8W3YXJXjyvIkDp/umNsno56r8KJln8JJTZKAwfR8gzEqxl/R7g
+2hOSS4DXPjPNuAAuIYHosPIdvfiiGkuGf9HEz9/rNE/II1qf4lFFeaHWbixYPaD6vu14RJhxNGo
aZ3O6yxE/tT49IQ2ZOVbNbMqx5O0u4j9dhK1g2Qa3gWZ7p6SbKHE6o4qtTOzTfEBF5i8ptasolFb
lzdRlicjcVVmHzmtOMCBLIUCPoQ9PPWTWKxOxoLcJY2Vm8qkH8rss5DlMYlo9LXbhs4XK6e81xTI
rAo2UjUEspkxoBHJRHt68p08r+oOK3NnxiurHJSb/j5xDqDU8pCGtamzHw+C99ViQ0UtmZNrRyIm
YbhK43lWDlznNf/O1ahRdTf5b+8b8ScKaY/lEiw1T9r20kI+8DfBxw+1WCYYpI0pGIo+MCOBWaPo
lIyG4vHUUm6RmEJc0iPekYiFdPe2gEzm+ImXomsXT49uHomtTl8hB8PwBmfuuzcAtGZIwJATIq6/
iU9WxCIn+F+hOtoPMuga4TXKu+V0S1HwYTg4Guhnd2+qTBOPXCy3SNXckETpoiAg/iBF4KOFE2nP
ZTT/Ok5zuOKPv7sB5FUoIK5A3HXKj7r0Ves4kfcakLdRTbwhU4QD7jzzYJOT2bsxykoXxSQbyjCj
zMNUmgWIaxCvb72eAyjJ5kHMIeM3gMRNv9Oy4xd5e0s9Ra+cFNpF04xXQ7AnyudAxhzQK8an1BDH
3kLJCMATPBukxrsUoQPhCDz7lnCD2yIdcwxK2jkg7wgKM6mpEhvlSJbUFe8ETs4NWslYWFwunbBR
wodU5z03SsjYOat4nrOZOJvgSeb+0D0/r7WUNFyJ1iN4hGjAW8xgnm6FNXsGXOx6zjpFjztz3CwJ
B+jFCvYri2B2K5e69oqnFBR6MjzukcBTcVXYAP6tLRO/dgO1dbSAoLl8VLE+YbYX4feKvgQHAWy4
4cNVGLjVUOcrn8HT2XEF2BeMjwJgaxqBX4do3X9OA0+DWE72hufvZv2rwv7IodH40ebKgMZ7n8Ot
/5pLaryJg8NS7Zrp1P/MskiiZjODAhQtWkpEmSAPcqnz5tO/dgIrT+FuUL4Xlvjj9UuS0tJ/YbCi
xt8wWdxuRqSoG/iTebfBLvnFbu5pOFB9Hl+ESi3A601akAkqgmdzfK4hnpboRl65C/Omlv8RE1of
KXLoGdcwIfV0e/UJyYmz0MoptuwBdal+ofBwKWlAyRFAnLvS7PP6AL8WKPlFWeE1P/OhdXxl0pRX
S1ujWyBtHflJpJSkGFeasZUkuBSjf5wVNyRSJEn7bIjHCdqJsOla5QD60cU6PrQcim53HqNpfRCN
oidusuBNynFa6EFvIh6d/vzkcyh3nqifGySzdXFOyQWjk4VKh/GSkEdQfPr20j5ydTgREd5XCPA+
dHMqz1mNNgYoYmcpj3n3/PjJixEqyzjyRUegvBT0NGxPhb27WzBIomAveG950yuiahtMw3ROiAoD
s5LiBpkXG3MPg6LDT7NHNkP5WTqylat4FwLJxZqPG+E3vwFXf+teK1fh+DV3t9U2HKh8KVE/GyH+
hKpfncZWwKlIWWzeiBgl9kTsPNBLh5H4B/hIrnvl1XPvr8aZjddPe+HF27W/YO8j9y485B9Jnqcd
SjGTGW5/lBKocV03wN2WXtECJu8B2Lm9mT0dR9KL+slM8JgX5nKZ4tlFbXzBiC+Y9H0ktEw811Qr
1dyejH4rLyLTuBopc/mcLjWeXNop7IEvy43rgqw7XPIM4EC3KKfqILoB2leaym9AY/QAwEI/2NDX
Yu132qi7UWqoM4O0BdTROm/lqd6Makhiyi7WFKSbtjUa/O1n7dFBCJrQE4hjPA1yilLlgqBI4ffr
a2m1SQuGKJ4OQxIrJaXEts530HJqCjgMwxLx3dO0TAO+6+rnP4Ldo4cWcov6YyobZbhjiyRrdlcz
IuzUqf0spoXN92d9CGt0xPS2FK/k49WtCi2z4VfUc7KYp6T/9+4cPC8rBt3E9N9/uwGfK4I+XuZN
ffFDKhOLOeI0k4ANitzH5WDbdXUq1a5vYFmeMVj1Hd+CtPnqv0cJCCtjjaoLysAijB98N7ECiMRG
NnuyvBOeM3S4mFLdg6DJreiaTXFx/xA7keW+Bvaa5v84U/oaefHOUxxrF3IL1Kn5wHcHocPQFQWA
KM/4EJlQbIrqNX+yUxnhTP2a3CAqZPL0nFDsSjRaozHz+1UZGUU3sIw6LwN2whd1mYkhfChfZdah
f1pt423B7PrBAnEtgnqQF1YCGemaebLXDlxMRkFVMe8G91IlQBoorXoZthQ18x/g5jjSBS7nSJKe
c0PJz6d0ilIB+Ae+7azwHuFgLWRbdpJw/M/GdzIj9Kq311Exh+uB0nAADjNRLSLakJdsx49PqMTd
dbAPBLPYsFdwg/Dg3EnzBm0AorOkj4koelQLc3ERR8WXBbIUkRlPsNwZUDQP5wLVB7oEzxHzKcbu
iLKYMIMFo8xj92BFZ/4J5Yx3paqcmf6IIbJOIdTIartPoBb8DuX3EUR12XDXoco1qNoqXZE0vnGD
5yZZqGeU3Acl24L41m0g+gGoWeSJ3DwXWaTzRpaslQ7oQrK2czxzMGzOlcbRCDlTf9c0JZJIUFfy
Qzsja3QA9kkBF6FCfoNgOxv0uW2PzKvcdY15JovyBdGlrry8NqW58ljad7RH4rs9FLqliuE/TQv6
iSzrSLjb8PqyHnfVdFx4NvRBUhZQ7NNxGcHzxPpKrZFpd9Up6yQHbWCvVeSHWsPJrEjQlAO26Ckt
xGosVyfJh2dOK+b0VwmBknQLrRzuEO2Swsz1rX05x22g/RLgogYc5N8aO+S+jzDIQn4PDDs3osMf
UjETa7+QZj18y4Il/EzOrs6ySpdaAZuXJ+Z0joQxszC4USl3XVIXM4WQcPNydIUb8oeQoNO/i3Ri
7ubDKAlr/wD5236FpxnZINv6J05xR9lF1kDy/gpALn1IlVtE+gUpS+VVXnyZMG7xbGOCz1kmpZIp
66ixMrrmF8n9XG6GHv4MVMx2rRR7ufLmLryfTBCW9XPrpN6n+typl32brsk9RnPHbLcdZAfxDfN8
guykX5IHldsJqISjmT74ymBx8dX9tV0g4jGUlH0DbRm7NpBXA9bOQcrqd6b0fRz2JkJF9g65Tio8
pti9AX0bt8wRFOWv38HeON85Jfrw36kPwByWth6o7n20jD3vrEsoLNSmYdZ+JB5AW+YQXkuXkOgK
4k1zdX0x/9CtbuE/l/W2v+EHESfFQ/+4KnisbU64VkNZwvsyh/3N8hnvCQlxoYMBTyLMV8DXCugp
l27ewS4EvmzWZjnZWwtln8hGrGhOhm3UurTVyoiOcGuu6UAEsTtIqiGoCEVexjcG8v3l09eySR9p
mlZjf2//PaeWC0sljyXzBaN16hQAx958ylC7F2ZbG1kwmrGX29jMjQ46j7M9AT3fDOx2h6XghIlg
cYTF2SKGTmh8+Q4kmPX4KKqxN4aoW1T48mcqzXrr8mETYJj2c6nXcMu6zrSbb5XMw0WD/jlqRgR0
CprSemnXk2vYR68WzqdGiWWp5WqvqB+kgHUk2lK4GO/FvgaNfV6Y0+2eD7dUrvnGQOxlTfbz3MJa
CFOsQTlioOMk8YQc/3o4arPJqEwUaKNVSiuHyvLs1Zr4gJc0LmeHF67+VpKMShV4GB4vkYN4E02f
iwsDqH1h0k3+ei4Gg6fhRVAEk7DCrdpivjUJoXeWJwLwOWuJ9YGxSpOeWfCNQuji/T2WBdYBRyMN
vmmdYA1CwEb2fEglHfmUcyakCF5HGkYP7gbtHyM6eryfj8Frp9oIBI+/xtLwqGp90MiV+8z51uXv
DHZhXXcBLNF4JUj9M+dCmz2fuhu+NS4z6DkGqFCEMV1Mu0Kkfld/lrY08xe/PpLnksFg5Y9YLuVF
IxOMjKXFgZ5BMn11TjWfGHRAI9tiiWIyYB+uG7pRoYuYyq3pxp4scOxH3pCFdVx5i9UEy4/OqAux
GD3poPjDso77NA9MnlRdrXxlN+Jsv+cJA8ESkLvWDIwh12qvq/pKihXf+x6I/kmke7zuIBay0ToS
LLsGPkkdmrrXrhTQCaSSEvHqy5KEK5BEMPcUhZ1qrfRsIrira7dVOy1IgWtcHSEBp1v765qSdayF
JqWrDSVcKPMfVSDPUaDg3t+bRqxKxKBSQnkHlZUHvVpA8fN53Oo2FC0sNp+3nFhH26pi5l2LvCgl
aNG7c2XMBcTEMfxwtlfj5C5tG/ND65Y8z5eK6igK36iZsp7UgJ4tyPZ0kc54pcaw94aOjMK/b6xm
ywIkhl+1zjbp2GRFBwaSntW19osRsEJLNk+n20Ai1Mr7UvZqngCxWrtQkEoSNegOOhRXsv2TTuvJ
CL5tjmc5SvQ+MgZmzfhQZPY3J2aiUlj7dp5t3Pu1pl7TubePSkDcWo3DGUQA2/OnCdcjJ3truDgC
CezklYy/6Wb21QUmeMLC7RN2GeR7wYApYFs22BXMSfH50wSsM8ewaNVN2ERPmi9dd2ETPxVeXSvH
fMQMgsgcva+RVCGX1E6ilgqEABy6KhNnUrND6K1aleniXxI6MqI7MGdV/GGL9+N12M5RAAc3x0W5
MXhd3SfwwxHaw/QhepPhcRgtRqAmYjfcwQvCC+KwqTceP+dgJJpY5HwKhsCFLGHrsKMd7kpMoac8
T/uVpTYiaqqawUV3TqDr3FDeDvy43RaPCVPWyn/9nvn9ElC+JAD01zpNwRXUhjTYV3HhgPyF4L40
/MC+ltl4xG7/vvSpFHKMxKqjmC0eCU3Nn1LzGKnWEpQHgniRLhmcUfwbSPR4FD/pMCD/qv0yfv+k
vrjr0oNGAQuWIOVeCynlpkfLeGZKCQDaI4EKeQwUQl2KUbKqkbIG75oK6OSSg4SPTkleNkQPQF/t
UJ5BBaKESJNCEcJRwKqe6pUVqTDHND4vdqq+UBlixyby+8+i2+BtttYVBuunXvfJI7OoBmwnKO9e
sQ0+0q7YraP8ANswHwBBw83sC7w8euzx3DaKvccDkOrxZiKZkDP4CmLxS+a2YtZ9G3KS4Gs/ky9y
ZAlbihDnb4frJQgFo0F6yuhoWR81FIF61OuDxBuO44v6iPdis5adYr4G1Gnsx+Ond5NcW0ekmKLt
kEH5bSATirSZLmFhYv16NgwdutwgoGZcFju/0HNFgmC5AUrDRnBIxs5qOud1ONo+GiDpLKTXdBee
WV/a0sNqx/fc9dTDOAZRxW5rvuE4kojhnJ+xUIbRaJ6vKTbeFzQekZ1k6jzPij4HL/IsK/9vCl5Z
kagJeICpAUv33PhTDaycIee+XGtAFKpp+o3U9Np5rj/tcbzgC0Y9MgAShgloJmUJEb5d6jo/DUXM
ftYqKjQjzETsyAbtA1i41n4FQ8TTKpEnfjMi2g2L4h5mg9kZa8rPbVXBcsn24V1pxnTqnQfHfuPv
ChxGIt2SuUULlbh71gTUD/G9NpPCkpDfCFF3k6GNAhx+kptmDwlvXmQxA8ltnkHRCn12dTm5epTJ
HLhD6J2ZAUr3SwbGhoowEDvPgyXJHZqaVBMFBgDrsnCn7eyTVMYHMuD1awNpmSExqoddANosZi6m
AmRZfCx/npxNQt2jbMsFtZDUoIiY2VZVf9lNhAIqG6f4rJBfftdPbND0mM2oERGgf+S3mcBEbtt0
7S7hWjjB3e8go2IlBsUJdPwtTve+CsSPSo83xpbLgBzcktxVaMh2vYXaVOhoqU+uDGFmiG3c44Gj
zVQMtxwu3LAG7/+4lZcFu/t8CtS9KjXkqGOWVSs6zSOu1AeXRv7UP3e37/pl0j1h0KpEJCziyY+Q
hpnrPBUL84hFa3FOYEG5EUFFsv1NRLymHZt/hvurev8GqIEJTVcm/UoPThw3XmM9gUTSnjcKhxV0
L33mdbQ9euPtAJYmVj198ataX5dYX42lpmCAAKn+9wR+j5QgpjH3SnQ8mARLbQijAppW7s1AyszH
tYHmyB2c2TREW9HBFNwYD/q1RHGCbmGUXu36Mhp30Vb1OEXEX83l+6QjrQX7kFD268p3+X/DgwKi
sRLYO4YDfU1/jC+VDWYctGaSMfDGJlNUEZJXLjDF/GNWp+9PzxVuFZRcZOxUHH83cIyLPXHOKQU1
TOWSG8qCsi5k4USY6kkwFjpTV29mhruZH8OTF4Yzt0wS2SJCEEXdFq+3i5adRhVg+KRFl733VW10
VqSpobClKXmHL2bkK+xeAJ883BZSRiu9pb7KnBjUp1zWsmp0HBYTDRI8E43D4vtOD9Boembt/zt6
BkTc6ZRW2zkFX6MX4IRPLmbV2AZ99TpVf30UtR2k2qnrNEIWF14W50Zsuc4KaKi53Xg1z8WecNY/
uGkraVNNQHxRz8+mdVRuyQwyzS3OYsLQcXq2HsTFUPinAFfwyPV5Wvote/FM/QE8bCJOxvy4SLKh
yQDdXppZTKIO8mS+KSQwOFFvs+Sm7dGKyZB4QwDzdwivhDTuFA/LT6CgeRZFEr4glvKF2v25ZOF6
yyNmo0Z1qDhIYHwipbR1n3sN6fu9kvEe6B0WhCLz/j9eOssJnRbkfdXSbPntbYCHt3anlfyKCc6b
bymlSHBqXoakwJqCSscEsaZOt9KUady7axHXS8o313wAHbbSD5FatChaVtFN1+ryTfn+BAs85yEt
scIGMeBAblM2fNQX2xO3FUrU4SkfJA4Ku2lnFJQLZgWQLV3F+ILe/zy+RjdQZVoVkK0z8/whYzlv
Qy80bCVKAjR+Je2dPLN3AzdJqwSqfU8srChoYFMgykSKiuMLIsgIxFrn8saKH0h06eoHPLvCHEhi
BVKAieKVpEPqMftkfj/DT2Gv6yGhW/ekQTpxNKtdV+OkphLotE/K1AxiIUE4QoULBHGL8lqYkT9Q
txXlfxIfy9LSkJS0ETi0ByIXEGk7Kzvxm39m/GBXav6Bm8VB85H4TYcwVqe1pP6elKjtnrXK5KrZ
GwHnyy7JPohRGQfI3hrTg34Op12ModlwkVk4jBAbe93+33LiNjbUe8Tx8B+FA4YlM9Gm5IZmD0Bi
7LCg57mEltcRMCniUgcE9x1CsAk3AQ+yS+2uP/7juqYLhJOdVZS8p+wyprvG0Gp4Rwa/sBmycHdq
0F+7IO/CsUzI/sXjCO5M+H0as4TTC4hq9+4dCZ1Ufwb9E7a9FUhkYPFV8rKh2ABSpqvTqZFh4rlx
EJsLfL5JfOYIWbN0zVS3IbYli3rJHsoOe7bKfLl4Bmlx2iK9mpBnfOdjZZmfYwfrvo5MzQ3vgC4q
Ak59ClemJbCerDoVZrGaU1WhitwEUT4NmxZYJ0jS2HVWMZNZYmCkrq/LVSs6qasOTG5Zr7R30RTw
KiZsdORkiOWcZeD9NAt3+NpA3N8Z92oE+OFjFi60S//4v3qPtf9Ca8cDZq4y1kj4CryiIxPSb2SP
LOcbndU2zCHBXsFf+/M8XpNSvk6fo/9uUyO2BOfnLk+Lqiv/EgWs3H24W4+uXaiWUWnWIA+3ym05
nS5O+UzyLnKEFuXq6ZGRaS2338pgcjYfhSdCRN2kOuAmsTdaBFumqE9Prkscxx/XI7NU+rdPvvR3
nk3LiK9JpE6nUwZDNCuMLYbdrHlcp9n+f8xwntgDOGKmCJ1lI8e1QMuSEk81Zihd2WFWhM5mecnM
nNn1t/DkH5esy+zEdp8pXREG7Z+yvsCBDjzIyHL9BhX8BZRXzygY9PEQl8x5J5sVxgCLmQAdA3u/
ohWVD2J4lfuvMFyIqD0U71bu80jKAeWWgLZ0kvjrlsTLBQrvfuYspkj61/HVItbDvTpRlm4DDZJo
hY8+aFQrg4406MsdJ9Cn5drOpzRdeNrjMcIT6AHvD9BwGk6rrBfKmc/PqbdZQQFoDEUNgq4VlnzD
LvynPWNUPnbCKVtdci4d7xmgPSOmvpmkbJ+oCYPjl4QSiG9guAxMre4828GqQ+xF0CCyo/d0qcZr
Dn/43qf7TxIy85ZCVG/S5haeepOEXA8YTJVhA9yHPPaDAqoIMeAcbBihBIKcxo/955uKlPlUMGhG
5RAtSZOMdpcRuo603A+Z923UnoQ+bKXZKkJTssNMjfe0FyiicKq4eJlQ7o8+EWvPtsbqEM7jDgWt
l3ZsT3rz+kFYcuw/3cxKnUo1QuswbrrkOBB/y4EUU5bD1SOr5puYKmknNgl5kAdwnmhiCP+KsiYT
JwCVHaxVs6YRwISX3igCqc88qbsAOeByeJrHZy5o/y6aCz3ZJ1psNjmdAMfXs3cNqB7yKBkZqz//
cB6fe3Vi6IGPpAsh1BrXr2oZjKcGKF99bgK6aCDyU3XJf6kItKopsPwtK3yJfxbKE3G8R5U6ePw9
zwc78WB2OtVsVaTfabJ//JWPHnA4R2mYprTm8rdtC/Gx7zLm2gXd4aTm/GRAWtp24ycV7jVzfQQ6
1yWnb0truf1l88uDzoT1rFeJO0VK/VwuqiIdSxNb73oEQJmgXBknvnTGKnNfXc05WwMP0pDFKGoS
4RsxQC2AOfrDeRmXSkk2VmRI5v3MA8PRO9j/zkfWgoYsjESlJWdw/h/Dts8AFVQ+aOuhBQYTZzQ7
Mr36iwW++b6tRFasfEaUS4wIFy0jT1O5qEQyEy9yprcl/ybmJ6V3AZGRbtR3rR+fMrGKWGaE2P6h
Lm+NEq320jqLpv5fzf+vBHrGrd4NPGSkcQqAUdSgfgq7OurCzQSz6I4EvQ3EiYPpfLAVrYQJ6C9y
jQha3GIDmevc86BhXGjp2YfEO6BogHVVmA0dE9Ro6yZTQC56Zab/xTp0wHSLiC6iQchM1hm5kScO
5fI8H9oaupOcR4k+A6TdCLl2149lwmMF4eXhmrghdth0/75lYvxrj2sA8BIiBauHypq/uXYyoGA4
0cqSQgVMgvS/9ObeAT1zmQJxh1lGoA3b+IaP9oDnCDQUGOTHKHLX/PJloMW7LI3kJ1u/41OdOUMz
mAi2AJbZKjGx2ZhvDxNTslP0vYAhN46bhrHQzK3bGaLmC9YwPRrGIXrMmgsM1tnFtzOv5I2Ww4H9
YIs76sMbSzCaLDuI4Zfenxtuy5+deJRNHjamrGTNQELbLe4pUC6yrb3tHJX/u9J/z21fU3uCDC88
7DtcPNe590Kdi98yu4jnIEUptAwTgzFWRH533YYt82t1zH1qeF9L425zVwZGAYhA5s7VIBFw5D/M
L11V5YTQeKkzgah/STS40PZ7Hh5t6Jttakj1+R2sTu5UOxofS1Ut35XRKfeJH2SFqY6bxqunuL+k
lDTCWqgZhWMLWMaNVlaWKaiaG75JVcB4Sbi1sPAwo0l0PNFQll/JyJ6/Z250UqCe0lsMVA6r5/gh
Zx46Dn0bieBjqobkh+OdMBaLLFs70heM+mnD/dxiURJB1JR9QpTNmf7K4adDWF63vUaXOGDnp9Fa
Z3Jrw/ZIj5MCWHfOwcMl2lvGB+PeOWksLc0UYIrt+LXAyfBmQ5aAk9sBfxIpOcVGraXo5iN6iO7P
eBT58jqBhVDo4vsEB9ZiElTawZRC45nPPV1uX3jdJVxImu2kplHJk6JuEXhNMMv5/gbCM4JoURhS
Q8Jr37yUWgsWBYcmTCN5Y9LHw65rH3ZIywSearCeCgTuwtBxs4nBGgDV3HIxdbOV/YG1jslfqbP8
TexfatLnp98q0q+OzdIPeRKugc8bcN1Rxw3DFEc/9lBHavRUYyyIb/lS5hAFpa1ELhTPMMzLC4zV
X4n3RbyrLHqHhUPk5wMsuWM8b79B9IKQtlQxGxlKx774iFJaoKIuwfjZGUY3QrVVVtMaSPClRoC1
ZDFpVqnlxN0VtLcApC2fJ3MApZZT+1a7n7oQXOUefpRymOWXzmlc4MZu6vzJxvxksAYrkmOLBPP6
nEygYi2LVbc5YESbH2j6K8BG35v1k1ZKGSTHc8i0d12LR/E53s2KQIXvIVSOKVy0xqnuAwi5lN2c
5UwMdPHx4GYB8SnehHRgp/j6LKva9izx1s9ZEimgXtIUJvSUNdSf4cjWa9stVExEK1tk7gJVqnjU
YWQSGPm4gCBxYDOdC09+bxw1mZYGOozN7mC0HDw/JwGvGZxw+z8OcfAiiiFxLOSmKpa5CNME2Z5M
YkXVK4/xcBosJ0H6MDZfKd/8ur5NFanzXeryJsQig4bAmvWLtGTg5D2zvWadpVWG9xx3uDUaDI4p
bOwWwtj9IIiOzkqOfSa+G5yCtPm9DhjL1z44TK5aA3cAo6yTXuWB/XUpkrPVPW7+nDH2ndajawXP
bqeJo5Arq7oK9/vmdZFKhIKN85tk/9j7/uXnDYaIH6Fin66P5NKtEGUu9hW/AzuwMdt6S7lyqXUP
Jv6BKUCfPrk7/RXwlk2xZhxsuF2hiVIRkpaIcdc77WDkS1oUAirdzsoU0pBZ/emihZlONxDwbhzz
ZIa9Q+WtyMLk5vAXb42n+Mc6hMoZd3qXycR4bahGU+yLfADpBKVf6B7HLFYXrdOFhvt59cs4t3nF
Eb39f10khEWwNVncWcYcBGICkT2Nt86zFd/8jSQc2C9xy3+j8vDCWQjDpLcXDKRNudajl3ZBbGE9
CFYWdk5KP63NB4sVejf+8sZdFG8zycCec21o1X8Z9A4gQnK1KU6stbaSPjDYJW2CRu2G+WIG4JI+
x3FS9eTZ9sCqFUBp//dwp5sTnmGbfzK8BHzC4T67EsnjY7CfDOR/APPPC/EKOCoBRxI5JzocdJXG
gPsbRV5AkU8ecDVqZjsZWIICKkFIYgUSmQC8plsMoVVQThUDfBIGuDJVYw2IbN4EhDVR1uh9GxZn
Ej8ArVGWjZGwa5OhmwQCHQjAFKRztRH9/vKgzPgBQ0BjmZ3UpTN9ml8l5WY/T5YiofGcycUR5dzu
heYClcfVP4VOLL2l7ff2YASEygg3kYMK+OB1FBdQBNdhr4RRKlpwGyJcjWey6zYhr4GGJQSPOPwU
IRSUsZ7Z0d1aKDntvmNkaduK0sNlWe33c6J7nV+cxZcqLcXXolgIoHibg3Ymx/cTGEMfumZxoYJz
BXrQkTRNJLjwl9g3iisLXyv6dn7vaMn6fgUV86h8dRHn2RdJJ5Sc38w8PYYt1aTuDW3joyCDBcJg
dKDXt1eBc3k5H5vRnf0HFis0y0qXrh4T8ZMYH1OjUCjjYKb0eFuLZkm4pJMEfVCQE+Gv9T4rl5YG
/wi4Wzfrt6cIh6JTrZtWRLHB2Sb19+ibNlbjUPntuVxY8337A9uQd6/fU0LZ2ivpCvjhLlMkbIJ0
9Lvk5Ec9kaR2SljdYr67is31FKELsgLIOgt43WVM36OVAcH7Jtx/AdqnqtOAam39FKacO7nwsJ1r
KD1Wc0b3Rk0EAtw+2l0t4+dwSdvYu6vJALGZVyuCpIsN0sR6sHUCVyvmeV7o9df4PZIyIcOe/Wjl
uoI1isdxYkFa4ir6pnE0DN6pfByiEUJ2vJYkLwZi0JgQHvIOardKD0KTBKzjTEgy7f5oKiXgZOrx
UqOUSwuufzrbWyInxG7HBAsLwXuJtsK2blVYQR1WxLKLsSWDqrSeJDKa4B1LrosSFTjNLVTtd+fT
ZRefsrw+/3v/QnKxyJQotZPsxRSXExmQKhfUaJRKnPVupEEzg3zkPiAaK+vzGRMDyeHpnp0IFfL3
6fZaM+r4tglJ7/yKEDsSSfFA0XhWCv5WYdIa8jjoOLgAVrSzv1ndUO64Rx+y+ta3IWKvkzzOXzKE
GxicJ/QRqN/hdlFyZ7SY1Sg1go0uXta8373VHmmJ+HUkg/V8vGwMqAXRtx1JpgdzM9dcNWQQbh4Z
VFdEyTuWoCvzFy9s5xybI0m7jn09RpChZxmndZPukvCJl96FAhbc4G6EosKLHdVjSupgLqVOOLts
470eXhWDrH6n0fOhWQJPhpkpehfhOCPKDfs0p9m/UoOvG1+cRxXIPurysHU5IholVx4YaWrRXNCz
W9WYfwohmvGCSPX0USk4gsEAYXITE79iNX/h7IZpSNBh4p5OMg36SfOsfIujh+x6R7tmq05JFtJM
QUWGoMrDhK21iqIPHh5Xkzc6R+FKr15PPOeMAHqUDDXBCYpYJ61VSI++N6BMqQPiDLefpRbisviU
AcMzDKQFlcGiTBjUl3vpmgr02A6xyzq/o/RNYmS+mmRP9SHsQJpqoD1Ls4ebLcO2qNgwWRY8pwJ7
LwRQN3ulHjHtnZvqetBvPd5fll2V5rTM8wTmEdmsBbJpWNuLrSZvc6bROkM6Fc3oUm+BP3eHvEGc
cxOLOVocz/ixXafIghRMMTbdsE9u4LZvQlI1JzZLZEUq0VxDp+LtnGjYFHzvTyegclwcayGPwG+m
j3biTsbhJK3i2VWzy33qkWXARbwW09Zido+kCi9M0RoqtaBajiBvC5bz4x0giz/Ql2+i4WHqjv2u
aixz6i8RfyVZVKzC6++dnFKC6AkC+xUhghNpIQw+tIGf0BF/3peqvED+o6qHOZkoBakA4qemR52m
a3xd/OEVou8rl9qIPcM4yD5zaGe4v8qHcSDh93xP412bmiq8KDv4yBqY7qHPnYL5Zft7+glyH/0n
AevJfSeB60PsCJ8/2aijBDLD1WKPviZzcZ3f4DqVya4VAXgnibzcpqGJRZQHMp67jq9ZntSdHaH6
Wq447ARk6uLtEFlXAopRJWyre39fQhQuAV1fOGlaxfwmLm//LGcslGKbJi5Whx6T/kUcEn9YX5o0
pRQFAZHMFjySyjRIuPRPD3fIzG73RxtrbTtN/4X3S+mazl89uKIVnkGeIJN711oHBLUmRqcBys5U
yVB16lGIFuUix7RTJB1LPQ10ujvMy2cw6mYhl8tsj3ILTM8jVVzpIDLdYFcCqGIPMHvc2a4oiduC
lhy7RHMdGUrdqnmyyAEzOqqG2pd6xPbuqwCOLFORXLwXfB7TLGGqjYWZOVvIGRJ2arKkJqeH3cVR
eg9UG0dvsmzI67daoV13BMQkHpsO/a23JkMXH84Bbe43XDq7NPp4i5koklID6UPdZCoUvoAOQMer
PmA3wOZN5/9cNEZDv+Ho6Q5nKre0Slxph8Ll0BpMF21v7Kt4a8MZ13wFpiwmGg+7s7q46bTL3TFu
7jJYmzb5zg9qNeuN2kCGKRuBSXc9c6SfVoRLaIbiXzLRwS0peOwzZPk70C+VgXB8s8y48bnXUeNc
3FKj0vPEbrUkMnzDvZijuhfDeK62UpaIpdN2lGcvDsrnPLx81Cv1hTGGUUVytDvZQpgJXbiPTryz
g+mAcZHsYSlFgSk768P3ie5i4ZM0PWBfJaEfiPTA1R6sCVUnHXioy1eScSgYl+AR1oHXEdrwmtgY
LhCPaCembZBSunhX1nFjXehgdNt8VrLawi1QGSodNnXwsHMkjx0Vw36crbMPgHUg7O1Q5zKRkFJw
z/sI2xTS8vrB7jDZxaWe2wvlw3MkesiAvfuJ9Trs7HRL49XBS6I4mWTpFCzRXA4o45x6on+EYJld
UL5UQbJKrKWB3HB8au1y5Lsd0UVFcHnI362bPoOcaKuWMAN7hf31KWRbjdfvhu9mhTtKloPUheq+
PiPQr+uLF41fCAqEU7c87W5hiO8EGzFk/jBKmOna+O6smwEy6KMajOhX6DbQ+SI3VdwTTRpRX+vn
tddvLw1mLu4a257XcLCNcAJ1FYSzDY53BvCr37cvPRNOJZ/9CuyLe30EV6tTCeuM5fntzsKkLLhF
75WujGBVJb3Skb0tsB//V2Jdz+agtmFILFjPNhG8Bt1PhhaxkubPhHoTqsJ/t+8fFCKla7cYOB9A
TkNtj97NGCvQ9fuCwL7g6nuuOsr3uCbYfqCd/BWrIIyXO2YUP0GvpICs2oN57/OgKhSdKhL09HtF
RDQpFNN9eHCyF+PV3yG4FSjtg4sttYZsYIa9rzXQffdNndbYKjKF4hYPFbwcRokMAOapn6grBT0C
BvX4D7wM+iwnUocSxuFmU7+rEPdmQUbiJYuwD0mOeqyRjItpudPndReiijjE5bLwRt+Jb4UOZF7c
xcZMxoMtNg7AaLJjyWXQ9wBk9iRrg06l8lv4lPc73wZQgek9PKuNRaQRxNkcV8X5/ee1T3N3kEcO
OyvCgtc2xVczxom0mz39+K9SSlL8ORthQzQNeze4opEEa1Z2ds3jVIjYaIxq7ecCznyfc+xAsIRo
weUV5fOXGAd7PLZ4ihyGX3jmajP9kpgA+x0YlK67Ef7AttZZ2p8xwlpfaq4JnGsckFlk5x4fMv13
yGGA+ed6v7DkUJe0eWRad4GqDDx8n+GwzGyzG6IWGK4RRVxozFM+8y+eUl8TeFnscxJgdYpChk0J
f1uAx1gXVM8rxE2H9VpWPQJ0HS4PaSkHepnODnXCDyK2y28es2NlWgeq3ScQHAsKmR9VmxXdDPDY
YKWyQh6M1D8mSKbJcteo3Y4dqmzc+ns/XfnoI2y/KUzVfhZnYBvWEDWH5Pf3YD59ilpMqFGrhJLb
CJdJv6x8f2oiChqZzRQJb2PFUP5d+z96IDtStUPUJjIvqIIMyzrLMyLU+J/dC6h61HkEA3Wkv1i1
hYl4XrxLLBZ1jLEzgIR56ClLRkKQjw9h9cu0F+1r5l8PET3m07LaGixu+aC/EXaKxcGG0ms6YWVx
oK/ke1HW3qzZyElX/CWac2IlQ3FlSxlf4o2GX6hcHgbSmxA1ydP2QyHs6sn8NBv8awZys+rpZHlS
LGcEizz+JidbosyTk9Bh8ySJMV8G5KJIjdC0j54piA2XBrUAlVL2B9SJ6Q3owvSb4lxzVPLIA93z
cMOKzbh+z0z3v3R1QQqBbgB2gB7lqZam28HtzAiunKypjvBbyTJWv7BbUebKn+48Ar3quwJHrCAs
ohpF4bdwoAxwcnyALxaxnqJlyAHPTNrErMXkiBp8ZxLCWK+LxSSbnpQZxtP/NlsJ9iKhLKtEvw9c
v3mo4BngvxGRjCKbeTfv2gibq4lBhFMZQInzRgjDB8Ukvc62CX4PW/jsemy27ov0pKRf1Q91uPLQ
sMV3vRQDAVWJ9AGPmpCoah3sWXmIEBDedL3leOnj+0dYo0tb2bz9nw43SPgyzr4qED8EElgRsmbI
5pxUBmVXAsaB2iS2uIznUJH3pk1NQeWxMw7Rv3hLB6U7+64iF3NagMPOfpABwWNae0fDxNN+jLLo
TrsYoCRfL9sSqjEOxNaxKWZZeIO1AWvuw8T8cFe80NOd81Z1+06g+ClvKrPzzy21UbMw6cD3AjnS
/VYbksu2ZaDsITDtwhWe41YxHyc2gthv9PwW4zwmCqQj6dPN0A5R5TFtQs6U5RpGax6+HW8pZ4w/
Ypds6UeweiUR2WKwGK6pa7dl+YD20GaQhGhtnuQYT1WQTIn11PKDFbrdMk1+Uf3vmhAqWX+fJrM8
6FKYOUSFhJse+cLKGN+E6C7h0t/Ii7ZXqS1dbNL3GNlEdt4LuJoqhcrbWKIbggcaNv0tRJofcZqG
/+FKWIgThsKmcEDe4hzFslazeOF7gWNgT62EBC2RqFqLXL8vjgVXEyj5I0W8jQnywOqTVsY6Tv9u
GLO1yCi0nTg2nsjYcEaEpYSqutzKXLQM6DQfBlkqJLKOwLHDvjtjCrtGLQIso9atgP9M+GUJLtW4
OXw4wTcgl0zHTT4c0gmnZMmBA29rVQXlJ7n2oeN+mD7Cex1Ik2Zkbg9HnH+rZEhWiLpkQEqSPH89
l0IIAczEsslFa8InYpiDeU3rif8uopJOyCZ/UPTM/d1AHbrcKrJkEAW/8YcAfKlPz5jdBHEnmvGs
H8SG5lOStnRXEYaxELVEV8vMN/HwGzYlMzcw7SDr0r1vu62bqjiWlQmLnj2WGNUMJJAmKqC6gCXx
UaI3EyrK655wHYgSGKeuleI4jbfsjcsKTKdZstl426PJptXi6Z44+qwNaU4hsRx46mDGoRT43VYL
pcLx+WhzSkR4aA4f8tKPGxTicDp+pQNiTOxhu8D073mPe1YQZ3OBq4D4QiLWGNQtrua3ZzSAmzom
KeRpEASRg5oNodEB9rEE4KdHunh+DBbD6BaETt7nXBoByBPP/eVdHNoFzs0hQklheeG6XOWi0TSt
FMHVk0sF8atSKF96l02B1Ton/D0mieMpLbh2LFgZMW6UgsUswQRG3Uyr/h0brOmnoeQBTSz+xeWw
X40yff24Lrsz9TD0+6EnorKSS+OizIXgDrt03L7X1yI8nu+tmZFC/0UbBb71TgfZGDlLYz21n2kR
pAvqf24hy4wKrY1Ex6FS1IP3gLkPUXcMKXw+bw4BCMX0zJ9rCsE9+fuoDCcSTpoD9CwG5WsttY16
3dWWFRLaW7mLz4leR92xEko0KKUkQxdGls1brNAhRNDP6pQNG8/Y1Th8dVvGbQf0AVrLSZD2AGlq
MkPlNTxNAmIhYdzsPMjQxEgB37VNshHINlq086d2rR1mhUPXr6GF+o6qOOqhEqwLipcQrXizO8O4
vNu4TV4N/RkslQ5vUjLDTUzm5e06vz+i7mtkvWK2n4yWLaDc13PgMMwqDOrB2mCVrbHKRcZqcMFP
XcuuEEB4Flo7YNb9s2C8Hm+bvBlP6xsc0rZ2YJ0XFF/whXoKGVddmd5VB3k/Wxo6X6Ylq2SPlFO4
hujI15QJ9c1fwZuhrJt5FpATp4B5RdRgQwmv3UHulqzpzMZookngiCni8kqMDo4nlZRIRd4XQEF0
E5KK7fdwEyOt6Oq9qxjntlbrxFCg1q51A/cFZweSPQp9znWszdDxjscZ/J6bya6jZmtHmWDNUIqh
bpaM/4tt4P3A5OR0t4hYWHfUi81QRO1dguR3jDTZTQZeM2Ohhhra1hjRBaUuKye0zpwOG9RJYV+f
XTYrUnt26TudmY3Mzt7TcVYs0VCz4jluFGjOACv3BFURSskywl+oN/bUsGX1fr+LVcTjmCcxMZNQ
ozZzwHvg7PjHX3tNFIUAUDDVJ/tYxW2stn9FNFzUPgobfMXAwu766GDvqGb4ywEVgRRlO10S0K5r
re/HXFSROlQ+N9qB/4eM+7T+ft1P3ihst+U0mA72kpadFO/OKocPAVT/5P+uj0zapH1h8I5ZaHvr
v/b9pfi7rv9w6xRqbau89gSvB3YoIbwQxIp2uvfVsexPmJbPVf+dIOvM8TgXNkDsSl7F+z6ph0S9
jyJTaQ7K8aNXg08DL0IDgLikWy+J/TUDptPHgdKcs8/evXfiAwQve0VVSuRBuvtU2VMxmRWgd2rT
gbny1yx/9wTrIV77OjDnR0UXbGRPYdp7xybsiBtcNox7AbZrLNs6MvCBmf5xuH92AWjk5Z4udo2E
VyiPCm91ERA1ozkOaSfPCI0jVImKH92f+1gTVc4pCtpCuzUMwSyfuq7zqIJNCDXySLPWepulnDw5
T4YtoGeFiPpq4yvoeyArsn8Ea4B43zNNu+YE35bZK+WcKEmlhAAuChW36qIw0ws3jpU0+ac0PqoX
3QPFv1AmDV16DqfWW0aOzl4pNXUXii4jtfaHZFBVFmFQuHjsNItUZ0+NiI5PXogYaraG5tT/l4TZ
0ECSRIv/Excji4YoNSfTfQK/ochSiAoq2NAd1wF1l9flcy89g5xPj8cQESR/wxOZcIJ4UvPgZv8N
0DnJ3btetZdE2F07yHx8mBxRgewRpDgJbAs7ocbLWVYNvhTPgdhJu3V+JUKjJa6dvuZyTx9E8k7y
A25SjHx279nGfa/G9HSpriXwgtO+JmE7YbhxHSdICR4prKtfXqqwOxCWkxKRvccUM5P/p7AUG3Mt
mcFuRuL4zvrUFRlQy0rHUS+gltkUfhTrpiL7KZHNY1/pXlvOgxsR6VJOllQbXwe7NMT5gxsoj3k8
P3CiPljWFQk2GEmiMSgIZtU/b+m5JEr2et0ljUPZ8MPiuys6Wrmhe9WgY8ueFsZoY5jRIrm8MGNU
brkhWJ5IfHIvNvq32I9RQwa6z6Rj0XRTVko0Ppxlqu92/H74sQnFmEXsbRebUDXNkPh0n+uMPfPz
nZeZyXZW5wc7+UzF0evCYMWwUT/VsB4InANWRm+VOsmcAYBaVP7x8WSfD/8QMS5lWEwRuCFoToP+
JTXU4iTML9TOpmWC/VAZA5B7VSr63VXIh81TkzhzjdcJ7+uya7B/yiTOfjFyfnRNzMAjekuhp8Wg
awseoNeTdoHgYUUn52r5Ffi0m1dxS4OtZf+HcvKzvyVWngm+nW32hQjeMx+MbwPU+hi+5uqwF/sG
hs4xUDk+T39ZJG/XbzUHoP7/8M/NruwuCnG38WEg/8EMq3TLJT8mouIhFwtxwE2mJXCJaVWB/5/a
+JP1oI+B57pCT4y5peC78Zl5SQM5NcGhxe7LaFVPpaobCwo8p5lxWS/FkzJ/3BGPFw4d27WB+rzD
ts7embn0fHOwVDw/D4mdYQQpGVTHUitGCaAYTbojgyUu8596pkKeqbFude7JWGeE228HcPqUGtYC
kU+x76rm5ANHXYRM6dHWOK83pwBOMmLoOcxxzIDjMmyR72SqjCiIYp11srL0Ye2bDk0nEelUorw7
EzAE6ee+FHcrQjX1P6saCLcHgdsAoxp/UwJIk0frsKQdROsFOdDN2bABs5F3QHVljWOM6Z8OIGgw
Zncs7jps7tsjDLLsgn2nuetN3yn2upfonRFAi1/N3ktbY/pZLMW59Pz0U0bIUzPppt+Z2pY2cl4G
mTw2x733oMux1pMkNH5CpKu+fzVLg6orFna31zClEdJEKFw6Grxm7g17fpfSQV/mg2Oc1lIoMhIJ
cutB+0B/Yy9K/tH21Fui7PtWBEzjl/egoAnKyCtEfmwg6EOEGSZ9VThtuH3T9GLXnoNFeiLF0VF0
fEt6yehBGUMjv02rofl62U9cdpoLEQlCyEKbnCrcDO7KflEUpPb8Xis8Dlqf6aVAAOTSVn5dzdDo
7glZKAD9x+3+GihS+CHceMQUxdMVJyaeD5Z5P4ZIRunOsORW8ha4hvTKDGLHCmieS0YlhAxXu1j3
qG9+axd2juoMqf5Kj/7O+pbgrHPKkh8xMRroDeyb2gQlNhdD4aGOeYSCYoPISfuyCiTZIwbGIZzF
BP3aJtMhQ8+F2nchnFobnIL7MdV3P36HuVkeIJaAw76j/v+DCIfbSoGlNCAq/tRn5Uc2px2r9Fex
v9Ik4AGqFB49DjHEUR6lJ9lURBXi1Yuj4HNTJs1kqXAYRZhpueR3KV5tomnVRUYKMU3zg3vmWFZd
Sbw3leUmucDUiHqIwpB88RWraM7VUnnk21ltnv6WaUep08XcBm846vXw98/GeYSeR9qnSFHNmwC8
4TAgHMJcCZha13iY899UDvBHX/h5LeSj0DkRj9pfa5BMUwrj2+YGofCssxHUpe0oEgx5NjxM/gEI
19KPw3aG++4l1M+HxJECilS4TK179tmATct+r0J8kBbqcBvCWBspRJPjfwfHuKXwi49LC8MlI9Ic
BvC9NxEKTinbA4TOa5kGX+2h/5uo2yoQC+lyeuDPsqrcXb1HaAUK1QnTn8H4y96WZNhSsSXYPcQ9
mdHbEnA/CujmpTN6xxRqQqpWWB1zbiQ/CKlGWVnwzYZB0yNFxx1XUnqDDXyqGajT19gBbsbp5ur/
R4xVkYWq6mQZHGFhHiZNTfeL1E/OmRh9q7xr8z6HKxRFzLfN4BYOoj4VBuQhw5hSVt+PxF9cOAV9
W+vTVfxL/MvyoQLH5fSzoEvNeyBq99GkDwHCSDogecvEd+OcbW5mKWLX2tDyCSqk1oA0dsyRJqWo
w1zq79KPdmUlqzD9eZGDMwcU3sMKBDsDZsCWoTlHeBMYb0aXabE1sEiNKybtrRZtXlpgaAQjE7gG
EMGmnY9jNUd4+N/ULlBGl5CE2AwNt0rHZ2Nye8MHxjeRdfM8xckGt1cZPszw0Yb1cWq0wC12CmwI
PMQkCmDjVA8nCWlSaUAfhSt+t01wNR4TxLBpfveIjwY/uCg56j83qc4pYCR0B0T6SgwMIZn2akB1
ZEBbBnN8y35nh4TdY8EdDsC7iIDTf8DrYB732zbNo7r0fZy/biTUT9wvoV3SVshCFt3q1ypVFJyD
Cs3OfA+eUBOelx3q3Xs6Ff+xaykYSgGnNWlXMadCBwEtM7+g1slUh8zoVO5Dqv2Ir4dd43D+7shB
QFdG5gMvK/+ZtttYoRTa4YDfpg4PJz4GIO9d6qQ430LP63aS4V82ixGWfOOkQBbqFp+hYCWKkj9V
7bu5W7Ulogdzw7m+f4U2PRLFXhpPJWnREPGI6IAh7vDz6pQKt2NYTJiP5ef+GUK37NUyQxbSTiVJ
x7gTlR6d+AUwExxM4DS7tIbfg4PDkk1eL+Kqhd96rNpzLy37pAVy60z/L0fSU74kHYRXNkpa7AYu
HvLqy6FeO/0RzoWWpLK8kz4etRVGxufxQzUoCpeulP/jDFT5bGuc0CcaSahwFpbd1cyhj+icIXJc
G5iDq/dhowEG/UfVWegb9J+j/R/CPwEXhoF1WrM46JB7gtlnjWOPmtio/twO4JfWYfKPKm2UxNap
X2NsrDD6rbtGXc7dfuNcw59/kcrbNsFk6M0iuJ23WWP4QLCoiXQeb7lMbNXdmbRAj8vgBF1Cf+F+
5YMaBdVbN5jw65uxuz4PczPFTXjWmzsKj8nz4vsvZFhjgpLJEOCqqCam3s+H4pCQA+WPGUsOirlO
lTRBGvCFJ1yexTrDzzkahSBzYxEjDrWnZnEmf3X3yrsAPVtG4HqGbm6VveoifFTn4StT6s53joye
fMwano7DxP1fzDId68hRfriO8hojTmhrFgrBOYmhMm3BJaMO4KQwAEYCl8b5Op0o+ftWw3FQp4jA
YCcqZJsq4+kZeBgt0rOkOsPD/AGHNtp4nAENRvp/ITK3XxZHttdGQiDlEmoFMQOjwmdg8eziDLar
cVuR9tYbGK0EcEB8TazWONiTjjMPYK8H5KtJKcpxSDw1RGoq3mO19bNB932Yspnq84WwxLVO8M+W
yVE/7skMlCp6tFOz+KEoF3f1xGl7GgyKJPtZIebWmWLOlfdUqaEVcaTFdv486xO430A/Nx0pj7Ql
3TksOOPldgehm0842lJyCNtu7MxhWd1GnywHVqYDGQmy4pFMhshu1mD961vFyD3dhWqoPq8F7C7y
+HjTK3kihA9hqykzYDdBsvP71BbLPBTha6BmpgJ/besnZXKh9xk135yJ3gEFFugMeb+u3yJb4+WR
N1BZHRu2/QI5S6SYLZvhpn9JGDNCHE5GyGAV+TI4a156dN3Jr6advBFM7SHNj7RP1gdLgg/uX0iV
OUqKJadzX5NWdPSj/fndbBI7HKSumI9lhs461STUWPz2GZIPoVT1XJsDz4FzVLU4sbHSMj6zf6tf
r8v9BBHiOW+jnq4cJcOyxLao26XcxDo27LFcRPFWixsBhvCh5uULRLY2z8OuxLlqA2arI25Exicb
5T44G9ID139fgnuDvN9bXc8NyzXlS1O1uaHMNe47zDXjYUb1pNn0+EkVmrzCYHBYE3oaJmHnoPU5
TZRdtYQ6poVmgM09BmfqvHw/5yNWdGHROv0r21TpjtxgqOBNoZCNLTBlIva/s1YDqx3HbaMeiaKF
pIhNAgiymYalzkNWTvF+XC/FC83UiNzStoYCNx1f6Z/64HA0DnueFH13eOlGKHHX82o8+K+PPiQP
CIxc4Bs7kGQVPNF4keOvPWnIj73MhiaN30Wl74NxI9jGTumrL/cOhUBL1CWok4ERMykghsJ8wOfy
y6Lm2l3FYHXQB0AjCHpRiShIkBJn0ERiQCvnCt96IvgKJre1DyQFtWc6gC9yW/KLR3GEcvoDvv3P
G+6p/IPhHfJtUA1LuA+g054CXaspuIkPhZFs2Y8nnjpJH2QgrprTwC/czJWgC6yMWy9e+TxQ+Fex
oq1D4EsCvUIDsh/jyW5O6vOEA6bna+QFlhNertlpFOGrgozK3/HjGfHqKXW2A0OWJAoFHmTdvGrz
459t9ebiHjBX3/Azs3/QHB59mZ1jE1Uwlcu1uHjUPJr59ikjq8kycQz+D/kKpMg7ligpEuqDP8wh
3e/P9wUM76bxFGXsAKqqfFWnFvM8qXEREBq7daH3L4j2zCBbd725eBzufrK7xFKZ2uDQhQWIBFFS
NyNyNNC/P4QQBjs64OsV9hb4Zgmh75MsO9NRVtznnfhXvXuiIal77RyULOD/8RFpTQjKVuhSk3Xk
05pHQESyKXQMoOn91ZnIliDyjoXfNd0MCU8HF8PpE5GxYPrlPtEdTFKeXCs7a9LlxIArTOGpQt+7
28tkmEHedesrhQH8GIKjp/G6yb+PWKWhI4EVlqEWZ9xgTRFgN7KUc6U58+p9evnaTOx0WQEre1Rt
P1SWiizwvBKwAnapHYj3lwa4g3HTEzviWq5n5baPLQAeswIlMfvfwtm6+lDUcpRnpeA7qlBIYNo6
cSYZV1bKB0siDA4K/Hp7OifbGnscUNhUD/1Yk2NGB6MkLlcTIxtnbeQR4RrnEG4pmOYCa91lvPMY
jey36tx/jFQvEXdAoPcEacmAiYmsEIWyGUmls/HcXci0I72SgOtlVsVpfXJNaZ+DY7P6hvl5T+du
NXKmNVgDw0PIt/b4kNpdanGJubWx0jVQPgwAWyEfRPGpM3wcfwtVHrdxYtyloUith60aaVV8Czt/
VR0ZZWzyJec9bMrRG0QnMUaeb7RqAIYb61xdXzP4a13tVSIVWjP/VP9IYpL05UnLvWbAz1CczwtI
6XaMdD9G30ZGhe8Akq9UjRMuImL0+8eQrf3qhblyhtxeTL2uw4zGqwwzAKC0AqqiSe3NoDfBE/+M
fepbO2NggQC7NPvoIsH62Ih2DPDg3V1ZoOL7DY6K1bNgd2apbqKLY0CS1WE36OeeMmkoTKaPr2EY
xZT0DjF4U8bJPcND7dNHVSSEofKwFQsmgtBOJbCFTRIyjIaBePPnJM5UeiQIKiBPIT5BSDSK7DMX
IAnCB1K0CgiHp+K9nMOCG6Wk89/J5StTQSUcohVyHdFO7Yk7WlQs9PbcOXKKxlQ1/gLAQrIbglMQ
kxRgBnKwHHfLqjTlvw4OmUi66g7YIR/we8UEAcC3HhlDTcluRYz84RdwdyQVtw1xDTEWetvYNHNH
3GOKWnKccI2RGJGC9YCh9i+FLMYupo/jSswds/u+cB1PmKmnjYzCeoFZnw2UFINpTacrQfPdkKjt
SrYrYAvD4LYUcrhsj2/LrBeb/hLuyMoRnnxQwPtLmcQR7GepmenK5YBvesC9TXL5gH4ldf7Umu/O
5yBqHy5yj60IqEYd/7mC/cuPTIuZOSEjb9BfDr8HP6VX+f6gskyC+fSasljfNs5w8BgLTXKJ8q/C
yFCC/RQFe7s8TY7vRq/XNvCa4OoAzFZTmlml1qdWQfY5Cf8fZUg6o7i1XvAHs7g8Qxo6RQEPQxhD
pcH7eRWH6+W8ZlQCjuk06rgpRT7fX09kkhX++bKRblDVQhAjMgny6ky7YeI3YjUNJakVbprgFjvk
Jmhbr19v/NwVzeBhKq97PHiYacJ0ST6S0pMu8n3ZWkL2kkuy1wWOKWO0gJP6G1h9kQBnHjOVKdB8
HdmUW5OKjt5Ev8JY+sJG3nsg3x2cRVDj+XwKGwDOLYPnro4u51UrRreJffdWzLZ8e7MyByPhQWwL
3jdccb3PxgttQH0CqC9SR17dojCKrpfZGryplEJgBWhM9Wf0P6lVXD87cXv9xZQIpTCsXhcYUq/J
T0jfR79EPuezxfkSjtT9hdtLnHUuQk6Z1VANsLs9f3l0azKdXh+ib9pNEWq0VVDuNiyWQ5B84KoG
s7HQ3ljOkFvqqtRgPOnJdtWUXx0o+nxm4iNc+/rDxw0660M/EVB9Iy1w981f/QqxAMiiizjLJW92
7dZRnBsFAQ4vJimK+4NkDHOxaC3QMNkRsgN4SCZ4XDvVHBcP6EJqFDKnfYH2n/ZMbXcnYAl3aZmd
qwYAHOzISCYnAd1yk7bdrS4eczOX7ffNl3102mi7baLr5JWEE5dKHb6k8SrfdYCYWL+9Zz/VJSBK
pOwQF2aUT2LfWW09KkxpFHamoHUjWkOWMW/kiGsjMKt5/JqvMm2ytHBDrmX4Oh0u+gB6aNQM0/2R
TJIotu+tt4LT3fpIDhQVe1CDO7BwXPKS8bUNvmcpleMAGrfsvkhiNOxS5SAoosTnu3bd0D/+UzNo
T0VO7g8Ev+EZTdYyAnzcQfcd5fMtuj+wg/3WsTpKudb3/FOXhhqSCv/R3j39OgNLa33j9x/og9wL
jllA7VZAKZIU6wZlRNRCqZeHDZ91ucz4pLsdbuMOszimU8HsiQCKuUAVXhgl/V47UoJMIP9WjokW
5SDsG2X9qOmgOpEtjFrlOqF9YKzHKLXHXYVx1w2MeCGcrijv3weeBHLZ9FwjZt7eV/FTs4E3pewQ
+k5gPgRwDR/g8UWZVmATl+i+vTgOQ2wp+AMWFpZf8GWpgnavsP3ADmMSzsfCB3xgVjwBurHZEJxw
6SZiZT+aWSjfpXfaww2RP+Z++blT3fFlG41O0zknD2BPYYhXuKlgT7BGhckVggDJopmKzp1eXNjx
67ZN8ThiI2hMif0U8NqCc4xwJuNXe2varx3Dq9rgcD5+9CFScuk7h9mgrp93RSIl0mCfbH7WYodf
oJhxHU2IkTKazOvx4ArokasxwmDRTk+j8zriK4gDb6OeEd+7LkMaTo1g05ud5jKhvCfNmzZ0EBof
N67U31IJCb8fE6VKamOy6VoKK19tdaMmx8qVQzfaI7E2Vroyj+YXTYsu2aGT5sKF5ScGeL8T6PJt
iNEvyhgpiI5GsnMybPnrntyQ+PzbfKO38udxmzRnvcPkce5R17uQXtDQMrR5saKrL3skgigfqdOm
ssqGDwG1Nb5mv7m4Bw2yY/Wx5QcUdI9t6aMTtbqSkc7xM/NF1DWD58JE9s3wMt0FPgDllkj7mBb/
rReQEODCiSHnZQL4jUjeAV4353HWyPO6F+IIPMLd15lOuiU0omHu3hBWjlNTw6c4k4Z91TnIdXBa
Oxw9HHa7lpOeDbjB4BM77Uf8a9i2Selc4XdwtiZ4CfsYp0p9u05+ZRKFJQ43hHNC15qgbbwmIKiW
57+oB0ID6qh/zTcYFOXVyNCR2upDQv7cDHoOMh2j6aIb/Fpyxj/DjnSzUu2KWHkAuZH3IyS0eUPt
o8vaLblJ78zJaMIGu8p0u919tief5mcjehdpo9zuqxTI7DMRvH2WDBSRCWq7g9Xw4IuSPy4ygtcP
LIy4+zf5g1xL3Lj/D3Rj7C6LnMc9O3cxTvoT9/AiUe88evRgbK0LZSfP9QkhRiqwnT/yyrEF2Qbr
bCPWSTiHWkt2uSTRl9K1M+S5Cf9jPLcEBpbgsRzrcAHJy1LnRHBEXooTuF5xbJMtXSICnV9s1cWS
BuZnGh1+GHM+ucXeixODXl8UrWDmvAue4Zc6PYYagR4MxD9XYzxc29557GFhE/Kcj1pH/R9mpOXd
5lofqWXQbZofx5YV21qOQnXcRkwWbLJs2Q/AQs66X/zK8yxlDAfpr+sa9gpdhuzcbACyebcH6qEu
a/dtAn+crGY1U4qezPWKzgQuYUUz+oEekb+9feaVUh6EbNsAd6rY7f11rPHrC1auDvS3+Xln07Rs
dlVwB/kGowm4VM08rNH2xnqoB1og2PQ90438H0T4KoHWBN559ZEEilCTuwZat29+obV4dmFfUP8j
nnvfkQSFWItZQi4xmy5AGMA88zV2qyX/cezKbM1xhT1S2fj8S3X2NrE7GhnEAHFq/NK3SVCQR/aE
RBLaA6Hg5sxbcevPucdypKTBYTPA2IHqscWU5Sczlp2ae4VFTo0l2njVxiCFaeviD4d9Ndp6Q1en
Ym7p8JQfDUtmh9ikaKBAfkVi2IRfnNmHlCviKIC+sHgUdy1VNQ0OPaQwG0n0AKBj9tfKcrC80LeW
s8PYTyckquyT3BxhPRhEgMZufHmp8dCnp7M8dox9j+69sAUxKMUWGrzTm48nnwxuPXh6owk2p2Co
HzZLRb0ycAy3TMkLb/Z/0IAvUUZQMdV8jERju4x9IKs2B9qIRCb7vD3ZYXM4Ydl11xMzhPfKT597
yEjdTOWLofsvL8UKTj1i8w5cA7xrUAobAns0srXt/41brOMufLehyzlhJgznQKbGyRkIVes5te4z
oVkINOQT+qh5Je5AZSjksmj6+cvWQRMSXkjxVzF2BkGp8YTkV4o4y0EAHUT2ss6WpfpBQ3BZIcMA
X1bdOB0RZW0RYKtnK1Zm4Tzwb3t4uMPSquWBg/NINBfRf2US6/AfSPxtAadivPKao34rgSApbBF9
IB+mpY2zapkgBf+j3t/9DaZImRi70MpCO5Grj4ImoQ4aax8JZrTCXNoXrTItBHQzF76QYQsmKkbL
sQMijKW9SBfqgHgjjVFbxry9MHy7E1nhtER0t02ftcQQzscsAY1hcOIXdXWE7a19sJRikYBW9pa/
IV3pDrIRHn/6xI6OBwTgizN+63G0C1RYwzxPTUNYvCN5FdnamVzHN5qGmJrx8J4IpSpd3MsXOifm
ewhbPzT0DIowu4cvun5nqKtqQaG+tweYZrm/NYFQtaftsNnmmJZLYPDLR7tlNEsL9ZXl0gvKMKDq
T/UDNB0/5Rq3D/mLm7jGKKWdAfQFcVnD74AlDRfhDO5T5+kfCSeU8kYlulqwzYsVexqS4YVR9nvS
AvPR8YTwtXZbE8MMyNJP/m8zBQBxexvqM/nAMHEakXcJ8YD4bab9qu6jdnsmWJXRFruGjplmgb86
JvPK2UPnAYnlyu7sxlPFp/eZGQ0R3RRlt15fNOtBJKQH1RzKf+ZDMtOxawY94EJipvjlv/gRx8Yn
XCAmy8gL+5wZB40pmQnaDr6dwju4IJfmyBtAoI1iEdXhdGzFCfXGLxHRJIiteFq357WH4XlY1P9j
0+J43s1DCsbvMlN0wZ/GwOG0U/SA6PpycATHhwQyB0JHtJLBE6Agf4H4AnaLqiGXZQ7Nr3v5mZ0V
vWuJtYQhwMwtoFWs45YRIa67EIHWFg0tgFtxhLGuFphoB3uzKsQtddN6TmKFLrjBjuJHMhZpH3Yc
f3BtICDVwpSQ3BTNHcirhdgPSKMpHLk41R8iIVGc2kdd099r/w7w+irBUdpmzngEOPW8NGPzUJF+
WWXEiaHglR+fdDwd9PeX5NwsiwuBQ4qEdJeZraruqkMfRMMlLJqaRdKbmKHD6nqu9UebidBzlYlY
eWg1LrQE8FReA+/u1EM+jKcV0w16Lm5od65A54cIImqQ1VSNs1FR06se2LFoznOnC8dqwvCzv0vB
rO56I90cotprfpc5GZsYNd6ACXIbvMPQDEoVN6fsr1Kh2tdCW/rtwISyJdY7qlyBMS1sgIO7MbTj
G+GmtJPCV4SfgLhv+viXEFdIgNXzfo/MtF9Ia5e3M0U6cFwgrIwZXWexZ4xScqVTs9S3RWSd1DII
mNhERd9JwRFSGEaPepDS5XkK0DaMc5cOhWVR/NFG5rggsM+SR9+DkJwrUVUd1ou8PjgdW3IGgRY3
rhwRGlSz8mZbwSj1G8mb9AKJbgXz065HXW1REujLqGKiA7SlHvfOvbpkRmA+Osg/UwOO4FjGI2K5
o78Yu66VLB8DeIfKYli/DJzFPaHx/Y3ERB2FXEMj/sHnqQcPxyiiFXKEchjSuUddSAdlGZa2Jir+
Eakclo22VoThPHGTGy1kGWskrpppIq3gq369lSBc8neOm1xTSC89IFTmGGEU/F+TGlIxFEjPxsXl
UuV1ekFAAgT1X3dWguXzxiDjoHbsiy472YZdhiTmWmPfRe13TQX5zPtKCHyWwrpeiDmWaEc8m4pH
BpuNDKdlksa3T2RyFUnfc3QM+4fY2B8QzuAS1I8rZiwb0xQI+PmzWHsMPB3Vqv3nc4m+b8vk5JXS
nnK+KZbLhz8r1XSwUa2QRAPSkutbqrAYbPnHLiNTocbOiIOL55CUxxkrmoaSR+YyUQ20t8CCM03Q
GMWTs79OVjkvZnj8bQbUk+2/M3IFtWY3zig8lbI+NGSJg6kR3zTZZjYYaVc8eL8+zXl6Zpy1LhtR
Hwv6i3gMI+nXwylE6czNZRbr/vc3Ik9V19WeRsLdEeprMhFlTeQKOe5mfcBfezI0fT0BTNYAWrWk
rplhTAWDOyI7+h4/ruGZvk1jFOyADzV2R5w2L7L4iSNiOjDV+W6Q4Ii+rg0JM1U8ZJVOHifPkzRT
LzTj1t6pgIwvjQS6MCKCQeE+CHFx7dCqkskrrpzmfr1YRvNd1lws9rFYScBiKIykmxR1b/WGcr4o
iTAp+Wew0wTSxbd5BHYHHCEMABxq4J4oFGtpXRsVUit2H3zU5Wa4r1JqRwP22E3sLPqEMXJbPdow
MmNpuNqdIcgXeGYc8MPpjrUM8gUlyx/TZtF2+R4cauYVLqUQW+getNcnJfZvLmOjiUOTZ8evrwGU
uofv68IaKjFg0b/DAWCC8GK2cskJQog6U8REIX5ksUT9LftSOS/ch5qHejgN2VVfHcbnyKJE8je8
0Vb51Vh8oYCCl5WMzaVz6YdPff4b0A1X40Rxh+Q8le+qJ5/FynDsbRWWqwQhAHaY5Gzp/OKlyb8g
Z3iHEaI34/Ny1Tl6Uy6TsPKvv54XT5+hC9JPo9am+9K+7qMyHmT1nSRLtYG6Nhlr+UcQxM+rn5ip
IiQa8jFbCpRGe7OlOC7M3R2IMZamjDWJiY8jLkOfVZfCfvLDlKLz7h3t9jP/xV7J451qEp+VTtZL
oqcfFBKZ6vXVEX7r0QEroGbwljIUa3hu6n/94ye2Z85rMtB7CMR12ubCZcqm04ySGQwzPUAa6L+L
cBj71OHplLwP2I58OlcypnGqlkQzoVFJ31RY9MrQJbdB0XS1V0nGtOM4gtlM0L8PEtG8O12OTOWA
F1i2A6U27tc34eFl8Lia25Kx71A3P4CZqCSPh2+2H07zwFnwEeU3VSEg9vfEumT2/rTAo/du9H1e
WmnGuegK/pEbsUwYySbP1VGf7qnQyXp6mNqWYv1sooXANizZB5Z4SDKOtGEW9/PantZzlANipOJN
EJFkOHt5mhbQ+n/LZJhfRHKfgAFUAJTeTyvBSaXb4VFm37CnNvuzt3+gdVV6Ui13u909PmuTWOUZ
fj6ObbX3MwLssWgvxwz+lwl7/OkpF1rAToYQsW3XE7/e2yghh6YqRq3ixVNxmJZvyoaTxBzb54k4
omQgjEZeN5NNev8VO2/DWfAhFxLgJ0Qh7ieUNsfeLl4D4ozO7z6CDDh42lWBD1IL6yzWVYSa3Z0V
LY7/5ACrk4JtEU2jrSRVPTUTTDQJj1r8HigpcB36XZEFlz+4IyK6CmCZsRfJ9xCPudsYuaq1zl6J
xc2Cm8aP6pRSNgubB2kVTDAJwjgVgjH29W3KSmj9kvwVWZ5uUQiI8bxiM2CCkMjyRERsilSa/6+p
ZgMF4anQwJQMQU4gLRSpcsdZnr8qKfuq7Mp1pbD3Odo7N5vLA86OM2vD3cg1TMm2sofKiuJ4OT1u
sfcRYUabUG4wQGnMQ7vAyx7K2i04Xig7dFipw7bcwfxnaiurZP0wux8IDtrDc8Ms5tBsWuHYfppr
9Bv0Nr0QqZ8L8FVx4FjvoNcdxrVCUi06QyuuITu/V+M/VfPityWXhafr8Ve6zbnsQZ0rAG+fcak+
Hg2pjxZfH8EjowtHLoEAVjlZP2eTlKuUWATslPnJ9GuObHYuHZ0n8ZVRmecvrqT2wlyHlg1AxyoJ
HdJq448FxZ35swSNnG/yHGLDeo4UEI1cGwhVh/fbsGgMPV1AY5zyoW8xW3jT0XZCK0lYUqUclLgW
ULDQ9BgJdOLgN+JZJfSYZX/KKfKTB59ZLPcHEL20P23CFP3n8Whv8y7q1Xpn6IQjU6u1L2jTbIC/
w1UTn7ygS7quW3EZCQSoPNKYFVynQWnGgUJ/K6o7qVD3GRQKFv1bP7ODCB6340LVrrQ1hL/LXhYe
xZQQ5ORdzq6gG6lYprh7hrl/IBY1LLJ3IBo6OIcpZCeuJF/WW39uxURF3Ur/RuUZoxFpAhAPb8XX
aRvvXbpjw5/ix/dnJAdDoCtGMYU/2DKdwhvhnwiEky2VlHdqO/IKOS39KaksWYZ6pIZD42LqPdZL
nnk7D6I059waZTF/NMeHH4KbE5SLskH0sx4Z2C5vAr2e8Bj8iOwpGiXi6NKt/3p/y7KAu7Zh9ElV
9DhKNJ9YDwXowKaKdkQpxgaKl+4cBYjIa9tzRFhr8YHMF78Peos5tmEVkZ5HKZhAeDxYoZhIpWo/
6wLPWJk7h4oBvRdskDeZ63NwOQo72xUtrSMySV4zP97rZGpblh7kMsvVOO9L0A11KIphq8A/k1gp
st8gAffK9gKZ0uucKyKF5NobdDrAOC+fKq+BlPP94YoDrjPg1WyEtl1/ubXsKL6BQjYedsLGpAhX
BlBz/Ons8CJHLjTfZRRa5IguJXouktQK6SBCOznZBLBy3/iSlgL2F3Kiq+/yBD5YqjEnvY+5nd1j
+KlEoZkMBwKvV50u4pNyuFCSya3sCEOI9OoT+EMpdy+Yiak0JBibpIDimTTQR3U5APRzOZmHH7+V
hQH3jwbUPsRDU5l48Zks8gysb/84KDoE9u0TJKZiKbZo9OA00zx0s7UJgmn5sJGC+R802ogNAwlw
pD4kESZ5HK6A45XqhQKi7F4B6btdEdSsVkxl6JiFKujdwpo8kTyVJVRPZmd2j1dFeB31jfqRjMFD
v0sUssGQyqlbX0dNDyguvnLxLJPLnhiqzGfWJXFJEtRQo6nGm06M9riZjfZGCQipTuiAlai5x63P
SxWC6Qmict3SybfugbrI/R9k5mj8kDmF9al6HWrOq2nt8FYYpVjB9lwJBSeQ2TMzageX9V06Mtm2
DDajHt9l8ErZVjsIaKytqerLaas3lIyC5fiEOYOMhieVw2YmyQC2ZRvU0L+FLEG2JJwzzaQPlHHG
NQ/d+THrYA/e6bUL/HGj9/q94E4chZCilXUYZO39D105vphgkm34gv8rbLo7TsBzIUeFgdg3HDAl
8r3Y8N2azWmJg5yFHtgIkkq3aLwgcgUDmWT3mMp7BNvp8lpj16yQ+HljmQ2tgzPxFUeU/LVLxDAR
nJWmTQbC6y+MLIo6wqGoNy70BZaoYrkvPXMuzOea/AzG8NtGRPFUn/9zPsaR3bhCXaOLMLXX88ts
hgp+3aoHUcdg7Y0A3NoNxNFMukwltfKY7UOhG9ViUNo1QLlopvYKGAKMCdRqsD0o+kW9aHhrqseB
Kf7xZwB2J8ZomPDP7/N95pvF7Ouwsk6KnDCol/Zb/5A2xlRP7zFVL5xKqoxFFqeV8rWXAHfJNxlt
tt1vxcTcjVJcwHxKX39BaJF3xIeS+O78F/QNsn3lr72V8K3OEVPJgi8QhWsgd4cdXBe7QQmJuK+L
45ifxPgT1h1oZNlfMXU8SDjk8tK477JptfUo0wN3BFYua4uvox0xR2Zv79UUrph5Y/TfYvNWr0xB
/SAjzjTu2FAvai79yvUr+g/F0xOKw7sVfr6dLF5MGWJ88fA9S/8Md9PUrlNjlwZEHi0Uxq+dCiBn
yJhzfUipcL/SOh5WtTl+h/IY3QrKTUs5hQSLZ3gzDDSPaEnIiws/qR/yA9zdfILRLcSvXlJkhh6f
sPA4rLCiR9FaSqsi//3GMznKinkOpbUhPEG0aaiedJ1hPJVC1UnkJ4ctmET5I8Q0Vldom87RqdLQ
4+IvNWhxNEy1yjNCFXDSwAY0dgTzlm4UdPFszo/YHiwcevl1vqFfsoYsiob3k93/qEvEQwWsbbu0
6C6lk24Iinu10H0LGvbrpByl1kCJLOL5fW5neY1RimTfszxWYUZCrQExzQ7UVqwroWaEAACrouVG
4RcdZ3yw8be53e7Lw9Hj+mhJRBB4QMIrShNBDA7GbBEG0znu5ip9CtW6e1Z7z7x4+PkrRmfJBLzK
V0mYXtAvB4RstRQFX74gR47Rgaojnx46PCPYO2KrbhARHn/8AVO8DsOAX350RgxCHrBCbASdST4c
BpfGZI5dcgjjtHLK38Agh3vpIACy+ZK9thFuWkqIvLzeJZ1vlnba5lRwoRbV5nO/pOpY5k40PU2B
byvqma1piN0Fzj6k4uUEpOQRZSWWdsoIvrL0BBKGF+cU+eCbw/few27TCuzFWZW9ggpPZtuyRvG2
PzTiIUhNPau0N6KW72fvx81MUfbGxo/X9juAzXHpLUvykT+MrvwykfJMMuXH57kRmssXzAtioetb
LKO2HDwYs3HYESOJCLgBgzvq5DwzsS0SjbfT4fmOOtyf7iigoRJvcuUfOa9btI6+Pdq99jtxnvvy
d/3GnMwe71kwfOmGnym72JGIoOz8SDIMMplGzZl3DCaXROUx+DnWEXXfwCn+yRXywA0gtDjC1xyV
53iL+g5ugRuH7+QLmnAii+KvDym3DYZZoasj9SAoRI6R/5UpLSJ+BS97nOhjmHhWj5d6U9iikZjg
ovvgrfHpj7kbL+Nrpoz+6bTRwQQ7e3D2PjD6yJw/w4E/gNWJyYdED6I3tmCtU6gE+i8mWY2gajeV
/C2ENuyCoATQily/2eFXEgz/g4N14rSdeIzrh3qsSqZPI320VYbw9PyrYyb9mLS/K1H1lBTMxNe5
0H8ayaZkOxjEQVgrR12kl/Fu8wTohEybXV+KGDjGq6eQIXIwkOeMQ0Sjv1OvtCY83jvcRIls6jap
Qhs99GpLNc2eZYsgOeXmA4eULUjfDoBujur8IGFTbQMN3Bkdenks15c47s+nOSY0tBt4ye7cfvEg
+kK0oQSXrFtuMFk3z0IvHqEpQmQrKSSffqX+3IofVphfnL6w1oXjstSWYhY8OmXJZpi4O0CYH6br
JDAO9OLLZbyllx/7G964QVT/Tz9OGllSCga9p3Ys3JDW8RQfgoWvqowG3ZkbsBb6ADB40ElQ641z
NAjvWUd2DPXg8y4muTW3s8Fk2RAN6NkFNMXIHO8/fBGfNZJkFmi51VoxkuUz8me/7G4h0s84+PNd
yksLG/wj9dT2Ml8ukhKXV1AnMiSfxF2B06f0/IZrw2G3hGFBX6F07VbF1vIHVv+3QHrngpaWS3MC
FGPwpw7tSv1STAvmvyaIpvSaA5bluqV6dZkJSq6UBLYMoGcyoITnIhyt7/dd3HTjiszbm5Z53+4p
R+Mw1KAw0DuX18m14pN31cSa/1Cl5ZI1vpV0wjxC7MHINYJA8h9f/20XUsOgBuxBFgrij7NSJvBj
GJ0N9ddUnDAHsFpvn95PYHo/hqCI/dZq1c41j2a7yzYD/joWdH9pJEi/4FuoCaLllofPajAhkofC
ufCFKiTXGfrI+6MxjLWwyPVX0BlBcLfILsj5LPWI/CSYswrrXcWaygEv3aeueguw8wNp3RNjVtIw
+XIePBzrv5m6eemtSP7P9/FSHkxgQD2MVRvEwNSCfJwSX2vu8GScftH91FV5C/OFFj2c8I1IypSR
XMkhOlPffEUjZvstd1Pi2SD9mSFC4Grw5FURTImqIx2Y1STWaFkhYs++0/hwkwrJIAzMRtbyVovw
f+zicqLxkd+eBY60yERe2H1qpj21on1gWewN2ldXeH3hdb6YQlwawVV/ymhvtAdg3fbSUN/wHX7z
/cK+imnotZTilduHxzJhWRIv24mC+AotfOGmy1+PVRriNWjM/Fj/GG/U85m9b9CIIkuj5DldRur4
EXkT7rIDYanrC0jvwG47YyA82pwN3Tbpjz1ddgoDaG3DkrFf4ID7ISKQ1vmbbrUUXkKwBQEJlwCm
z4nFlFzT58QF+gWp26gHnwBm+1TC+MILLXVVs+UxN07/1N9zWocN9oLUP0uCyeHZKD0rOpamyuwv
o4DBogiHr4UggMiioBW6YIWzrwNGjOAaY9A46yU3gzAi/FNZBfgmnY0tEx+S8bFSFNFH48McXAlj
jOs7b7ubvYDCpUgFtqp26YYLlkNG9ixCwbEI9kpiULMg4/f3uJkHVffVVrukfte6c0rk6eQrCpws
+Qv9qVhwamQVwNrqWvpLAkMCdjzWIoS46jyVI3jjak4JBgQA87qOgZySX7/dfSND9SfZfHhTSYrb
0nCxpfLSk8U+Uta1PnY1aXMrFqq2MceztXHDfOjRVE55OxKTnexAUzQMmqmhzjYIVuoQNPrSycaZ
+Xs4qkNjU8qvZpUP1RguqexEN6M+69p6xEf3o4SNVql84nT01QLMimf6y8/bNRn9j1OvfKfnh74C
wq+cQIkzsd979DnnHdhNH2umAJk1rL39XVjxNVX69ZAOJMgz7RZRsyG1wfwfHKiiGIcCFB68ZeCj
eQun6RlyZ6lq311YY5KiRpMDdaUX9TTfinSfCsVC1dPesc05NhcUyT3KdgOPET9oAdLUivy8klOU
AhzCdJdBx495VrvMlAOgo+frQuB+YKoxclOaRWbBrjklAUmZxz7KPCLkSqoZbXAYp8Rg4KNYTjBv
7jyzT/FnA4v+vU/Ebr479IuhmiSIiSGSFYaZUMFXEakpuOBZHdIfmihTrM62obmVxL/FUMSrV/7m
4kDZlDbvtlCHRV28lVXz9liKhxTgRu8UYt1cI4Iwee5cjmY4NBAqC3u1YVHA/5atMH3GFv947Wl+
A6YJg4L25G1ZTrfbdisJfpFpCIUD9uS+r6SSPmvgebMpHhdde/5LikyNIZGP6pCv0ZUqxxrDZ25J
Vpx2LxTcmmTPcLCWDHnhn3w4rG+Ufekgk9AxDZXAoII1Ob687wq+er/tLgNjAY563FE+wzJv8317
9XfCfWm3HlCRnegTWTkAXmCKqWS2vy6k1yxU1riGlLtT8bTvHg8Pzc4OBElIDqZYFiZsQjbG0U5m
cImi4xFY2AAyrAF9UspsHzjVl5fQ8262hrGSll0XJGbCqoovmYWORywhm8nFfC3YiYh9tL5KMHsr
inyRheEeVLkamKNk1dqGtF4A1Z4MAWjK6PBIWjxGQlm/QAywhvZmW6fQG0Qggc/gnIFfdx6m5mff
7XGN3B7p269/HEUJ6KKKbzy4gcGxdqRvHW35qPisZ7mEscD7FZS0tU1NgRCmeOu12i/+BLSoJxNn
J6is8Ga4r+1PLuVEjhCGDZphjQORM309392c5+FlTwBKfsA1m43xwkAH7blNWDN86QJpr+de7vUT
dJ8/k+gRhZDMXvShGV/yb3OebP+dhXGrywO7eEr0hUbcYu4Fk5VHz7BeYnI+o9pr+PhtljjZfNJ9
liB/YlDDLG4QhYaEuFj59e8HxCDqKGXKdZYXsC7p0jvUjyWhtnh1s9sC0fBmPkxJx5NO9P2pe9Lw
ZHcRujb9Akf1T9ko8tHB1gSKiHa7jHYzSHOZX1uvwf+IGeZTkKR422wgwSjOSET/8BfWCP84Eeth
5L8EWUZ7HucuI+QcLLPzz6/7ghWyELWBg/j0L8gWGyeBzSROtEj8SaqEJQrfScwqDUo4vfuyPitc
kfsGzDiINMzoyWU3UdjE5Hd/GayXk9rrAUEcSmcfMB45pGMK3E3gNu7m5paeJwv5/G9mwhuJkn8C
PDteExgxm5PVRwgsIwdtPzmDuu9XHfW20/QTOSGG7m1JSpA34yIVWXHFUs+ErZNKrMSxfVagjlVX
oNhtR0AzkqznWDJLUrgcflTnd2Ck6j1VW50Aqjzw71CLcTAWliQdXWCSZE0rboa+zZrO65pLraiH
gN+5hBANunsO610oDulU3MUZboSVNx1aZJBraoR37Wc17kEtlvBpM+xDsRQCoIFeY+1XO34xxSEA
VmN2qZTSP7OTT4Y/nk7vbaIA57vgsXPy7iHwpaZuUTeTr2jTaoU6Hf1w8gKqOewuAWw6PrDdfjqJ
dQufs7WhX/IkiJJbZ8Uom862CrERJmG9uU0I4DMYVmJ+wokK51TAFyjc3itfsKOtJ+l9KL71PGtp
Eb6W37I6M1WQm/gpfuhsu92QsbXaK4hlZFsxBoMIDFRu7L0gYkSOSarQpe6rnUH4cLyIjkySMymr
wFjR6fHCht5OvwbfoVqsI5XimyQTeSNde1P0OdPhzpO68tX9YrkFGeuAP53WGS4pcodaVvhpp9yR
Vf8R7/4baTAjstsxBcHzbef6hjxzUUGkJ1WHag0dt0q7HNTR7ykIq/xLvwOkd4WMQZ7wKxURVt3G
ep/1ZjQPZ9AMglJAN49DFY0qFUWuAR1Hl4v2+1Dn5UL1b+HxDigV9depEuyzuABTB4m+c1APkCcN
LbQxY3mtY8RBeD3iCCAHdZWJnWl5YFT4k11LBq+xL25WfIgfoVMvh4gV/Zm3GR7jtzfPUdjlo9pd
lQfVexYebMVHGr4CqASBM+Wn8IOuzeEw2rPGd6bL8kBwxN7yuBqaf+32qJ8vyUFYl7JiyQWtIFPE
nC0xzDjeSEMHNUaL+e0y5B/56EGNcjlR74jAoHlABzOZ29Gs4J2oSr410PKJV1ANI3QO3CooIzJw
myuVjklUZfsqvKufYxABJBtD+5LZh7dp1v4nLgFpJq5U2Xue4I4o3MlF499RsOO2Xs53RdmuaRjL
lT1i5QAyXIHe5nTuBtgyMTpPlfOrX4xoeVHKMYRU7uFMJ5qRsPiIynQua197EgPyZ2FECnINFTcX
sLQr1bl14n6EQsCN5YOOa24pgGb5fRWWpVco8tRAWjRpcDsah2lvI2ZHlq3UKN7jHEyMiDhT/DY4
NH6dVeveskifsP3lXHA/U+th+zmXX2Kw9zru4+rQ85Gt73iVsBC+majtjWKO/IEm4dQGHTlra1RA
KU598tkbeb5sVyZ2prAf6He1HzDRRN3ybt1wnlEYEFWN5vbwc64u9B66Ua+U05fx7lXOf0DZcZ+Z
GkrL0LNoK6i3tkck28RLxl8PCwl9vWrkwWVPSMMwtLaw3C7P9jnP6gc2XEYd+GXM+8Y9wsnJiCQM
3V3Pmp2nkKpZKxHag4kjAR88TKF960yldXsIPsOo7JoY7lJIxmF+mTEtCAdK9XZ+aT3DbdJs0pyT
4ijiOKJfcS2UDVeDq4lPOeXZ9LszcB33n17K9ZKBdhoGt9cGI3+0EqP+m6J0hQxDrEgZin1PN2cV
2j9GoIBP5/swvbSqjhe+na+dixnc/UO75n87l6K79oethNDDOhvrBe3dgLUVaCEwrZPCTV9iBDr1
GGE3xghqfKECEIfiyISCJrsFGtrA7//OVZx4SUxM1kni486cAvN8JAtRjkB1swYlo4pv9MEn9KOs
/jOiA9itF08Eg3SLRwq8rXgz8OMhWQnKMgW+coF6lFsRWKxVDaaGWVKGRH3RiwFnOMvF5bblAGY+
4KWirM9Bq6ADCuCOloGPYLgMslbkMSh5XqgJIiujyZekocXCqYDaNxyBy4HWDcxNiCA3OK4s/MJF
Y8AATIycWPwtqKeoON+HZaYOSYcGcciwUOW3S/qSsySY5T5QGuE6yZkbjHVU8Bgswvx1ZypAx9c0
Q77zeE/NeCXgl9RPc4lDsPMITlpfD9W9ExrxnecMLhL4ZcwhD8QFVeCo/u829PCBfY2bR/eeguzN
pdH1k04muSEDm3Ihn0gbACQPqgUBLmHIG0CYWw4HIwGNxV/H+cHaLXijJVMJ7S3CQMEYxij/PbmI
Rx5UuVlHPV8Q8qFubyJxwFFCGaf1Zfr3pk6e/Upt0mZfrE7ESu5eB+EsI+6FBDPhBUE+3R2GvYaC
OxNB6EgZ1JpGHqBm7fGtvgXNgG8ETgFHeY2ENUakV33u1ubIfoM31JEhL+L0Y10VcB6WSudPBt+d
gU90wsNlDR9FZMPtnWbgBEdgmC4+IdJBFgNGpqcGL27BJ6ippCsSneBVOk5fLMOqlfoaFy9QN2lN
LFzraxKJPiPtF+qKVjbqABVgpkIA1j2oXYbq4vB1EqGRnZuSifEgBpOFyq2G+jn8HyoKALS8GMfQ
DN5OGF5vosviOEspmRRxznNp8u9DxvjAXVNM95UZZkhWif3Oz28vrx42wytuMCQj0RkzFOaPoEHD
UMoXWBdRR9NhBcB2MzFYHqbIdxPIVlOqQPYJz/k1mCRgsIcfM8z8OgkFU5Crt4i49dgejp+cA4WO
hC+uv7zZbeH802uES6k8/pIdlFVBrvEOdbHLfezzrpMwDltMDtRb6l5aVRZjSmVS7EzYA+SEAPla
aaIG+jGQsXPnANADc2IP2YGo0XPGu33igAJg1IBZ92VJoBZ9cUSuvjQFwcx+ipUoXMyulLv1mhjs
NmR+gjZkaNFYRf/QnTkZsr3LKB7l3z39/1+zfj10A6tSx7GdYNAff8Yk7eLdiwut7BktfX+ArGiI
3/ZelHX9K13fs57LltaH54dQQiZtYo7Odd4dTcID0oxQYCOsp8nfqYFAAdx4TDOQ7uBDH94CigI5
f+RFCccKCtAwcCLtAuIIa2poBg1Y+5oFAvequXNp+B+eD0r+ttf/oY93YOAX4hEkYZwfZTrP1Jwq
7IhCCynzdASvxbj6rQF3VOyogqqOlrMq/YShm0e0PhiyTWqe7mH7vR532JlBmtbDZFeAQt5MfxLG
KdDw11BQG0v1c/umCmOzqEXwVsUHNvNHm7SzAyaDUDNVitlzwyFBblOc6Pufiykf+0KA+FSgzybn
LXgMfUD0ehgiTZEuF5gTnjiIY1T7S+m/xCIyCG2NWx2SBfTKBaXsKjjfoD2dvlWYCqmvTJ8fSSFH
lKoTl4rHEpJY50jQcYrZWvRIg12RgjdCUrDvUE1fnsy65/fZA4raxLQ3VZCaAdyq+wBB1JEGzgIO
P8Pq2hp0/uYFqNAdNWHI6jQu8UK74X/nPzP5Y2Q/z5t2URZNpyCWg9VuobnspWif5Yp3TTpHQddY
+pkL5WmRiyvGSEuuU6xHzNmFSTiyuwSQjA5tRy+NQpSFRSEl4ASY42fDHI5q/nxLlgDU1QUmLymS
isdXzUXpmIgVQaKhxJFus9XeXqF4odAUVZrPGUtddzsGL1Ate4r93rBWDylbcP/qSZm0jA5xOHf4
2ioerk/O3XtPpH7hGD4AbM+wF2Q41V2uK7bBQpviFSjIrEPOy9B/FYPM3A8DE3TNzI8hJ9OtwYtg
AdZuxK7d2oruA7uqY3TIFDjOiTYZJSASZLInHTOizXFFyetndmLfe++jIttKBK5KJsaZuhMUUt1T
6IpqddaTbdv3/lVq9glHAFyKfQv4Nt1irMZZpa0FMHHZegEVjJScN6A6rLJHPgT3FErplIpRc/6U
eNae5Ain0kY322GaFdzK/siAbv55p9iDpj0AaNaAB/5GPVB9CZF1k5Oe0ySvBJicG83nLlCO1UDc
fG1P1ceeNaePwY3p+8O5JXPB09aIL3b8YI6Fu1fxirsztCK8PMOgX2aMGpsiX361jr1CUtcRx+Vp
z6ceOwuSIz4ea2/BhzAl04AGU75VYZv8umr48CY8MhWHMloCGeD7N9qMPbOI8waXw7I0eJcWofI5
f2/CpCy+u4qC2UynRcud0cXg22BglUfdi9avnpZcA/qRt9Zqmg0CtDJXF+iQp3yH+qZg3uMOZeyi
O0htSxIxiAO2dpNCHjTukjyni/tOTBySMgoKJIRrnAx/TcKzLZQJstAy0NpnQ7ysnM7734Tdu7R7
2FJySGvOmkt322uIK7p4pTojT0smfNdJG+cvfpD7Gp0yypxnxNcvYGxmXA/7+i5Q8FyHY6AzQIcp
7VctAdNufLAhT4GiWHi/1meigiT18X/rMQYWtbpFojwIclGH75MDIs//sKv7nCvQyfnF6tnH+X2c
I4SvwIDwTVPNdpaOeqHzw43Amd4YamDF3sAvwRyQRcEz5IT6Ds9cH5oW5VFGP/EfbekYA9XESHKL
AkejWUhD20Q3WkcKlFQgA7P2EMCNBKnbISPCFo2Ot1mIo8caESy1MjgzmmLmTQuuWEXPyOOY2/uq
M0wfmlwFvkrRKKVr9c9ynz3O4fL37Yt4Rc+1MXaQMMOQPqNoozvt4Fvlb3Q9GgkyNRs8qQqE5T/7
Wmho3O/jO7g5UAE7CeoPGi7H5uCYqbVK31Uuq/NGmZSlrPICBwR/EW0NvBE+F4P0zJ4nxfWrBZF6
tlv4yCX9aPrg+/bc/Jh6ehGEnyzMWedILTlXdbTLGLc7HlPgf78DV02bbpxqYuOK7VOI/yD3Z6Ut
t6tpZv61E1eqDZ9ftBj0pd834vYKwEr5JuN9f8T6hxowZZN7JCutjoLZLL9zJWniNO8DJC7z3uBQ
LznMmcHoPbeMkmvQP+fec+OyWef+qNylB5wZI9bWESwx2/5iaMqoLgRWPDNf/yWWBlM0hu22/wCK
nbVa0L9zBRRvzelCgjqswmvOan3jlcIU8ZoQ27R+f7DxrLx3muwXQ7DDPU45vWWixl/ZctI0eU5R
Iu/ISTJ3He3TfpOgiwjGVsCosCv8VDuwn9sg8rk0t4/b1nsRYeW+EwcmGaZcJJYQDZxMmXSWRkfS
QE7vO95z/JlgmCMv9ltI52hV8DEnMW/gBm2U0v5AMiMZRb2+dg4tRerlTtG1KVtX6RmakQMVsDom
gG4XT4q0aIpgGRuce80ADXEd5DNOlpECKoBhCKKzbBvZIxvs5BnZ1a2gZpjUozWAVcre2DcVun6t
H52JmzhLu/M2KMlOqF9KNAhskMpJgRkbekSLrxw8W6s/vFQnW/GAYHTKZlnQQR2wwql2dSy2W0O+
DkSj77n2W4cbZOBbiPHgum/cPhMsyTg4Dz0mN2wMwt4Zow+pV1nDbNexQvHDySFQbQPuYd48P2wO
NmrDbemj0wm5Ea85tMPx8+7hOUsHJ/84tkRg1mirV3PHYHNWN+357KLQqvlG25yuq3UK+i1Oc7ip
ovjWeDonQpAV0JtcEBrNZgSoH3SJJXi3C7WzBNY2IyVbX6IPVVunTTIzjw0y1MLAXAS7p1zB4dPE
i4+SNHMuGjg7ABp6s2AU1RmFs7TEKw1DE6tRz+zyYvvnlV+hgrBk4oCFIwnpsObsfgyPjFsV2SEM
F6BRFn4po76ffwjD3ij7hi9MMqMU1+uBofjmv/6b9KNbMIxaM32orK0KAKxXFvZ3C2KQnrJaQ/jU
bqGETXFHHKmF7/dyboINYJqtz4tTPcPWDQTlDDzXKLi0XENqhuWYRJMRNr5R5BD7gXb2eEada1Nq
gRmpBcPMQr9lsCELLD4oeu37ZveszEr87otglzaaEP39DKNCPrKnpTJHe8ufBPTr2jKnQ1JCCqTN
8ujoHO8Z9y/trMrzkOZdWYZqDGu52aIS5z4R0/dpD6Wj+3k846EVjHx+xR7rC5idW/xRtu8eHjmV
5kgDylVKYThLmmB3bvXp+rb8T0S5eYjprwP5tbL+SO5Emunu8b/NUsEpsklQoTQ8fNuiM5k0oQfA
9RNCL14XSE4u9oxhz/eP1xdBMXv1sjtY+H1ANudkxm1YcTdM4YUaaMbl+6x89y/E80vtAZAXKb27
POw8UFQwJB0lQ91IbW6JCuNedNB0lfV/Gzex2iunEvz8fKsj/Au7LhWVlvjVqa4JXgL7uWhOy6GC
iqB7cLF7RTNGPW15ZZ0ThJxnCzHUeju+0Ecxd3SbNHOH9zxB1GDW6IJlTfXXuMjECaoCMlFOc5TX
3oyYraiIlKDqv6UKz94us8YUzXHlyn2LCUgRyNiTl+Gv4yvH+YqJB2yTNhH13wL+5ZZNTtABSKqQ
+eE3H5uel87a8F10nAP1TzmBcLCEccob4nIPqF+tPnrfo71ksT1KvbJcxSPRqrB7qdG1uYaW5xYe
0aF10BcQ6PSvmKtzMVr2CpxaESuZmBdS4xkLbEV/D5I458FWsOGS1krrZ3Q8/zcHL0Qy2qlHuyS0
ezox4/dyjMV/34R2S7/ey2lvExOhbUwL5bj0Cz5J0qyzbT1alN9E0uS/O4gYKd4MvVVZWxiEHjYa
nxs+UBRh22buzZkhyeZui7ine46J4GTZdDnuwmHPPJMjDVfl5Jb0rBurPqgj6+qKKUDEFurSC850
pzkVnfDG4vAAjeM/BlgGc83fEkHW1UNkPOnDs18c1bxWNrbkctUBrIIi2YwCuSuyfCG2OKw41Vg2
nn6x2dYkL47oEULm0Nrg9wTDGF6LX+0NcUXIHbE7l4NZoDcfBqpj9om3Kg2ltlxCVS+T33gJfTAp
4/YoepVWE7O2lYrt7ch6v7Nfm+QMdNrnE3q8v6Mnp3SPc71oYbjpHc+oCIAHvz+ajNjp0CrBMNOt
I9HsaAxrDQ6NB5tp3ql9B7PBCgH70u+mRofHDfrz4lMp9mjvWvf8TQ4TGSkX0bnpPpcRg/bpvmai
6ZNtMMmOBlNqr0jO0X1X3eth3C0ASgKqbl6+I8DqSR82NAviFGLrsthgvJjI1a4Wv773R6YIjX5c
mteoB+mrj/FS6B5Czim1QSq2SzPtaPsrAkQ/ToOvEbzymu0xzcYzEnFciezKy5uIf1S2xqqx3hh+
Qn0GhTpUfOJ+WJlclmOBfowxRj4lfLqm7V7VCmmyJ+RlMyw2a5KkNDkGXHpo4+fnqfqrzziXiwFt
9Zlqa1rZ1qr/QQfitE1SM8kvK/ywykV+BanEigDb8TlS8nB9xyTe2qC4N75tK0gI7/x+m5X2PxHA
Bcgo2gqfrHNpWh2ii5fJrZqFfHYXI/rv0Luna2ozgbjnj/cjxMxm8BVEBD3fDPyMJLQQIdDMwtP5
T5qPKYigvu6xuOFJZYS/7Cbyk2JH1fi+aB0AK3bgK8GaHX4USV0d2nqkCcLZNKKNm/h+ClcjNyvj
y8+5yu5eIQWj3k3p9A+53rXKayk33MJuAJVajzBkNTQ+l41LqTf7qC78l7TNKZEaGa8UtaQMtMwr
q8/KLqvJTer32A1aOZZFiwfBBGIOet+2z8GYIZNM8TKyLLtmYvEV2qdPlB/svGofS8pBdbO6Mu+T
mGWDVkaOW9Ds0yuSKyvewSm32tbgisIc+fQWiFk/Ndp+3ib6uaLe6NnYlfBvgQ1IrqlzGTCxf0jp
CZLoDEvQRszr/E/N3KUQ+k/3/TMc41dym/SLrjnzuDixDVyHjXc9MJUeJTYiNY1yMYcnn2GTEz7B
LPfPBwtxGro3ASP11wtnh1iVj2wPhK4IyRwcAueHRCE2jprTPPHFdEoP/iIo2FlU1tv9M/f8BwjH
p5hF4X2fHXbh+O/vt2qmSS1huyGKDeny8hpoHIAzor6mCmn7SrhFSidjGtm3Q+zucW2deheiwmab
yqlDGtArSJpOJjYSghQd8hv/UJJVs1G7XHPPYPvuGTVoNuwPLunfuOOzC82KBez5jDWojzKYuEjE
nP6N6AFy74WvAxUAmzra0jN6UmtBLy6iikR/3MQJNVr3xBwm+dtvO/WzQOZp/TBACtAsS+Rcsjpg
bZ+CDplXAbUQGroOwQZ9w9PrWFgiFeQzuJNL1miPfrCLKEKkGUu+glosJpvyqRiBx1tIW0FpGZ5K
MGNwr+TyvsYTiZKFOUl1UhVoIuOGebWWcOK4G2z49qy6o6sIy0CGjvub4TwqbsYYKQhJuqqgXQfo
hdXg5Bu24oy7zuXEGpCmcZoc973KgXAjpdmOZVDwqigYnXjKdTvGwoWuTJK10X9d1A8D07FesBpP
pdsS4fPSteoIisJQU53OBnaVuYNISaphTT2GS50t7dGJ1PmGKGgZgnEP8JZxkapYwYa7zZC1wFRD
I/fbj7Jn/u0EwPG1kAeKRVJd2JiUqmbxlrLo6+XpYwN3Nknn5cMhLlgtRc7OMsV5yP5iAcfh0uE5
AMKyuSMVC2HmdreLlSMeEQC0ZMLpRQNzcWDNdl9C6imuRPEL/VZMCgAGqORr3xiMerQWHQ7t55fU
MjPyN5WknauM9mV4ZSd0Fwjhypkzkk813jK7WfC0283srcGKpS8mNYeaBkcXwbcQIS80sOMEvcAO
avZYHse1ohOeQdUpW2w2uQn3pJh/EFEi7lE5DOTBMgX1ZQH3S1vvX3NeKZ6jWVkX1rxUW6aJW8h/
NJIcGBMrSwwDIg2toTC+XEQpUXDbYqJBaeYzVmh6TIfy15HPOmov9DD5/PU2PuKkRuXIqAhW0Yf/
1nirHyYo17xprsMnPveekLiv8Xp9E+aRZPiHHAJWrxf1aSfCaCfExejNFPkpmqqk06uAy1N4fODs
9czlLaizPXp+2Uv8F0aOU8KkvtOC3IzzIIPScaz3++O8ljAyvwNS7YPvw5qkJRKLDUb+xb7M37KR
/xkeTeJO8Q3MKehWLYAuEgwA3QzXW/CoBcEM+vxDlk4GjFdWuAhhf0NrUooG1CMyR2c9lX+bhvIo
RxEaoj/lxBWg8RSTG8yFzffkYQBzmYBGoQxlzlofjmNWuWeuDKK3clwIJ7o8KbBgel5klZzuEiTz
rEqJQNcGNciSZ7RvAZ/j37z8wwWaX5VfqGvrN8rPVB8rPKD0qc5OwL90NQ8mkkUAqu6il8l05bwe
bwqV+AyyrbiYjTDetaR7B4TUReeZWqi+orTMlA1PL2QxxQG8PfcHdo5hCVt7uA1T1gClxJix1BIr
ILAiUP9IvfrnyL0+sfdAJRnzmItwHmt61kQ3m6WUppTHNsfCZoxh53bb4emQZJqJdBk+tzzrJG3J
zHkZigP4c9jTOKmSxJsmoxzDjCG4+lJkMKzGp8FMm1nxau9KeCL5dANOgUS6ORL8KkUHgQ1j/xZ4
7R0qbMKoyPNvKYwAXnQzT2Iplhgm9GDWZHeIJp+9Ch0yCswijt7nxV799w50QWyDKSSZF+Rl3LvE
cg7NnhdjyqzG8WcekMz95ZjOELAg5rDQI8/qOn2f66Ef4j6DO56YkLmGNkJLYqo7/CIQm+xa1dHo
Cf/mknqzj6ld8+5VVrCYTX7/bOLGLSw3GG6RW1YOZx4aoId17VSsLMXgFLIGHGYTSHx/IY0/D3m1
wXLx8H9Gq56Yc9kfKIVGwFRsBD9YuHA/TrG7RYAvipR+MFrKmeoFFaIMoloAN+eCTlKSblIbHR6o
dyVo1ruWeJbnzhTCtl8jQEu7+EI1/5o0ATsvekcO9HOgDaoe2tzDCD+wLzYN08So81B5YMnjYtuj
2qIcRj0FxZSOWBPajfQaNA8yIUWx9zib0T7k6rYqmiyEttrV5yWHFkVk23B6mI2L2B7ndGwYeMnP
xFXrVwrXexX2PnW2LA7sa0PxVj01dq2OmoGN7RWO5+PoT21S9O6VivU4EHt3n1bpusiWcDmIWX9i
qDbLm6IZvsD2Y9raaCFn+O0zMc+I+W/rzmJmaRCzZovrv2HmHs3eEd+jRkMRBLKnRUk16NTSUVhf
7IeNzggJVqeF3YkLmPo5K1Snhfz3K+lJ9iH6mWaUP/rHkT7emiiSgp2Z3O6ETHBCZUHiYEUG2Mv/
1QjCY6tEMmNHIWAHzWGFNdsHoSOd8r+bZIx1amRjp7I8Hd3cvJLycD//nYVK65P8jXSJ/b8e6id/
5a/FWdjbEPfe2ewvYBV1xvuxN1d3NwwjJmnEzgQg3AkW3tl5bRe3NyIZ0W2Qw36IB905iBrAAm7L
Jk7ecg6YrDFkVim3qJzQ+4BDRQ8WXm9PwgiZ9LSRICcFN/CH0sEfh1G1C5tTWlGDJysebe0Ep6uh
3CIFrY5VV/YGs2fYwlO1Ec0EQrhrOdmaKwnixWmzjK5FysOUAJHOQB2hb09JUg+JU7tCg8zYt8k6
rR0bUEcqIh056fkzttFtd0OC9gjh/NNFEl56LFuQ8Mj5GrxH+9Sw+EW4gztS/6e17K/u7Vw9tCCU
vMvUamSTuRMMQZ/fVlniNkmVyTc/ReP2fh3e7DDfRoLAzYU6slK43E0i2Xzw9OVF+Xt098WHS+nl
ALRBjVCuI4X+S6F1DfCJUCwvZ0PXsVdFT4RJuxGSrhcDOjJBce5Z7vVr75KOOKD7cfHXpRDDYzc/
aRAZp0WeEHPnZEuCuTISsimtAyTNxYWs6kCggiFUDXjx0FzakfRgmaNBfwaxUtiIO6N8lNd+pZGw
QCN01K5fx4teqpVe3fuvrjW7WB+KAqXAGec2AJC/cNvaOBl1USeVXd7zMSPzNXigE+J7EvsZXhsU
0POSpnbwQw4ePj902X4vd9EBnMXh3zWWgGw569Je7vDIBl26iTqv4KC9EV/0aAXpwjBWgj0K+pDe
TFO/+fe38+PUJ7f1/aPuqFA9m6S1OGgU1BdhtP62uNzTRFFZJXgp0kbHxhLmdL95KbNZb+MQc05u
4aJkATmHl9HT6ZWJeRlrqEE1Hlu+G+rnZ9Du/XHD5DeiBS9gbwfV6WLzK1Xhac4DaW9fySluziFX
5g1c+OPVMtvh//SS8q3TL/2qogUb17jdBzm/BbR5r9Kineg8zX4nVDD1zSuGuAoy/5fe1FQA/e0v
wl57Arfngq4rwvAG1CEXdL6rdc2WTk7qFl6jSvQYKQwzbLqay1lvDNRSIHI2c7UyYisg2ZC/qbVN
9lVT5cCMvgatlye0yBF6lDrYbAH2Y00DddKB+X27Mx23/sNIAePPMXNIePzJ5/JeBqQ5qZgHGRPR
F7mIKNz99zCCyYNbUxb8tgCzux35XyHyEW63mEhjoc29IHcAx1Ox41D83WL1qzS0WY2QT0Huh1ez
WNLPq5qKgzXScX/PfOQYKSig5pvZUtbAp3+FPOFS1xkJ47eZgNE4A3skA9YHO4ETGWz9rQLfKB/N
Pz8YDVxTmE13eYQceAYbNlUZSrlALSsazR1SDgsUVP+iAAbEHhIU7LjsWwhbWWqWWicMfW/GXG2i
Vz86Yc25t0/rkOYokc6zooLK2/qHvBt0fEynVQuK2kTzh9s2cFeLigZwEDTxDB2rHDIjV095o6Nq
hpCV081v2kTXEOqUmBL+peTaN2+8TSbxaNOY97F520kTgFlRf8Y6E17x9BEMe/7gBKjAH/aCdp5J
l8d3TUV3u54iDcky2UxbZ476iZR9Z0/o15DWgKPKkDdYPDTjQuBCpUxjIuoNrcmOtD9sQwt+7FRC
JgL4Bqfey7ZIZ4WQQ9o91/5Cw6F5qR+4z20ZM7g1EaZ0QqUzkRiUD0bhVowiXI+UA+FDRieloGx1
9rMmy5AODQXj6kZdnOPv5hNPNYm2Iyb/iPHvLSc4Puf+1MW0cQCeCbZUhbopb50DexlEIDad2DEY
+gosAQ3W8f35O7jbFEkzPd/M5LCXgmKzYi6VYe8fZp7cJhondo5N13gvum/q25gHZmcWUPH8VNFg
88HpA0HP6FR7NXsCUAlchVbwtnmaCwp625YRYojuqj9vNsau8uNqmZpfzSjuY9m6N0ibEAYypYYM
VAhgdmw5KMd+UPuRf4bl09L3nHx9URL9+0lWQEG+p9j3cXijr4le6MdMCCLMIL+VDsFlJ4CzX/Gj
xYMKYPqXB0XV3UB1zvprCzt6318ZV8AbqZ0q9e3hdRlwUtxUkJacc2ZTE6A/vnQGXievfHRfyAkc
CA4CPxY+mzjXva8JrZ85dUsbaA2HgoeuEi8/ge5a/j65eWGqUatkIFh6jeky6sCGsXeVNiKOvX2K
eKOkZarnyF/9KSGqLVcnBVm1jcFBZpbhyeoAFcTry6YIGgo18kbfo0n53E7NtTQAMeh9hkp9KyGu
yf+f0P3aP0CuA05oJaIape5XvqARhVY7kYVihACLkzgL5uxwovGThQmTVrATGM9+cGHiqG7YKnUh
rA4qn/+o/UjgCPS/Vce6TXBiaz2JtrySA4C8DfJPZedFEtQXY9TW1GQDsofIHAzLrhOENMzFG3uk
s3/aRlrIW2vZ7cqP6VSEKTeuUZ7nq/krejeITkSlFCWdxoIYf3ykgY3oA3atELBV46I2NbdL0jS2
+njq1YbzdZGxbQjHoa8qaEma8Tra+ZdIEiGF/AAFNdGBJX7f+PdkzmejeqPeZ6RKxPwLJw1tXM5R
1wKkl7tRCG73f2/E0x0j/ENxQD7OLBRt6BpKOJjeNnnNxj+D5H37XBwUB6MzU9QZ4fIK/wxFNRyg
5qWoTHUCM/0lZIKF92SFdQiGpy3JiVNY9Z3R4DJFUmKoq0e00GZ95hrHOieJNy+Y78beopcLQsUC
1jDlamsRxdyGV9Jjj9C2MxNaY5TE6lCTlRuZmbTf3r8swQcQox+KARCFLGV4ZcjBobh/ZoaZ5usD
BDWrzswaESfxOa95iJGbu7uYBQHu2ax7tOjb6AXGecowfEn8PQV0rsPGAkax7rh30h9E6JVqRgkQ
JWU39KA4aMjjbYw79FMxW06OUkfJeJX5ZPZ3k/5graEQtaE1Fj3sbKcLEBIN27fTUs0Ff5Zagl14
Yp9fT21V3wCWjb/jNeXIKJQZhpUCCYgQbeot7TIOvvei/XwS5HXqCGNVFL14JuD+E3qQZ5Zi4bYu
APZsqJO89fAbQfaBjMu+32CjeStfVYCJv80zljNNdZSyBXMgCPfcT2PJSZBHxWiwcdwofl3wuDA+
SaUn3wDThje90u3UF4pwPyn4NOu1XUYuAJwtmpxXCtrYcquBT3ZrSsE9h6a7HmLBuP1awyuD8sgI
RnILA+tg6mGETJpDBPa8r8CIW79i34bw8O9wGVIPD4ycSAaNCaBNlYxSMY7JBDqne2P6H5kD4Ov8
+5SGp46nXTYcCVMOReO6TteMX821y1fXDLi0sH6iwKr9UlooBgEYwRCj2fEqaoO8oahHg1HRy9Z/
s9K7+wZM3wLhBtd7tLXdgYcRe8gR2BWvvpdIKnXPWwrO7YMD1Qz8K9FpkEiJaPI71QxBrlSDzkfq
+5VGid6FE+BOKUk0qeG6vBGNmALznMOGNTS+wgkVKEzpiENH8x5jvvkrMF/BmPCkxl++tMQ7ibFn
temClWOyiH7M39TY9UvFhEflhsO6LTO4+ZUaRAsFxIZsCO2LZBPNv/6LRC9CFp9G8bf5c9PE70wX
98ZWtnk00lTSDA/rGOr8Sv8ZC+//4pg148TiiOh/nrTTiuyVJdTfH5rYBHHKHKdkcEiufOOG4gyX
R50UXG41loq9/YwWGRlAdGaxDVR+WTP5jZJxfaqWWM1PcTyRgnQBtQ/1uoxmWe/ZvEn4Gi/zy7xz
zVDx5hwX5v9/muj7IWpWvRPRC5lgdOCMRJP87EqDMZ3Wq2Gp2jM3uuPEdkTT4NSOWNUYeSi6+oI5
i+a8tWoNnFEqNsdnm5Lymbsf+MRbZ26Uowb5V4xln0PTyYrqCp6nAh02AXDoNo1Ug/cyliLnbQs0
0B61ANat56U9yt2OEtTM4xTtWRnPYpgwFTidaAnmcc9hy5RJCtY3+JzH4C4nYGFURe7WXh8uuU93
hgz/Xr8PjYgmpwl43bJ7NE75QdL6pP8lKc+13HWiH/752SB1ktPOVQK1HPPTEVzW8A4Xd9k2w0Bu
HAWdFaD3uZGECXqXsHpiyw2FUXDdPi7qkjzKhKkEpssgwzI2ZXrpqXPqivlajg1SXrqgVuiuH/PZ
GG3Nuvj2J7Mf7H8R6Jo11YFU+B7XAPuIB/z4w/KHcxVYQrrvoTbL71tdPG1L2pomLQ8iAvu97ENO
ZMUiga9a4+OJy33U79IY4AL4TmdOotttkd54Pm6+f/M9NAw092LDtaIK/hfz6xX8evG4XmrBFI33
xNh6/cf/m49fIrdXir13N96gPHjaeQhJ0sbFOAp2Vc4wG5Sj2dYcFgYxZHxfKFLboWP2NUrsK754
gGnerMs9uCdNOKuqVi8VNXLod0nqL+PrE6eFUdaz3nUV2Z2HRPYi/JHqmWOb9kp+g7PsEF7GSV0B
hPLuZbKRFTibhrs31MM2GGPVIcS2YELuEc4vIKySkmq3gRCHTJDMeCHmdpoeG7l8HriGPaH6K64f
tIsI1ScLe7O8wnyoj9ilUD5tt3CdUR55pWxKxHBn0DytPsN4LE15J4pmw8HsY5DnXgqhjy5Kk7z0
Am3JyjlbnQaT16SoHJKGfQO2hPrD+4Z5bZjy4h9Kw7apqillj5Z1ZXjkPgVLEPCbJRDEVcwViI6Q
PgOQkNRntW9UKV8W9/UdTTBGoMtUbHJDrZnaRK7+vuec3F9AP6/xV6wIDr8CCZv9eOgsvt3TStRs
Ckr0klOqU+SgCiRrR/xB+NUsGjc9lDX1BzZB07R3Rlwz7evcJnhXMP3eejZjtJn3ST6ZilfvYXzC
fwuGKsZa111A2o8DTMMN57/0h1D7lGfVU+bNBZh90wWRKo5Nnt8xYfPOvIMoxRY9/gysvgbq1T8o
hQpmC4yHC7+9Ijr+TiQ0zHde+TdBbGtsNKVA3qdpj0IkoIv2nbffaBoFTamnoAZ7IfVOc24xiTy6
RCVFipXfHIopy7IdLx5hEwbYi2xiaD4FJQJ25PZ4Kv30z2NXEZ7m8GJ4Nn/Rkm3yzezfTntO4RPa
k9uo2b70HGt9swv2zh5cexwFVHrtLYnq+fIIyepaFw/k2XyhQFM6Mq2bcpAdVM9sqjBO45uPQTcp
QbbM3WZXcJt8Mqx7tm6Oq/LsJEOgQeNnjchW0fuvTOtKtQCMPaYbX9Ibj5Vtrzg0YZjwAZAd4ER6
a8/86rfg1BBP1LCW8Qd2iEmzDuq0EYLQOXGlpK1WxOI/OfCOKbdAT6fHivHp1FZ4Q9unGd3nSkpH
C5bXJZlBKmvy7Ht46XxK9sstZAC1yAtM9lNsd3J1DXatMENvzF+9YQs57BdzqxctNp7+L2LCpHS0
x50ClvvglK4HVIHhB5wBaWIMjO8xEEhJYFAZs4DiPMzmuW/RgTTWtzAQ4z5fCXMEOUUNMdYy/xN3
3GNZwN2rz5mIjx1C1SMsl/zniUDWXBTO0kDQMsCao5lFj6jk4EmcK7mzszYhRIHUT5y5uUHh4yjO
JMVUoc3Y7Otw4UU/13dn6t+EZpWR0u2LAQnVGPvMyVWg5BYu/C/xD49JCJdnEY2aqz7BYtKcIEwy
TuSaiaWB7OoV6ghFmFh4f4KL2SpVqB+P/unrNeosJ4gLQAhDvMdpGxg1p04g1tTBSbzfvLUTKb3c
riZ+BceRZnr/J+6nfDwP5WeZKeBxK+L+m8QSMqOdSXXl0NFZ5KQZ0qXdwd07y0YHe7xpKH5dZOy5
X3ZAXTrw83dY0C30adbDB2s5MQkByyhgK0oikWIU3oxoJWicurYCGo3rU1iKd1ZyQqA6LhFpZ2Vt
hlRFusMJPVP/5rX3VPKyJoTdT9FDAP0VSBNUQLbc7Wf92xp7Anj6EkK/z5HdUtLHYg9y9twPhbxS
PzdXJkXyEFUG4qzod4n0u76eecZPPfFuk2H54aZap+7upiTaJXctjayD8CUixYy3snnyspMl1+kZ
KfOcOoQO7ODBzKrbCJ5jDZUbT1vCj560OAYXhBD8+/QtLrQVOJHYJG5OlvIz5HDs63GkpECM7Q6U
kqriB9lfFfgEmawqC04j4NpMB6BDP4YaG7myjyOlStrrH9MKNU6oOTkyaKRHIDZlNh/Y4uUSad6n
jvOMEiyK9B0+S3q78SJ/qwYAOKQu1gxHN61pos4MGCpw2mUIG63+yDhOrf4kS8E1Vcxv855If+bo
ara757sPJ94REWwg6eWejVdeumVscQaiwJkEV0gLh/ypamiYqGYn1BcG+9fQ7bFKD4l6E38FZfmK
hYbVdxDQKC/XnSiUMPfpjHDd2Tvgu6CwyywCK35AMHHC9KO+I88nYWGitrTsjVDjhFPIqaUFCm2b
9i7Urdo4svbYXZdnwjj0WsMME9MWxrTZXKpKTZrUi4e45ToxfGMprkW7ycOglCRu0vc4QPRVdQHc
g3n4UhNupFEE5+4nT/bgE36RUDCy4Al+srje6OY6yHerwJyWEg3XwU603Fh+Gm/opn7dAqc8Pc3w
zTjiH5SGI3gsAcEaVpbfPQdNir58peJ/3DKXuHFCrI8GQhukhAjmeis5TWijA0MCg7EaqZcWnnmZ
1Ea7r8xa2YTDzyBtxlBfaGLT0qrzUO1eUDaDOXvJJ6HBAY7E8+qlHuJI1EfCW9CBZtfTByGR3lRp
EOc+ljI1LkAHStQ6QSCbdKrp4TNXB7bVHnl1cZf5eBMF/6ubmz7hWp9oulQIvXYcE4piSwRNIXgF
wlVaFZRHIKyUJURwlz9f50E98dc3X/Y4mHq7jXxc0ypz3nJ/1+DPLlkQFeK7LSi/uoQVGLbSlXv7
eDJsg/cN6YwLw01snHCGEPIncNApZfG+Y1VvbcUwSY+xElcQV6LyZwaqTvJ9ZbdvPjAfTfBbVA3u
58wvg+BqYcuAJJl4Gz2GU8FmPEmCfFmTOI0T/HN0OjMZDtYeopTTEP+ZX6dB7KviGet50y7PnWkB
N67CaDyaDs1WGf7Cy0CgpjaxI7Fw3vRRWVSRagXc4pCT1lxxq01H078rMg/t4GRL8Q8k9+q/ISai
817+OJDy4JJA0rjg8DXB/nLwm2YcbRCs2iQsyZZ5M0x64Z34TcqPB0goS7dau6+kXkmZ/Ed6Qwh0
aehFzJWVzna4E20c1Zk62VPFdL8KsmlhRLYknhi6Rk0GmioEZaw51gqMoDjSccSoOGqm7vYG8DVl
fkFVN4d4JAxUS3+xugsoe1jMxS1gfnYlEFp59Ek33oSfEMgJ5hvPrwgUJq9a8CyDNobIT3PE8MYb
YUKhC+DPi/t8un5ke2Ds1qWdQE0dL/fFws8aDh7QswuWOB/MW/3KUb3uQJUKnsxe9LPnlmIMDkVP
Mu1Csdm+X6Yo2HNtRUAsjs4HybAaNuKUrAimj+njFGBU0RmWqjyRRO2o9H7X9WiZICE2as/XbQ/6
GTLjxM6xvU0GmsWhNPc00fcGwyh+FzqoMs4kA99MglYuVdiZo8QnnRKXSwiySFSRs+hb7d/QqLam
QjWzt6vR1BzKHjuJS50kJ2uuhOadHVgyEsgVHLFnH21OQgH1QBwki00uTZEuavi6bxBOTjXELxvl
B8NditlhLH+eSK7DAhZXZXfmBl9IEVcZHO2stYq32Ft3lR1yMSI4s5YWUdqhMFgUDsZJ9xNKsej2
suuWH9btvpNk+fA/aTRd/e7HiRhWFjabnU+4YFag/3Bdpg4ZXcPhEdOIiOeetkuwSgbHsyRDRPjN
+xuLyQTTX2s/5QHrJJsEECqBkwrGovCmDbw3o4z9tF+j8mElBwI1EmAv8PyBRjzeMbRcatra8eX5
2IcVKNmUKbPdPMmeqXUmFl8mZvknRMk1YNlWIj0zBKkLCs6NbJ3tnyj5ktgdmbyK55tIhpslGPuK
sX3tIkmw1XDx0JxA5s2delNRj/tJuEwSYueeYJPI/BTzEGxLosGuPR+hhbvbl5sV9JqgAkmTW0xg
BaSZ5JtQ1lXIGymJqOWAEiYZ4SftwgLH3ZKV9DCcesN7gomxN1NEoCMJhDgJbl0l7Th0wFmWFq5P
CJBieQ/V58Asoe198UIoNkZ6qRgVU96cHK/lT5GT4udLHbWXtyeF8SAMnWCUw+eqx9PjZAPEZHvU
moUpwyGOA4l9NlOit070nwhD/GhpLEhzWUTsmz9ONAw6pA96InXsiEgCrLuR5M3tq4JkCH/OYvjp
q5hdMTHj/yj3Ipd++tiJsp7FHwJYdgI/jdqoILNP2LbAh1+68Uzp5SZmMLW59ynPneq1MXRAoTU/
nrYwKta13jyomODPR4OH8sfhVBhJ7GQ4qL64zbiWNcvsv63m5NBI7CGmK0fi19jAfGQaGGQ39Cat
8hjuwXgXKhzzYnr6+OCdtyEYjLFKnneByXmYasrJDK94s2cDk6MmEuqy5BQjvmDs69vDfowgjKvV
WmP1Dm+NzkYuZHcHmjdT/dLlAA8VNFHd+uqdnEJenx3dVL7z6dlMcFI6VxLmfG5i3FyUrJ4Cm5nM
taNfm9pH5fP82/3TIJvrDORJ6YNf5Ita46v2m05DIdblhB5Agcjj5BYHkyYEJxSYZPsm57byxwIi
2rKR0kCntUdafU2A2WVfaom5VecdcaD5fQIFns2vkgvAzr5eLeO3k00vrtBVTD0aife9LVq5ZbEA
6g5k7wvdp4ExrNQnIlDucJBapYfW90MNlFsCLTnm1vSHFS8UFpwXLH+tDfbxyzCVyFgqfoHzL/uM
z5Zep9WON/F8pvrqMmpNuikiAnjdUyJ9gyHhnykqz7pr/gPUOED/ocmAQ26XdeTOaqlHn/mZBJxv
0enHgB6fBsjUF8wfUBce0GhbqBTXU2aUX44sqj2VXngKEGFJMpBl/agjHNei2NKYd11r1jYOYTC5
gxtuD9EoQQF8WwaN5W2mgfHSI9rRrg0XmeDREVXwB+V9AXjQBAlCQQkXSQSVKGnYHd4rjutaoO2/
h5YgItT7XMGGZLWPwboR4D1t8g9PTgxNaw7/LxIHotcs0saXesjiGV+I53sGVkFVOCif6ngHo0+N
raI2lYIq7OX/VK73KV6mMXrQRTrGmym/rwo87aOI8mLpv60gnMINT/AV+lwVKVgHyOv+BrE7iHge
zM4nrj9HIDzq5iQMOcmuCKw2t1BQw2b0oWEwiDO50kWeC8UhFddm6fek+VOXdy4r7gjs6k5Iy/r1
8o9pfrCHY3/bkaL/7W2qFXRPa41aJliYliDwQth7xdVCvAO1BtmqTajwuRKnpngZy6Z0y5kuZX+H
pYfv7gHYSHbeLD531RvpXq6XIyUXy/67FkP0yXwQA/TkklHUhmLbQXh/oTPr/CemMIugtOrTEWJn
E9x/jmBOqJ46vpFArp8Yc1wuzPziKzr6RB6qddEtUL/BvVnm8johyz0NltaIQSCi+NoCQ3EJTlaV
+aZnpaVuy+r7e5UIG5DIgWb+vlHFqk8nwbQh124hNRjXuJ+WRBN+FuDdF08Gbr6E4AeTvn5+ifC2
EqKABQz3VvqYJ3YPl+bWe8ijJovnLg3ALG5ZgGpZpX5xb4TU8nJnrBYoEbBryjwhElS4VD6LEPF4
cI/hw6W+JVTwHFS8m5u3lcFarCNoFlsX8mqEzcHy2nagTNDGLjhdCJN2oQob6ecRoYSywSbSOM4M
NTf6j0SF9VqhpfOB/dN7u5I05O8znIIhlvx5qxg66V9XJlG1k0pPci6bFN7OPEJaAOTUuvVJdQRi
zuoWuaQ+cwLVOQzJRrHumiOnDhN+ioeQlfEUEzsw2CVqYSNbDbC+cSlDYoIfjiU/N/Ixjq2sfEss
gOC8Ze/C9qV+IKdqROZWVrAIe+fLC3wyxPOxqAFYqybNMCNenZL5TIIKBOL0yxeni2ZXXfGgkQB+
YrBLwKpZbb1I/fqc5iPzZWU3ITG9GtPIwt/CszFwJB53CBVl1mYpprRUYwZicDkzh3ohuMC6yiIK
C/+WP5W1NVwWV1tM666vSLLYWQYd+NqHojjWWkE11PtncsrNg4LiIWFUTy8VGuOWaMWpaU+efQcK
VJRJg8qW1tcTxYiZk+JxQwGRZ7s8gvDVjEr3Bw2ZphygrcfR7FRTH/AxEg73FRnISLnKyS/+LI4D
ybM9dQhgwmRCHxcL3U+RvKyOcXaAOKTKebmwZHwfe4vhiZ8QosjPHf1QJJzkV0TR9FfDGF3qr3Vg
+IfgsVBaMFyVQzAqx8J543Lobcd6gQxe8FbhVRVq3DgqjQfPZcuVL53V12LsCdGi+CmfbsCeMcP3
UUa0pDrEzp3IgoZB5Zo82pbnBZmeB+6yR+173/M4PP4X2DNFe1jfYLn32viJFcmfbhv4IiL1kQVM
wuLKVy+kMq7lbDD5A4oC70pSVOj2hDNUYmAM1ftrYkBFVJ3ozQWJIbU0Keob9s4m1NuRneXuawa9
IQGSXZ9EtTY0weMXTjhsTlD7VUjFZv3mcKvU/3C1m3zeYQxfHV3FQsPz/UDEUMwAMR6M8w79KeqX
C7znCu2wfzW/sP35OadRKFnDVqPw2obHKkXwZpL/2lIw0D1a+D14mBSsXKb3ysVrEPM6Ozn1Byp/
jhsNmIG/GPcHm2XAZt2hqaE9NMM1uHuzg9kx2jn6aBZiRFgRCslgfgj3IlfTOOsFQhrvJKHSq5yF
FhrTh6AWvDZKEGBvpe8BgtLdIFDTDXAHQ6lGILWf6xBiReiOy3ihT3kDXaEX84BAzajVwj2nd0YR
/kNeTMU14b2hGJsCVpM5AEPp4g9FhuTs4dK517IUjCOTr9R4D+ZHmav77RjlQQ++SvmXbcQARtPH
4632xTtfHopzRgHPJWIXsM+TpzeueQloy7kVim3gEwWqf7tbOLpbHy9IyaUYTvqqPv/Hn8dYfx+E
gNduMEZG3bCJFVeISqboinXC6NCkdKD8MjoIsQ/ztABZfof2H6QlAlKlo9FOjHNlxqEryPK4B88h
v7QNpfnDoff6Hmuzv9F1VmON/6/faLZ6kC6UUfUxJd9Vq3q/eqP0qOtbhJnnbnOMBF6y8kJXekjF
EWGLZP1/Cfj66HepoxL3Ne6cqJ6FzLAId2daqcriMEOYfYUEk5adUJSO0itEf37uGniDOOVIR/jf
o+z98XABHEEbbiY47fzq+dzBK10fu4GRAEOsarsbTVT4X6Sf6cEOYL4J3rH+iB+nFSYjJZ9RXmVz
5BN7qb5AAhffTA+SOWgkEOqgXaIZIBGkzN/Rh8gMWA60xW1tTIq+Hzl/ajLUj7stVVKDFRYaVqpN
LPZNPeAkw3BmnweN1HCQIuVN6J6uxAxvEDTps4hfQOQ9wMZpPBjq7THHztgxOTfNEecKnJJz9jDL
zmddQDDbmt57IFJGhiPjg2zJwABDDZQv9ylz9vJFzS5sDYn3Cc9iG3iRgYzbLPaVavkU9Vocjr0a
7T+AmJJHJMv1l+0sia3rJjylOOLgdh/RXsgn8uX8aA+lrE4bLYdyGQjAheB5Kqd/8Hsn/i9Vu5/N
edWK3/aCK0Jpa6Xd2r3qtCe3/p3mNX6UbDqLeDWRlA1Gc9fyibUwFPTc/GtK9MG/vG3wKXHfXcXk
Ayx0J4JghH2AEvJ1EMMolPsGK9PRJUzR0oZktWqZ81yCwrOJJKpyXICqJGWibHNFIEUjNP+078G/
zRJ0JfwKufqlH5Xq8uWz7+wVpBWkjC0v2IietHmfcgOTkmYze1RcB3HYNLsHZTAnfgqJlr4sNF2q
Zu5ixpub5qtyEFHjH8IU8Qo+lBNGQA4BJRnpIiwsTQbpZxLXwMq2uCZmCdUWtEPR6jlVJpOseIw3
N0nLegFGAEQI8uUmPzb9l6NSObddqJn696LoT1o2Zl5h9ZbjNFD+i7msfzPDtzCaoQxVGj0AezoF
CNeku9XrEGl1tgOHNn71EFfKY2c3mkHRxkUVGf5LjEIsyWSlFjX4NsRY4s/mil214D16INT1ZV1w
hW0o9S6c9s0uTsBh7KvQH+xwRJtjihb0RU0MFm7im9ZE/9m6Ls2aVMfpzJh723I8F7epo6oXkymL
YUJghTQ3FNBd+mkDNSzOQD0LEdVLaU6SPbbHRMQXyNuythWiJz5mThVT01ieQSvF2kgDhiaMIhcr
MFka9f3pXt2jlpFnjfwEffEKIiYZhHlSsmYXA98N5WQQLaJ39zF72SVWKdoe0fDxoQyi2+Yj8qrj
OkzI6Wl1rcKCziOZvVVnR+BVCO4gROHrfJrcLk7+LazyBbYRx74KSDrdud4lth3vIXnfTtzZWWZx
mKZzRBxSasoYm9JbAoPybODBYVubSPeWwvtTCry6DlQzXLmUk3horISpv/8MKUGV+xAzL3IEYSeh
NRmh2BeJ0ONiLx0+XcHaLproJ197t6b4ub7tHFTj41t750HsW30xAs57Aq54TwenQDnpX35si8eI
4vswJYbno2YfpTHxgxnpA0Z0hfQtCpiwxUeNyB14h7jQpPbHBjpCDozPbEeGwOwu5daM9kGi3n13
fNdTZuma3LlHvTYbEJs5faqvurxrgOaw5/T/lj5nDRptS3aKsFTySQASiLt0drvI0KQ0Tkaqa/58
/0ze4akO4EdHs9H/qGxUaD9DB2JNcZHWlITUJbWe1baTReCVfZJrgs3bl7uLXm+u8RyIOP+8CSnf
8FKEAGAXl5e7Buk9M/neBJpzn09NkMQnB2nSu6SW657Y7Zefaop8Ntfkpp+ca5abc3xwuyDAD50+
c6hti6TFidEWQA+0ktWA6e5q5UcVTeIv6Rfs+UChWd4IgqStuSoTnI8mKTl/87S9Uz/jkOrTbfPY
tPjp3Gp5/IAtgfuKYy5h/3JyYZ016dCYYbZG9TrqTKpgiRB04euaXZcupzwEBwl/WOqTHp41x9/B
IKAewLZGisp53dZnLFdPisam8Y9k4lnDQQJXr70o9kPloufSGfk8vFq4BaVSZa3HfEk1MT4u4qUF
hUAq/RkmDsI4b3jA+Tt0tVzbha20GlsH5c5lFqjZlclP6rihrCQ/aVmGSTeYH5JF1/pfyUN5ts8z
uU4891aW6DVj4R2nKt2N/Wwz/1xg68ONcWs2JPL3DSuedPoNWqNaWFFzKSiokc5Pvcf/cEL08XIX
c/RotTuB1IF4nhyCb0hf5GsPv4a7HSmtXIL5a5Ggvra6NmeiFFyXGDfJQzUBgL8V8hPDnpBDAvl8
vGI6IK9PmnGhygj3RqV/0IZXVtnLp9uX644DSe6aYslCztBr/mnNMXAFhH6ysWfQA13QdZUAhJ6o
2CnT0SOQ9c0mkzIvw8vjnkP2LEWFb8HXFdLrDu6hPOBxRyAb9K2vT5cgG431Wm1v8y2iJOLdHTzu
pv7ZXD9mPmVuuk2pRcXoeFmq9iWJCRFut+1XSx5QBIPqF8TLqgnyfZBhslepdhCn/CeTeeb9ASSn
npvCWMT6lonLfrIrH9wRl8Hzm1ew6qZGCWiqmA/DGjwv2cNAK/9HVv1fsw+pyEJ+ns1bR9e2z50V
jA6btxaXRjKqBIY3KSjekvqyqE9pbkv+9Z6yL0V1lwdMYEYJCzE3kg3kQEXDZyiqmK799ChIzg5N
znHFi3HDPEogiu6HhvDV9ak5De7UJti/9U+cAMJHBkeLzElvE3pG6tAV03hYPOl9K3cx3E/WExZ0
mI2oi6IM5CGSvWac7IKSUUtCtFXo1yEEhNNTlv5VnFkE0lSdKiUR3qYsNUt4gDMqV3eGX7T9tc2Q
SdBlvjFuPJy7KLVEWu+0yBrhRfPkSfexMYKBzec+puZFKpukyehzS/F+4ead6Ph/j5St6g6IOIe6
FeajSqeT4v6Jso/dGlN2eia3+EyKgLbK1fkTM8imJnCw1pQc091uXr9lQTndbq+MQMX4+KyQHJO8
VF61brZr0IWPBnUtPy99dPRANKoLdIZIQqpfbqCNGUCRltJGXknVsfettxhtl8Eo0lmXJQaahtHK
2cYm3vC2JxjJ+9PKg52/Du0pBlCZAVrxH/Gwgxo/UOoZ0bEBzUgW0SP3ILIOPbqE2eMk6yfOP2UR
UKjFWFRO5sP/AMv4K39ANOMJezF5+nn6/4S2zagofXUbpBgvdCMRWhrZVCjfQHcu41ePx9du+5C4
W45QbEkAy2nzO4POudu5n0uxZZOfKg2mLV/7sDv+qWX1l4T5DMwklTSLZEtLXlz9ZVjGTg6gMpu3
wqdcdRFTl5vKQu5tB9NLCtXQggT+8Wzi62qPEMqCRg3YNpTeQ6BVwsHAZrM99xhKTEh+rPpyU4j+
VBO9tT480IIBkyYzRlOQQsAkoURDVzs9E8zKbP3eWeXD08TOlURSzu6IhAncxZi6CmjFG9t9upGg
lXD4VM88EFuzTH7tWYLKQQyG77dB55Yemw/q6AiB90KgFeSgB4NKbFkFd4CApbPALI6JAwMqmZ30
y2IKSWVnKjJRuhcZUXER+xI0QsFlJjRe8q9HvuL5snCIIu93PmOVcBv5gK/zACquJhetqwt76kS/
NFnh7WYu4dZYQimNnoATdZVQcDW6lObsbrv/0moT3lyrcJbbxu0vNf3qSRPokOGSWFPASB9YEcSV
p0WXjKDtZS/MEhoRAu6MkEd/ZPOyQ5+YTh/+c3GYLzsXS9//FurKrTlxRJydK10b3SCSKFg+fdBB
XD4Ne0g4uRFBZiObZlo0wHvrJ7S/rENg+dKr49dum7vXvDt4Z+fpyVfIKMOpDw2Ja3vbOV0GhmRu
yLyG4RR2gRThWnPZLfYr37s1vmr1fzHsns3aMhu2O1YxnIzoep2IF+7ixEO7hcNCtU/iGLnmxdhC
TMTtdzxsUdvV+gXHaRg4PrFsOCfsCKGwm2gVv3DAoOhaRREGUh6O1NzN2CijITV/9Ow9FOzLzLct
MPWs+EC3jYJVaElp392kXSrV31gtpOd5Af1HdJTjHOweiOG5UO2XsnbpGzSvSV0QWz8izo3s+Qtr
bcaj6FXu1exYR9np8VvWCjAwXM4dU1BJsFYdZQFd8vrz5V4jHRd/bP+V2tUDNCYFcEymZw+pAJdv
kWEResSIlmkjm+PDcmmqMpYBmZeuLPIwPuJrls6muZ0LHdy6q4+icK5JJM3K88peE2V7jvaU+4M8
lQF09J3d6dgWFF/FXc81qhbnOjrB7fC6LSVoyn/Zvupwk+PiSgDspeuE/OJqQ64Xl5RL60YjpEOe
PMtLFgJ8a5zIQooha8LptNiN7j4uIu+Fi8g+ZZRdDcHqb5LXHKekXixVhvQhar0Rvz9V4ft0U3VI
nlpQlaHSjpZyvUGJ+3xMxgM20ZwNFCa3zNzWiK4wClhqxp8s+u2seOotK9tXNf5W2R/7fDsBplPq
xmJn6KdyLik9E9o9BUJVaMy1fsSj9wJC2Rj4Nf4UMy4Qq8n6NvXqpf73UpXHD/LK6Qtc6QGQNgoN
xiRfD3/9pLuA6I1uKWliD0mZYDDVhkozAmNa/ZZdbwXvzApL+PdeLKyi1I0fVF82pSd60LlpH7Oq
36KeqLWtKj6SuNsDkZ6Hbm+7f8QVlM1vmx8iz4qnG2Z8Ah+WaOGEyZTfaDJqqAlJcba+2IK8ghgL
jKC9WNW6C94sADYb24wK/O4MF29jCcmONH663zB9/VUHtUkcB1OBZZEjhPFgcvCZ5XALN7B92JD4
MO++Qu0bQZmaWf7YEZOfrVCp+bgS4JUFPCoyOtZhv3uWQpajQcXk3XnFLATMsbvAEdB04gNOKHpv
0k2VKI3ET/bpcnTDaW1rzN+fT1QAFEibRavseFlRGDlEdAE1nR6SIYkWgKl4BW+88NQMns0aU3Iq
23in7GVd19Q0s9ufnjAu2agi1iB855nRJU27xCVaczuwTihKzU7eLbWUx+qYYJdGYlhyR4bzkbDm
h4POyulIqQk1v3Dr90tqnrgELII3vqm8I5+zkmEdlpwKznGs3TTIKnWWJi36FqVlLjqD/ipDfdP/
/+ATs2AQnI8lcMDJlCavutlt8Z66XsM9OSTk6WQ76KqqRyi8JkvN/hRzKykLOWjiW/IvXEZxOr8f
bDmMq0H51A2ol4dA+LkgujCSvez2+PKXM+Oh6bqL6PHkbmVY+ZEgSpGp4Yen0Z4xFXP/L+ZYTfdf
Es0w/Dne7wz5B1lKEJGMEAJI8M0zi+FRfs1msK+ltQAdR4RXd8Q49zxC0VwQNL/K/u6jK45fqB0G
Z2rv+G+6rT7zG9uxEHIv7fTaTJjijym+Ki8I2WJxfAi9IflQo4cvjynaOaKcVw8M8I+gHb4+g2u7
6zSFIRojD4KXL5hK27bytAAAWyANriyn3VyPdvX/boCyPL3tF0jy3AnKQXizY0vw0TOo3EoItLof
HN65r+55kldZzOBxw8khG1FaMOn1Kd/SgQgVbL43G4waW2T659FP6IE7LZNwGYqtNtmMX2R2oF0v
zJ6T6HGBFFsgc+SEbPGQVOzT2Hep/5AzQdqKbvlgoykl7sskqlcavkkR/Blu7uxBe7mBC3L6vHDP
OmthYByAYy+UM64Lje+aeEo2YKm2EvevmzL9xSn+ufyK3V0FfSMvSsDZ9+RGzCUXPK2DUFlGTlgN
zsDXkQHCU6dpR44/kx94lOwgfYp1Nr0zRgCJNJ30blgXiF9cBebKW7uLd/J9Oi00wCNnuM2+NgoJ
iEKJ7YDWrCyotzRNK5BjUbnvnr8f1V7AsUVT/RW93iH5q622L/DavKMqPTwyNNbiPsjljsB/WXS1
mIn9Ncl1o/ODU2sA4LNldoLY6ADxPyMKQjzb7OW/g+aC4niDcTYZ5Ot74LOuipvObTPRFqJMp4r/
IrAs4iVh/bV/SOb/oV4ozSa/pb/qR1+ygPSdz+5EMo6fG463jDTVNMa1eDziLh1z5NuhSOu2ZVts
OOFa8Ix3oUm+O74f1ZL8DQSF8Vk9sx7BYOXq4Jc9PpLcSuJ6oG75+8XchJmPkKoM3D7DVQ5+CiLE
Hrlb6VVxEbI8OKcnyZGfzPNO5j0ywbptggdkl3P2m2TY0WmyYe3jfJyvbXXejGiWdkpu4IlG0foV
YDajdvaUKnw+rDyUpZF5SX9Rv5RuLQT+t1EE4gA2IyFp9q7OdXhZvNhtifTgUwDtyeXoSFYMODIk
qqF0aGQHYb17ZQBH2WUHkzJcwYITO2nzl5N07kZMdmcxIZebdDX0HFJusBNI/zUdxmQy8cpwtzWl
qHPKSuv6IjLZIf9Qmgf2C2qH+R6lQhKSQCPU1qUJPNPV3uV9E8WMQBoGv7WexYp8K/2/FzgKLl8R
R89kHM1sEFMR6voUWye7j8JsLLYIydVW6H7bvRXUtUb0CX68/CblqLZ3o6KfDEQ21Ez9Yj3LuRe6
nqzderSxvpSR0YYmSk8aVUsUzPYRdOjnUYvAZJqCIEP6mf9n7DbmseFGc9DUH2vUcOmKGbpo02hN
qFeVR/dRqXR2hEn//nTechwOZSoIK5Vx4ycyF0KFnlJhkGQ/3KMN4BOUP8MoutQ4LkmnVcvGEVWc
n4m/L+HKlIYleC8WvXRH2yTc+oPhZbt3iCH8hz2YatssuhX2klacnSox1rZTy5ai3eN6hc3n2X59
iQkXmrtmi53MtvWGnJGgXmd2DsBsXual+ERMxX9YEl1JBcmzQQPgkUEy0OsAiDLxHrvz4XeXQygC
TGTP7dDxILkXT+e1etBZPac/YC/qqF9/BH+0T2FChCo8u4hfu6zecHCWrdHEa9g37gT0scNAy8DB
tXH+fcz+iMSobYyUaLNBRNZSSABqOwGh/lT7sQU75UGui73rTEe8S+fAuyT1C0cI9BHr/GT5Z/m0
DWtTdYkBaJBZ2Is2xaUJIBVxiKe7JMn0ZB4OlzLlb8wMTr4x2kboav2hjk9k6ew47HQrZTJ0SpvF
mVD9gqrMJYeyzdlVQ193Xs98c4X0XHbJ6aLNazkr/NWhBG5j2squNRBYzTJldBOj9pXOy2T/dP1p
NNb+knBMvq58VZkgtJ+lyjFJJdEjzVnFBgutRIxzSI8w2w1DXr3v7n+iWsD/mChMIVR12Gvw6bV9
OREkPzqeVMewDzrvjr1bWIh5yRDkJZV6aR/0ZdnVW/mHxwjayofOsAgHtvDDPkKnI0c2I5YwQ86q
1zMuLYeqn54PmesvGoNXRAqRICjgIDTMTe2Dva2GY4WI2OJEyopX3LdD0frbl+aCfAqVD7ZbWVyr
oYygPIslxzeH601IWSHTsgqpixC7iYfSvQzGZkPgbU3npKaWN9mfDqblHMHKnNgMR49Gt1eWxWYF
CvaHnCHyw+gahn4yQFD9FDMN8DoWrityeG1tW57hSZmgley7X6VGIzVXhDt1QLnr7ElDEtgjhImc
KgREf1GgpXroqcajUenXYMMMtoT0yWZSfoqUm8PHThaleRJabxszrW4B6Ab3+iFUTozbuBwcdgln
2BUzkvIk2FC4QtfK+lHijlP7HCygwKHA4i26OPAz7jQ+wawpfS98Z1euC2sbnpil9iBMPa87tRiv
5/QXvcf+LlZk0QZSdXozpKtX4W9CQ86JX3K3uxNKPhoiG97weyFqjkhZW73wwCox19GEorDj9ez5
HjCsoZTmDzgr1iV8u1KKtpe23HC3XtwE+DKCQCs5wJty0Lhhk4C452IjmwFstBNC0csjqqEb0LAG
+nBhXN9VVQTMbhXapquI+RmBLIb/mGDh1SIrIrDfuM/zRF8C/MoUbcoeZOXo0n4Oc/Fn2a8CiKL8
u7iaeH4kJkybPw9V4dUlIE3MQQs3KkBorqY3dZzbhVKsqBaxr85yPJuvIbfQcVHFgmCBwJWR7np3
RIwW0uUChGD75Rps3o6fLpFeNg4pKj+XA4GfnXbyQbYOd+bof97TlXK9wgkgErxm4I4qYNCbdB+3
SYyeEjJatCIAErwLkJ/RATmH24GaxAMrcYoBbmdqUILJOjhLK11RPZGQA2mUDQu9GrKfU4FxsfNN
0hPvwAmqDfA/i9Gkw0lV+Vomr0KqEQtlwEiPe5CvQdG0VfXcatzYtwjETkSeWFOVPaDL22rioKCv
brGgnttPWP47LPYb0k1msUc1MkQIix7xxk/7TpN54dMpYBORj8Bw4+481RQx8rJbg7pH920+SM4C
SmGI5/wypPzTZc2iFHVHTCvbmI8STtH+HONCHWwWgu1QdVnjw6UKNQpw/U/WiJpudoe1Vfaueqir
tuwESftgR5LE7QT8EMlIhtLtbbRBdnN/bZtfmSZFXRjb3DhgBCeyuIN828KgFy38a9eNYKSzeYqa
EFUJxuID4iJSWmjQxfpwjWwEQi0YXcMZVLYVox4pvQCmb2Sz/jFmQufKjoVD3Iyd58MQVpuumZBf
LNStsQworUPFo59S+bnjJNdqdyBDAs6I/Zf8J2OEqm+rdpbdNvZIRjk3ExqVufb19JAISB47nv+S
0Zrknhyrhw+NVv+QSKvLcZRG0XrlavN36WvP8PcxaMy9xauzBvvq6MYvxK5tAe/xli9pwl1/ATUF
g884+9qfF7vnjo4ln0Hjc2jy3WQ0INYHLRseefys79Z87S13jqShYlH0ZACmRYOsrPxnlpmgx5aN
l2X34FurqWaWfBR958C0dKAe0hzS+wWcXvxBO3PfmIlVRiDehXZI6av+KD0ppZ3c4nC1fJuAc8KZ
4fPylVWznoihDPLG3ejKc8/q/yIfBbsmnfiCPTsnFO3xxO0H+4uf5uO2N0u1ER6Zgwy68Zql/bmN
IVdq94gHfzn0fS6vA3DJdL7dsajJo6+cFqpu9YahJHMOUnDl39k3PbJe6sdb34NwxP3+3rVLq+UI
Uwf5m7Yuwl/rFeEdzCPSQLxus5S9+6Fuw9qS1GGtBfRx4GFrZjIvvV404F9v3iPU9xo4qw/yxImj
EyhyRdpOqRKjfGeAh/pi/emjm0Zz0+eXxlF5aeUuCC/K/TVah7hY9MaB29/pT5pBOckRWpVS96tM
yT+NYKjuoxZsMSWD9ue4bM+L+dhzxSTYmnY8HL/JfEjyEDD99fGagECRZ7C+0PAKN7+ZQTA+24iP
NYVFMFGinMZ7KvuW5u/k2Px4Ep7E7o+J6wwPHWZALFOiTigvjyCBEleU0I+T/8TGMn4uhItbNEqw
oKIjEW1Hea6jS4FqPMLGt8uTlaenJX1QmYUg1UZB1p51uOcavfCmFqrRgYTgnnqN1/7G2ebEbNDH
13H2xM6f3CGVZSv7erSDD5JZ4LBkl3MCxwStqTWWkxm0AFB0MkcCrh6dwrfphLeYxXulMRrkkATJ
0b0ViMhKHGbIxXbHJhqNwF4+INImfKpT6CKb7B3wGfwmdtmGf8WmAvjBuqo/rbfN4Q6/xA9f+Dhz
cmlBx3OnTVZraoTGb0fEwtzIYknpQF9ew5pPOvV8rWBBIq8YZXhxrl74wk9xb3m/LOD/h5GJ0mYw
mGsGeFUamYdV5guOs9Rd0eQzHS9Jg+cyjWMhp7iMZ1xbccQv+iGBxAsF15okXQmhYRzZUXTwQaeZ
j/1jVaHCEED3KI1Gj9IsT3zPa1+26Hrt0+sU+pf7qoXqNb3GWv7MXgZ2fzBH+Os7Hu1er6VCZ6nl
Sa7gFBVeClAn7bc1VooCS5w8QGHEUf/TaIa6+rG07xivQms7OYXXhmyQBUbOXVsCIbeWZZiT7zL9
W8OoXBPKJt2VuyJqk+hVcvDjB6UQpxsFBpDDEQrsOFDwewiDB3kJi6cfiCNAkI8d5q7aAsjt0ANS
ttuBVj5p4HxQWRHydVl+XMTLlLdZOzdfVgbqrBv7nW6bmFgtktGtLAlrvdmeeeDBeAeyxa99vPWq
tDGiD9lUkBohpFMv8SuJbyJEkl+VLjPS1zYtJontS18NSLxrPuNbRDK5sz6xCTfh7KCo65Qx+fzH
VMB2y6rvXFmP/0YVhqHSyWrNTkWqW67iWtxtd8xM/SxNwPiFJQWKUkiRr4H6EP0ny8KZ398HSMpb
RN66KIbPxv0Pmq310ZQ11/IK+4mbjuKm/8dwm6V7Dw9JorW6v2zlvfAnWKcdhNtWb2Riw5TztP8g
xsQ0jhrCrHa2azRvpVccvNe3JoyhSMU02vzcUUrWq8PXPtCKCgRH8cb6Pl87WbISrz2hHcQMuY9L
C/9KTmOvnXS7fwlaMjKdfFmAu+gX4lOF+iwo/PWI5nI2S6iVMDPxmLjhqRc/chfOxeIj8fH7K3Js
u90DT0YQpbR2KI36LdLmHVjquovJcVniOU8S/BpFttjd1qnfnSvMEgfZE4NOsEZY3FJVyawXl7vO
GjQ/Z+FReNg6pTjDdE0JqWTBJtfVC5d6INIyBCGQi0pvdrW7780ZajWi08qU9/YBqf3ssgd8WnfK
ZYa376wj9zjH6pNjvH3F5mHXQSCI4CNOssP9eOHy9H4aW8hBnohiUG9NC3fsq+iE7DLS2dZ2bpFB
RvDy0v/zgd1fryKXJLeMpCaWUNb0LgPpK/zIdcrFHRvlIpN1Ga1C5+3Zu6prx88S3KLmsmrVUYdj
0enHtU7ETJoXSGBZYzMdOaoRtDsFQao3h9UojFrRKR0ezHPvSOdGyJyG2jpuEW/nkJ419pfY7Zvj
sWBoVqvLewPij1u8BpGu5q1T+j3UIppYuaNjttRZXG7e56uEjZ4HOe3T2Foxj8xQw0WRiEyD1A5g
ChX2G69zPpwtTlrTAq03GxEkIiQs2uw7mb5LU+CUBc4cA++/Y8315JIgWleZibx8TnaBMdxZ8lSj
YBOAhtsTfDkVcoINoDVh4YkSVxHHDRJJh1lY2/6EKxo5R7GN/oVszVk506Gw6mLROBwpqbE+x3Sb
RZm15SaK/JnOHVrb0X2whNEJSsETI+UXNdDpb4h1MvDX1o/4bOhvNyBPFn1OwsAvh6RrCoLAy/h5
N0OFC+f3l2ezDNLi9RpDaHzCkQvT41fRCFJs7/OgRQlf5e2y2ly00DgOh6GRTPumQpCIsTEgt7U4
3/wYlPnGWf1/g8sePk8EWBKJCx5sD0l7pYRa497vErSo4OyQpNgxgK9/KmLQD+vX5uDmTgFNK55z
T1GPxG6Eyn1QGw6ZiFrcP0JWQxZtrgH9CYE2+wDF6X9VJcH7KKfKPvBKzz1Z+UtVXZUCZ0a3SUtM
0hOmZMa1+gobP4c0X/Bm2HuVrBpynJkhnjAaF4TuJA1YABRB7TMZFxhqGHNUDheau/2kAl73dNAd
Yte8lBcfBTrX/5KTCARTKISOuBRd4Ckj59CO9mBKgBqN/xYMEwz6DAZRsOjqvNsHEGMAfIKknamX
s54KMfItg+jdIqUr9sG+/vUGn5M49RgzeZ6qte135LS+fYzxaQI+2WaTttPbet2ntumicarobHps
wSY7aKJfpPg3MbTp3ifWDXeam4MLtAa0x6jkYNdTCvfKzfyNc+A9zCAc4LRAFawaM1SKXrsdqJZ6
Q5TcSqNVMzYAPiAhTV0r6eHg2Hpp/UgSw31TrEJ6D8Lw9jA+NGz/SNXgTDUESw0GBXLDABUx0vZN
rvWs9/3w1/GAN8he2VKVN6dFpVne/q0Hm2zZm6vRC1/VYtkdVfOStwWaJhIIBUqueK4vosfrU8L0
45N3y0nRT8wvJ8N9ILt42Fb/TjYDYJEsw2rtd5juvRufLYK9CV/exfju2z9Spz3r+tTC5Aj0fyIW
sG4PEfP7+8P3huLt60FDyyWaeQZPTD+vS3V7HNstSLag7+Q0STBsyACREzO6KtM26r3Y8t5UnwSK
+5zIQ7w+bLnrY33DjKkT7aTfwaKwhpzhehUnPENqshV8N8MYpzfJtMfUtJhrE/jZw4dPvQMgvOef
8nVZKhJGgl9NdoLpMeBgyeqna8ZucV0mciqMCEVEe9wkuGrI83NiHDwn4o+j+KyHef5pfuP2/xBS
b6V226NUvsKWpRQPDzjERoJJoPbIGgmJAPQpITqQyohJW060imfyAN9W9OMlpLZRAZyG2iZLu3F9
GNin8nXuc5UKSw0z8ns+dw43f+Bw/DVTAuQxhmv+filq82kZeSCGY6aSZ4xR34quWfMKc6X3s5wF
d41D/T1r7zpcVb82h6dGjKTqWnAk1Fnnu1vhsbJJNnAnDuYS78LCWAIGo8dcY7gHZR43D33YKCp6
QSv54RAUiPaSD/x3jfOKvzXg6VI6+ehFsKf0qb5pAhMiTTqPFPtfifD3ucZcCfk04EJH//Fae/be
mHgzv5y7Fjiurw6YOCYP5c7FxH5z2hjXYVD6Tf+Df3/JAyiFonM3JX0+VaezVXu3NOhsRiOVpTz3
cYhXstnuSsRcpuk2lgFXGkoG3mj0ITBnT2Om43OOBIAkqG4/5sIt9PyK6ikYyfQo84VTOzGY0CVk
YrVzShJaMr4WTyPp8l8vjFG7ZSy/De8rj3dNBtQTp+G8ZH69v50BNjaacteGYCfEtXRElcZoxb6v
wOWLxvTmApYtEoesUeq6wVZuPuBEaWnq3W9o9VSbIq34yH/PuncRZ9cI0uuGfr8FUmRgBZLMii4a
dFf8UdfzSI1fvKr/Q0+i/WupnL7dBrXMfz6KQahG1TqKyMg5S+dYWnHv2gTUJ+txzYb/t/voo77P
02RIP/eq4y4sM59KrSQV0U2t1Vo+5mqPZLlBJNo9P1AtEezj5iJWCTP90N8tgmMRwXbr20QOKxR5
nukVFyYzSmBdh6ntTXVntcN4FA2RSyL92Y/i33WeYSZDH10QvzqZuFrg1JuEmRGJeI7ti5t2zdqf
l+FSGxO1AS/bNUH+MOE70ts7c15cCuYFkAuh63ea8HjLKVCUiUjrOICPkznL/OegdQIrEsRiKjxz
KNPtMc4KOM0ti1dqoo6fGXgqvwR4jxTyJcn59NtnvGCwN6ig74sgVzn9l9nVVQjjkUW9WxJ9yy/o
Wz/I1ZWUFy3xWU3+2GxEFa4hifKc+NxU99i3yr2bKnpnbBEYaysqNdZYVyPa6ro9bOda4RWt/nDO
8iBuNJocRzgjwu2nk67EIdWqBIbs3CtLN08bTVJMj19jg8+8FLnWkpRudt3Zc9MuO3Oaa80DpSjT
v1QSFzcY4aI/7TgqWf0zRNmL/Aq2krXuRVckiWxpqKdSlk3oX2OE/M113VktYZpNMKbSUssU61y7
ppiv+3/Ays6YhxX0HoYR7RlWP+V5+DrIyHHsol/ZmgVzECYII0cZb0oGHm144FL0m7vWe4fsb5z1
FhHpG+AhLe+L27OWxbO2D3PEKWL1eQJRfvO02EJanVCcIgEL9+Xby0U0P9BYMMl5wplvNkjN0mlM
pRtRkQa3k1GEW/9DQtJOgrM1Zgc12JQc0fSTbCLPSEttxSpet3sV6EyjpocExnTihnZSBEP4AcoS
CzA62Ey5g0tdjEuDUT7r9orhxNzYZAO0L+/b2LHm1Ns4qG5qSBY3G8imCwyGfXYTGh2+Nhb2IBav
zVrNRT6EJzVeYneLgqFbfHt1QP4mpBo14urC0g3UR17RVtv7VKcTEve+b40hWVF0odgsTMa44GTA
dxxbTeX9GSQ3yIieHrTY7hrYtxw3DE8BJZl0fFC2e5SnHucovaQAXs02Gr2Xacd5pBCP1gr5wpl/
CIG4hmfItD159h0HLZTlGLaDIOaMBLNl5UuWk0j1+gmM74XnY+g28aVsyvfR8H4cYK5rElvR0CKc
nBHbJTdO3kAcm+hx84Hio0cH8bbea3jkX9/QqjozspyL+wLQ5v7zmuYkiCzNY2sD4CI3EJHFj1Qz
eZsJog9x4BxtD7GeyuxBsjICTOtKhMMR0hxf5f8ZL+jPg1t6EedSTWqlv6NjbZXqM+Mf7I7Eg/9D
DURnJ22LmYDLZTx0+OicPt9y6U+AebbboMROaaLeKLdedGniliAmfVq2ukUK5CUb+tM6IWeT9Hj7
UrLM4kyYcv96oO2gweBBWRT9iPe9qG9QaM06Qp/boDpHobWDR8I3T+wnItcWHkLN/KTCyfygo50M
6yGpySujc4DUGwKnMScaqdE6oS/fXRz6mWjvXx3xHYY4c8M6gVwIa2kLQHbLcgfiQI0yULXPhx+H
Dego0x+Nm1lpjMPfb14NV/dKmY8VtJsMBlKY71bYhuWNXWdA14BkSfHlCK/ustk1msTrHyT0NfwP
Y7s92UDT6R6WgwYSmSBDQtR07JNRONSzD80b9GM70v54/iGM6lHNSOnAcSm6xQSWstFG3XbWNXSi
c7SIJ1BeyiiVadKq9xnBUL5fjueMtzw1jWyfGA9t7cIJwBZpSLIY8+4G3Ap6ub3+36EAOatSGaco
/CZv7hAM2B2SUuZe30pQr4tMPurLLNtWBha1+Gg26rnbbtcFMaoj6+L/UtQASrUvNjHoK5iK6SHV
RcgHPnJDxIKvab/vYGagesihgmsX0nycFDp1z1SIiiX7lP7SgasQqpwnKASpHaE5I7OnZh067nWD
2go8cQfHfmtc9hO39Vnfltq3ZjkJn1piMH+E17SwLRGHPKjEIHd8DwKsbz7pCJAsqGm2VPYVdPfK
ffbsXDXxYhJoFmEFfmnq7RsH27xF7OUXXmBrL7NTgXFf7pkK7B+84yx9ZATfjj8RvW5PpvdmAy62
KKpWqO5evxIKdsYipNdANlZ3GxjWCBThV/e/+L9uCy50WEWJ3bXoUsTPC9WYfLVCHAczB61YxLQU
eD+rNlT6mjV1k6OzutalSK8oyIje3uBRdrvTxz9uVD1FTCUHRx/adHRTP8vM5t6sDgBtu3urnS3p
WTNkOsWSzE05wMLiNfMO7uHsrCictSjX3z8tB03CS44x6nlnwbCQ4Tg5SX8CX44hM5syqQwxeHtt
qBjj2fQRLr8bxdRdTC134pLKnIVo/sHf9rQVCv4f2O2aqvCcxR7I90fGIov9+GfqIv7UawADan6K
3gc5bD9GG8Fa4DK3oFKphyclHiQaPBCrd2sxV3o2azCFIcZXa3DO4xuz4C43kGe+LFXCYMD454JC
jLDYUwxybFR/CunLJ6j5s702uU35JY1SWE3+/sFSnNGoBbGN/ynSZ/N0pzuzEEKsCtaNUSZx8ZnF
oeVwrzkR+VAVxfOKzZ8R7UbH7X4nFYil+Xsc7g8AqelYxzZ18gDrFNgpYfXwQsQC9DuftZzRHv8E
+/r15/ANvfQ/+6Ogpw8jLczl1bvjC6jJvpBHdrIqo5hGhjL/N0Xv0MvmRK1Od8J54LWChL7qyF9c
PtaKpaNVZZenkyxOO0V7bV9UHq4FdHyJYOjfTbECpOM6J5+epdv7nZPn8SpG7PGEqhOAYNU32CXX
WmFso10iOLzBNlX61f0oP1epNW5Qh3463vetzYa0TX99aGuw+tUz6iXYmRnRAL3dcawvVqhqkBnV
QiDyqYZG5AgnTuhrbX7jMbiFYHFIpZTPZ6V88cZKVn1YxH3DofPzeW9WAjOZ2kpEc4+LSdn3babE
/QMAQ+nbYBcFFwyN+9j6ao5Fc4UcyInDzpWZ1ft5pInIQtwqVVINA+qtstbc/bKbVQoCLrKn4E7O
+aw0KGwMV8Ash7yL483agAyNqQD8/eDTnHG9lcct7d3jCfpNim/8QsgZFJvcWwa44HWXwACP5zTH
emStX8CxpwGJVi+Zx8LM+G4gixLWptdVGVvcEYfCjWZj4bCXgAg+VxHzkYNArGKw9Erx2cAH8Q3j
8whiCymJBeFSZ6A7aFxjIZGXjiftjBtCExcWSljQQdvueREQn56Cqr+juoDv9p8nXIpFiJ5SsSHh
j2MRW33uwVJ8xJdRrAwtBXScheJtNmp+gjze+cYhppharLUKMoBYXhz7T6H/SN4cArJn7dJBD2hb
w2Q1z4sL4XNRQbZoYIK2r+XD8uh0OTcO5+YY07dYLTcqbOy1JNBgiTA8VuIyAeMa5grOZyTwh92E
tOxpjvsg59Bk5KIHFWASnJON4+bUITIg3dAhcBR9V+GX57KWBDHlCKg3eriIiZuGwQEiTqTOzRl4
UUrw9lhxOe9+WRmzNYliIMe8hGJgf00D9VsTf0ubRpnh4pVtLfzCUT7jesKwqIaFzjt/pZsSXAtQ
FZf3CoMlVzxrSK51/NvOdxJxL9kBvqlQCJtPLFUhFh7Y1xts4ACmYZHsK4SeIcccz71Ycj0sLqbw
CJTedGfpN/Ht2Sr9KsjlZbp4Siy3DwQq34U5OzkiNKLaB/1IVTW8RXaHINdD6ucZWHvfr1InZXZV
h75fbfpnjsRRpDVU0lzL99EbJLbhEUcE+YqotZSil2i3K6mTlQb/+2RufKjhO+LoaldTSTElGOiC
NYd7GIZB2DTCh2Jj7/qwW1+al6EjQNbMO6V17nmzLbW72fdafQ9KHxT6rQUZdHG3Ffky6n/M89WQ
8N/0b5gdtvgj6rvJI4X2JOLezW7iijD0b83EerWr1eioxbAhgoEHZy4fceAJstIg5i0xgfciujGZ
Qag0yBW4z2gDYO3iKi+OBR6r7UdeNhcvoFqb7DSWMhHDxpFReWwzao2zGdLegPJMinnhje4WBtEq
TexcqqVwFvAJjD3QCMOMk23K4T8BPvmEIcRdhfDknHplNkYk/4SlR/GiyXd+4M7BYQDTrMXxYMw+
Mn5qhCB80ukYwPTVfcUArK2v+P0cfWq46DF5MFwJFg9CNx1vZUQRFQc5ojy3F4T1rigdHKTFDFzH
ejngNOKUjta5p9I4sLYYp4gQrElJztQjtFLj4eNoAvYA+TDYCKw0aGhDvcAt8x/X+2NWp3dOQWj0
DXEcyn5iCL3xlILvYfDDFfz3Luu/gJd+R+sMsmwf9//ObMWIH2D8AdTUPI77dYvuIJb5nQb4UFhE
8y37eLQF12mXP0Srut2vExZov6bZYBUmr+0sdZTyXXYbb6RnqZqlofIRjDsZIVKSQgs8Yz9+SzCh
RuVXN+4BSzcmAfwu5DZnXETGoLa2NjbSzYxi+XvTK/tP/sICsoIdpAlzruSwy3N+2L0AInEaZaIH
qgt/S0ES0LpsgetNYANium4em5BSH1VmH7D1Etu2zpgRMZTfEnqtZRD1VBP2e5HG1zTr9bU4zadK
NCBQw147H1kTo6Ca0Lx5UT0ghNkOgY1AF+F90n593XEYxfQv2gkzjuug1otnfbWrr83rCw9NsR4K
pquhjKH/j0EKQWb2IYQ9cQXz1iMrJm84EEa1hF45Fjm0rXBC1cyUtPBN599iuOj91HRFr4RW1VSL
U/ZOJ5VZ0bJtVBc+REna6JKkeH08/+gF+H7wGrVhCQeFrfj4/kDuY/vd5OZ2Z5qHO1bL7qgKLho+
sCGZfgzZyBH+3QbTlEqYXlvud52v9mKXjipL7pruoCLSyN405yF8OVZtmQZYeMv//6VqOXSDYudo
JLxYN/M5zpcnFP+esoIMnQicp/8vCnmD5YYnT4g0MNLgWVUH5Rxm8KReNSBxW8COIpGrrhsqpvyH
CTKhNPr2+vDpZy8HwY7a7pQTQ/eAk7RAuXTq+X1VWRU0i59A+EvqEQE+yrGCZE5qBvvkg4XPLYIk
p4bPVPLivMMfvm8TabKHV2soXATrgDOVbVbxRjaDCD6hawMFs0XjPf5+lpSeW3nicQ3CT5TP8c+q
uz5TvMesjs33YiJ8IK+rr8UV4OA55lrPAlsH5WOF8QHZGwFvnDs1hR2fIHLFxibdyeloZ2umP7ru
cVxqlpGQ7Eh61sf1nF55GgKrzgw5R3lPFa4bpmQKc/MwTFpvjA/gvqZUwCMnPgT88Qp9AVVVH63e
BcX3xfUmEH6glfFjIkpNQRyVUmh5tI+T9Ko0SM79+DhV0ksoIfx0WnzRAr8WTNrYJX2qdwrm1M9H
dPqRhGMhr1wD6CWjrWrNNT2OnKbqaU+xHnDV33+ceFDk3XIhHRoKONt+6O2XkyRrXHMWu27zqqnK
jiIGwFadd/ijMwYVfkVPcoDIPEjPjOuC+1lW/lNTzZx9b6rox3zBhlkXuQ/kmaHLKxc4DqRgPNhZ
3tgfWqRFzXJ3LqrQ76zqN1RoraIQSwpjI73ja1BucpLlB2R1xCkk2KTrNR0JE2O5OgSxNUnL4rVo
Tg1wcdFdXsyaINiFPMJUpS7Ip6USAVg4uHHx+mPIjoOZFG0dkR4QH5VuOVzDFnxLaLoaxO5M2wa7
VnbUubTM8Pu3fkLDRKcDJkZliftuCbdGVbIvXZ6Cnm/Mhx54MFnVV5BPByRwvvEPeKNgNXMBCu2l
hjBPriIQApHBfWfvUdDRsfc+utgR1P2PZagkDm5xNK676BsOTjuhnMTrYy8jZi5WsytR2Q8uyXCl
+V/1n1e2OE+Th/0MtgNNSqIUddTi8oDnO2zHE+4Q6pIaMUY0PkrSoQENoqDMFUJVtqaaGN1ZGwI1
vIuE6W/YA2RiN46S2aG+TgV+hpIDZ5Xwr3AMvsuGRKdii089uTWFSIMnajMhnjfC+PIjiur6s8e0
YUseC0V0SGvl56Lk8xK9IA4a9A223bi/lVX2rZ8/kwGWXBi+GzhutXrFtiDs8s2pgleOudD7Bdtk
B7U2+esHXz3WKCCdyZR4sUvY3NnwJs5kuM51thHptBxvXDsmSzSmFRUSLTEPsoEaik5nYk4klhZo
8edEXHz42jbWPVunE4OjzFz+8sNx0seTbKqarUMbWexfFWGeaGS9NhqGpMEDNEoC6S/6187sOhJY
HGvtHR4PXdspBVAhWR8E8MVtIuMimTDF+yEetmC8Zjj1M96bpeSzkJAUqs/NzwGCnXBBY4oQIElI
RPQZdtFOYhSNAqrHvWYUi733epG20OIsgjK2sqk46E51793u4Eb5/8BR/OWYP+E73dec1XS3kWxK
ZqUz3EP3AnaPbLzpEr/f1WCFc8nXOETmtmIeFPCQVjl725fb3ppUxL4bOk9M4mVSqpOnXpBeMtFe
fdLhWig1XHyVidUmzG9wbBX03ZT8Kau3hqgC9W+PtHLwgzUBI90OC8Uxa9htb+igkYMeYg+U90wF
hUDdpAY3eaMsuDWHAcxCFuT8jrsg+VNWZPda0BnUU65kOkmC+zDCxDiPzialfu1uU8GXbtZo1LvB
leJhiZBxIyaDAnG/S/PFq+WLzSlx5RNweA/DljV56QpLsO/zAJBaGktkKISYtxG/e5V/g6q2EUmT
amRkLN9sBwGFLTXeT48IY5TRd80yEW6Gb8OBQ9LVwVB/ZAkaabgY9Wa1iWjFEeRjI9bOGwIPVfPO
8PER5qzmHQ/A5GCVNopmVpnU/SintoxoYCIELfM8fQLbpU2R21Dhv48Vswim5O5lqqfngg3WiW0I
KJ9pBrc10/IJcIyQ+jsmWVpCA1gGu50Jbd/9zWVUYVCnKov9nnmRUUd0XWcZefhhe8KC3cdxjcQM
pfUCKxJn0kesXBTTffPI6n998mfQxbfToQPokUpXGvJOaounmNn9LiYD1AZFA7rR0orY2O8gcTGf
+/rbZmAZrQEsafRmXdAkBRVaanACNlN6Q6u0bORS/9Ev+lpKcOXXRLlTmnhqE/IZ4dxlQcMM+JbT
0ZPqU62bPqAq6DNqUkB0tkQYKSdsQZUmsx5k0DiixEGezXf2y2GUU27ZohqyqHSgOqiti1KNyyIG
eaQpxqeGTl+KKRnxHvP8sCTyoypfUyT7mVcF2IwtNKOY2edqSJG5tPoVkVCTGNzaSjdx2jWYCW+F
GewqvVBVYWPVTw1hbDR9LIwsIGuYZRGqwqgL5lbD/a/hn9lPL/Ndl8/KzL3EfWUNB4MJXsa2uCqK
8Omvg2yGD0wuoZmBHttY9nrTL9OR+b8PcvZACI1FNLXBIWnAu6sRSDvUsHlXIYKUHkVAzOEpDz2C
CK+x9UTLWv+ZFF06YCDU297p0bIpp3GuHD+xe/juVPLwx4xPf9250/kKYqGVPbVzE2IDxTtEbNW/
NXbcG84bT5EMdIL0jxZtMEf1YuWS50Zfy8QIAm81Ni6AQ+4TWNDkTmE/aJmKdWhvlkqtdGZP5dzV
1nfcNz5kEkuF8/saVWVTHb3JbYq2tCtjXZdAgDgP4pB9Pes8x76YI7wj++YPyBllsQsPcBx5FFk+
29CHIKtcBTPBjNAAZmeQHgY0VO3hDamuGF8RSB+/F0poUhRGPsBwyHk0Oox18W5YjZ9JugviSpe5
VFkKuCGSSpJSobeZX6T/EtJcyzbcGp0ZKt6PUqtxZPnLnT6ddVBe9AN/CvNmEcacTSuko+LGnzpv
zBF5KUnpwJemz6ZpQvZXZ67DhRsrhILv8bXjxBjs0pSm33EbEs8sT55H1NCPdo35Uael22Y80Z4c
2HwS33fadiiPBwwcR/9jJvTEOH4t+LNdb8vBV3ctm1XcplVd2COicbR9xsANEmZb3hAI8AmHPznM
1SDuF1A+GaWI2+XqBr7mlC8PjjJWIK2g7PqEgK3MoauSjpeeUU0/M36uFEpgZnJh/Qb5ZCNUD5xe
m7WohoH41aB6n2h3ofOutZKVblsPcsZtFW6FOl7Ch3XDpPfVjCa1lvMn/iYVpqXbZc9MU0x/fqXz
PQoDoLw3WomYWCAUIJe3CvLpvRgfsrQ0pDRfu8085txDi3j5/2u404RBzjrIPVXzJ1YQ7Aj/0bow
lCQ4LcWz0GcrC24OZimq5XOVaekkM2hy0URZq8INFIIGnmzSa6sdgW94MxPDV//WNoWUCpu/T219
JbG6N05U5BkHtU8nxZNz7OlRIZ1B43/zYre8aBfz+CzrrWReMolQczuu9nVbpTei/exAMvWqJ9tO
AhThqhZde1875pPzyFjuuGLWUxW/JysxpetbFHJjW6m9EvrZ933HbK/xa4mF/5HUV1Lup3xJixG+
md0gnXXaKwE0hd7rC8cQMn8Up5GpnDtB+QxXO1OzfhjUEFgr+/JxeQOHJJgQ8NTuA+R02LJ4MLoR
mTbgG/0guNbehptg+Pn9qzzoZsNZ7DHYegiWcXhbKohX5Bw0ShT2cFKDiAcPP3ftHYM883L/rrS/
LQbKHX2YechZLekXtqFDRM7aEvPqMiIB7PQVNf8+cgKlYNkkWNehv0EZ3fTDHHb0WQt68zrlxC8F
SnFBX9UPzyU6uFqHGaigzCjvj4QZkrlkwL9kdmenH6Uao0XxDFZQQ6rmJi1Mcw/9vQVoLgJei+Rg
029BcbSNBZOTUpQ6F+6rpsl/KRLEFQ44bkMqh3PxntcxFx5ubqlV1VQzDmeOI4lAx8VnXNHHEfsr
OUBwEhEgxGI7tNemO3H6KqasYXzi6m5Q2wXRNvZtinI+0/PZ68buy8fT6hybI+nHnb2wpGemNKKM
4mGMMERKsfGYxgmlOysxEcBcg5TpW3HpwVCMVqkQgkID3WgYq/qHg3t9Mag2I68GtdejZBgwPO9j
x+WpOf7ul77RSFAj71/wAsRXUSh2wQx0NQpauxBEDqCOeLSEymUHTNDb34euXCVqPGTfZPMQ8AEF
NRKAHM8i0fvkQ0JTEBI1wWTT6K87sGExwKQd/wQQozlpEqCkdLACn0FYNINhulewN4iMmeoWXMHB
BIfaOK7IhxAK7suBfF6vG06ARwBYKVSJoaRwJzzXycIZpyIwp0zDuqqNUWGNvQ/FTZpw1pgOcxV1
sQSYG3aA00EzRi0u2RtqAt68lA+bkjPHQpRt8jihpd+Pf/84g/MHv3DCIldNZD4N/i2PJm38fIWZ
TEfuwTyrbJ65NO8AGzR9hubek9TjVqOKnmy4y/Hzz6mtAfz9EpiEziYHMNMutdLMln4maBsoBBFn
8hEvl0JEGXbkOT4/d3VYxQwk34EsQffkj0H7YqLxiGQ7RngDkqo+011asP7IsLeuKkJ4wh2iD+65
s5wPH8izIpSIbLqeLdMslTn/cfAAJn5WwedMx1QjlpToURvdI15rmFJLh4DJEmkSikaGihV6Qu3z
+mZnANRzF93ewj0NZUC6miUFuYcJ9M2wr/27j8jnW37zI+/mw/4qaJN348JQORZYSmOf6RQ5ZeXS
eM6s8tBuXl6N5HnAqe9XecmdBZcNP5GEyMY27U7W8qDuxWb9niBa9dObysVvl3twZuZLcXtYbUXk
ux3Tz/pHGKH0/nNCZ5rplhuDmJX2imkYd/ZYeqsu9L1UP0iQ2vHMuaY4uqImj9PgRrgw0g6RiHJe
Ui22OWIPJhf9WzkE/vElB3UQ+a8jDkG1nMsYzCw1kF88nRaanNGc8ctoQap9J/PtX0fdARUKJfed
R5FcU8kigd8sW115+rJi57DrS8S4cEI9DY1u2PoRztLuuFOLDHRKaDbdKuWmDJdr9eYo3mGoh0JZ
HyUfpq8sOtIa/KGaXT1iGPXGj5AxmzuvUfpRMgcuTZj45DPxIhvVJsbYtqjotChxGeadxtNX1CAr
t98BwUiVkT1/P37ZPSmingoK19AidQruSNQNaRVw//KY32//EaTamTQWKfBJfhKRQcB9A0nhkFIN
CaoZOTGhcr51JL/nzQ6xEFEjKzjdsDFRba3VKea03Ajyt4DSIxUpLcvKN+mWVRK/X1tXX3neFUF+
Q8PJgZritfzycfj34QoRJYMnTYR+0aQe7wIvaiCagWKGD8dz9b9NAogsXIlWamXLSYiI+QuXUkTk
2ZbGmsDdmZ3mPKk78a77++HCPM50JpjVYuCUTSlgZZsUw9c+epEriZgEh9hB3mVybmGqdpUA/+Hv
SsWPr1RvW8sj7qmmMxPjo11Y2P1p4k5VMVXNahJutar/lolEH6lJECYsAvkhyXCGFWp9r50dvbj8
4xnIodXr3/OMtjAGTMbOv6EjO1zKpcJTRTk6fqE1s6xwWYnTUKyVqWCehBeLHQZYA4HT9xk9dDPB
zEXY+heGJ81NIpY0oKa0Rk8PDN/paOGoDXsBU1eBopQEJbIjR8/taCkdHXKrbYCtuk0UAa8jBNa4
4UJnw1oJUCRjiKFaAdghBk9BSclHd1j1ZpkRnKkdVzj8Ga/3GrZpXruBRHYnP3FXTkXkAtjhYd2X
Wb5eAmEJUCSUiGS+8q6PTmi++Zqvak3fbHN8py57b4z9Y7RQuN5WU6FVxbHvx9Qf6J4nWkpTRlN9
UywhHvSIGdGME+a93wMFEg7Us/l75y7pr/7fISATE4ykW9U1qD5yd813mBHQJUlNilZNZXs67eks
NAzS25bKpug1cs+jzqTP6NkBbpWSX1Fn07raxlzFPV1EwYj4/LCnusrItYQgD+Fb8tSx+5J3VnxX
ZZ4qBC45IgtVHpChPaALU7YuimubrPJWJ93pU68jP3q/OuLHftTO5tWM5oAn48dY5Tu0q8Cdu4Im
e84VqHI5F+9sHFRioULL6sBscKCF+iarkXnPsiLPcD5FEKn9fO3wZPdgCLav6K6vlPIl+iQmGKq5
j4himM53xaq4BVcIlAxjpuBVk9HYqyaJ1pX7kULZZDKxgkn3LWGoUedN/U6Kee0eO8RwPC6fq7oJ
JNxndscuZe1vduDnbCH+oJ9joT5WmbNfsVA9+VPuo4Nhs/jwdP3VDKVp9UhAbcKs88Rp6GB10LeA
JTl5OxD9FY65Rx7c3+VAY+DxKF3A31Bso0jAi6ToXbr3GszidH32M72UQ5i/SCyH6ffKiaXiq+o2
KWuxtr8+iXS1NSIXvvnwE2FAiS1XQDVKMi68IIB+z1tuDc4Cnjbz3hyDMg1bXft7wjy5wLHRD8K7
jHDL9PIwbdpKQYTJzoap5eSvWCxl+Sjh3w487bcbAByq5m5HK38fGqNmgRqEgTuWMYbCaVczTJNx
ZejrGzsze0kRP+4gZBfvE9xRB/VsFaLo+frQn4Fw44890y4+qWHZQRQ2XX4CHczOnXU4qMnEx3XL
1VBb7GC2CcisDj2+skPt7BJ9MpKz8X9WIvVgTv8HDYarl0BpZmz1U7vm1q4f2k0vSWijUBOcxhSM
0M5qz7f0hAOBsVo9GCrexi/OjynocfHzio3/SBugQ+jmIWESpzcvLIMPumtpjQVmABQqRayW5qeL
eCV404BFkYtX/APTan2Ghj3t2zOjjDZ+370S5AAc8rM/eODQAGjkYaHstkvYW1UQyTJcLMYGhD9N
SD9NnBqwuoa3QMFjU53Vmm/rpjapGjolm84PGO7C9bxSgfZZ2/akwbSNiZGWgxa50iQ7LVlLJ7Dd
f92bR98PeALaPp7UHs5lN54fjH8ZtvcsLZk3WoD2SD7Zoz+9H2ntBXXGOsJM1No0DYIzEaJL/1Sj
mNlvL6l0By/8zcvvtmMEBx7kM3UhUeGnKN2XZz2aRfr/tBJV2Z4rBlOTHuH33oCsAHbH59EZYTjd
xATvnWrENFKahSaVt+2apWTv4DtcbHQB05mX4MKd2esgK3rvj3INBHuaE+ULqVmVP+Sj/zocAB8c
vRD4t1CkjWVKWhsb0UiiuZLV51yQDcCCDZ/b5W3yf/1QI7E4T0w/08D/A3tzUPhJCA1JnwXAXrcj
AzB9v7b6GaXYtI9a2kUn01woga+aywFmhmqLsow0JDDPtu3BFjdtaCQtet4YLkPAgS/hVYmFMBom
ahqaGQYb9DBIMW1gS6GYSFZ3Hgp8J3qizp/L65W+EwUrnQjnSu6xHO2/6443v1RW/XAlKEAgVIQq
RMOGHpvHj2XjbspcExdxFvkicXrvBZ8XbI0+8XR8ARnQr41TApXMoa+DPJ7b2DrDCEift9H+DfAV
Iz3/dH2r7ofb4ICrjMsWYQc39ePOq8qPKzWeCEv1MoWeIW55s7u1uWXrKkokQkxjisq7yJO8hHGL
F1NQ5h+4P0Dc7AV8TcF5qJp4m3GTK1etzW5P+P05IWpCqxq0GLa3dxmKzeIpvET8aS2K5nR/KV0q
/gJ7iph29PG+NlfWxL6Kltmh1BtzMheoRq1pfYsqhSQ1tQsH4XXGy1juDC1LODuh/XOQhTdFK6RZ
w3OU83RkHCX6O2u5d42K2kS2w7ehacP50k5l3zNESbgqO2h6FnuIxBJAAFE77AsvILRaOZ6ZNkTe
kiVcipB3DZVb6Bkb2IoCqGgtpbakqVUBwC1edTFBXW9WsqrJvt9ehCjgGE7bhRhzHWwv4ZR8zACA
n2Z0PL5MCgiuH282bnk+W3IQ+hU0GBBSSHHeFxjcAzjlHq5xJcMNdC+6PM7NGfmn2izKGA8PATZL
g+ufKFqqNixzBc9rj2UTK6xlRTcxY93A3IBYac6hAUy7z8IrDBQPT+9ST5hL1uxWBxW2cFAg2IrS
wTSFTs5ozy7hVWk/Y8NttloFfZLpGpnu20TKConRwK9k1DqFvU4kxFeN9I0v7f3eknf9Awdgm0uU
KCGqMR9t7LmhUsvHYpp+p8sbvQiHHSdvz74MTnm5JNylzyKvnp8k2qiO48c7iX6V8KrRdX40a7sv
YQKgMb9G90S1fo0qhZx592y/wAMFidMzHi5Nk3q/NrGxwBDSTo05S1g0F5HW9+HIJY4PzXYpgA/B
/y/b5JB92Yezgll5mUtY0dN0IXaW946Dz7FrxtsQG7KExm//s+dpSugJhKGxGRSeRKYtlSh/oQGf
uq4mgZDTDDwLl9IEHBLKYNx2FIJtakNhOTk6n6cyepBrIEOtH0cmtfYtveEQHJlzhHN/ZnhAwbKn
+tEXHG6bu49j5FPgp/IpBCFupGHTIUZpb+dHn2EFxwt6zlOApOG7SliF2toFv5RxDjYorEtztV+z
wqsjizHn8HjdYSQ4f3CiSR9DwZ69Cq6jTMoLnIwl3d481QI+3LgSPiZuYJ8XgzYlHtoPSSNNsA7e
Q+0HHLaUjE8qoA3XnZV3cdJ65OTn9nvmfdMtV2evItzpS9ignRT0aBXWmMc6tukeVtA0Eww6lYUT
KvAQ/RHI+1JmKTA7VFyjG1Des/TAWow8bzxbe+id7wgKKoQZy4IMtIzk3s/IR2NtNygF041Mixua
sg0SEmrXyRmABWfeeeK4VbiSZ5eu2MnY/bUy764TSkQwdA4+8zHO2VYtIbQz3uzUU5bBeuW1fga+
ghEwj6Q6M+K0fxTLjiWgEC5Zp978snIuH9sCWGJvwn+PJyT341SQC3qkB3OH3UkXw4uEB/7t93Tj
GNHYYqnzFZvZEjONBFJL9ON9ev4u1zaVxBIZyAWBk5IIgiHb1M9UXcZ7t9FRGpdcC8jC2lp78pqK
4H6nIze4UTsjA5GX7OFpRikNbU2EHRjRC5biCJykTM7XUU8wQeRbZArxDFYSpcYPrSmajcHb3y99
VFGYD8W4Lz8S97hpdz3P9bbhlXDQfhQWBpexhp74ZrA50XFbD4z3aSkNVZQCJSzNf1UJ7gMKP46Z
b6sh9wq+hHolr5oq7TYI8CdgBWZJg9Aa9PDrH01J2LdSudYy8iVvAhuabbG484eAmCd6YWwq4I0C
jFDIt1f1yHeoxpMqa21m42FnmZfwDVs3hcVn12loWCHP1YSUCcq6sJdiMqcCT11Z5LrFe+F8AF0j
mnSgKInLBSRaN92DUQFUoxG80nKDDdAAtE48NIVWS9GqwYM0jMBd+CX7WdIRdUuHj0vTSNUN175S
jM6ykJIY6wm8nWw1X/zbi0BflNFRMYzC5F/EwGlyg2EjqEwcZEYc7rZioC4Zzd9c/xNUyqYriq5H
OSJScNXLu6HzQJh0u1clIdXuBtt5khOrA7K2qYzfowbOAAtehjXn6gb2K9Iz3y/41e9Iow82YNvk
6jRpgOW7OxCbQgeGRlrCDQwoKmEBqeUxtIceoPO2mc5fExsIeQeUeLiJl/fRgOHn8aWjmwOzmj2w
jjP6/OAf/xy4o79YUfFMyyp75eZDHJFQ53FDZhTjGebLjnxfio1xlxIDFVADKLAxEOETuIye28Wq
K7OX+UdctQrOgt5Or4F6aKy7fXuZgMldrQkB5a/OEDIJWOoWseoGOsUwT1fu8xXLpVF0qIJsY+Wb
p3Ym8qEaCBPZO1N/q7z2zeesUdQP/6RHnrpgxryO+2M12ZBSgUtT0jwqVFT5cnLIm1hR8Jaz1lvF
9RE2TvqlQEKvOgSvucuSdgHhP+U0y9AZuSD0BDSERYfWhMzFpvSotl/YWY8CGr78wY8c4N3DypbR
dAGIz21+2q/EsH+MYcTn+SYgbiWtLPBBMkKnEs3s8wjXa2BIqr1Bt7WmUKFC6/qMjXRISiQFkl8J
yKV+6iN21CpQRhncagWcc1N6jzvIf0WSIPgodYe3Q0G6G4OFFq+ZQNnZeR+0HUasbJeiSo3RBTfz
1RuwQZEiayzqwuEv593HRJ+C0i5La+Dnrj2la3CrN3yFQUox4+JksBHrg22TR01fEZekfWtCzuTA
3IxUeTA9JmgXWGXjS4p6HTGp2rWPKZ8TCSUVtnS3m49M1HX0hN2oiikVQH8N5KAzYo6lRN9HpJer
ZjbXSYt7W5U3xCirLW3vmUOae3KGEntaksrNdVLEbnR2jv1DlsXIMzQfm8FmTlo8cLo31hULMqm6
NMlHJaaZpvDpm16Xaq7TKK/0Hg4fq6nefP7yRyF6ruLz6ZlgNJ5+sI9YnW1vV4+rfTYR+5qwWytS
41Sg5uYcAA/gjg4erAN7xpaBKWyY1965fq8JxacqUau5slI/VMSEB5RaYry9DmgOzQrTujESEfIn
6NemCDC7hzDnO/a+Zc0+kv7fm9v8NVlKkgAXE2yXf9xWQw0bPk9rkpinJpx0vPM7o4F/uwtBmlyi
xlgiXX5v1lI4+xxp4VXug4eqKTShjMbtlsFO8BuOS0lgX1YDtEKOBEm7w6GP+yXF+yNP2VxZxQvG
tsAiBMeHBTY1SgzgFieGIktDQFZW29ZDAy/IKRW/8Nv3s7ARl5cGf/uN2Av/N3D+95McBxiLNhow
MVaZWfPrt3rhDBhFA9kILMerXvijPw2GzQ+gnHj2BGCR035d6k4ibZI4xPrbndwx4ARmMuiS+PqH
YnKmLODRO35DaDvTDRzwhLd3POaHfbXugh0gqpXCdocf7LI32wxvxvUTQoOt64vFvjyF+hVmRakt
OKeC07TY2jO3o+qTRgT1yhKrhByFvnohLtjXQKxKhB4Riwoumgk90jBjFC3WPhNo+JtzJ7SccPep
TV/hcpn4cnivuK3upt2211Z8psb5h+PNvYkytmYDonpQJ4jtw/qNPmIT96PdrMxTGFWhkAFFek8a
oq7tb/r72zlu6F/dE80TSyqdzZCHYREqkHleJIl7rOX+8DNQeIzY2d2BM7aULREH7PNc2HS/VtFn
zzV8h8IWX0nWyzyFzUxufqtyqNIFRptpwYNQ9MU0r9/KVmxrjBwn0v+HgF2VZ6bVPu9ca64Xkrl3
pmZiS7MR09rt2cSjXC1yUPplWCN2iDK5X5mwK2IJAPEdZjsoMjyMlbTTvATTIGlB/ryHlPvLbDZg
Qx77VDCE+pSyrf1h38YPDNx9PY2WSKIsybjkhzxhHIeKIuUIYYOGNBEWMWOcLB6aV2k31tN0kvKN
HSMyieMPeBmh5k58TNs9j0vGeqg7xCdCwsghYsDaIz/qT+OPHW1Ca116njBMspnLHp0f34ULWJVW
/0Qrra6jt76l7p18QUJ6aUJCDUPbE1EwszDxRlS3ffPmYgIaiqrzVHWHg+OrotaO2MfDasGRLbqa
egUN/kTVPMMO7fWeuoF2/aTPUTymCfuvBCL6x0cmzHWiBZMPa9bV1bmWCwvsk0ZsdCGlxKq4M9Ec
DXXfYNSiCZ+2BXtnZaa3fQ/ytxbmLGlE6dxKzpXVSSeKxHKEpaypJJkJqkhp4XN3pAhdAe7aQtrr
6Omj+1xLu1QRqcjrJR04u+14N06C0+1zbhhemxfJwOwr/oJJndQIK6UMRF5Q7/VaVzjN68z885w7
L5Yl7drV0BrTGdxXqSF13nQUMp5c1uwpSZcFhF0koR2Dc9m+KZRFCBeuvm1G3H42A9OJr7Y6EaMb
ENfZJkyOrwTwTd7VvfvPA+GlRhJu2djt0PWYbTcirk+qxzhGtQTbHzzMD0rrW1JjQozLeh9tuACJ
++wIWPY4yYkAPyY0Ia1pFCiPvv3v4OnF/xvghOOv0thCrvzrCGShBxS3EB4kmaa7N77/2AAFS8V7
AnerQqns/pRIcFRFP/zPsiffKkIUbBWHDjsOqPMHmbvLvX0JieNwSgqqM7FnVzxDbvZWqqMCo2eU
5joYc/YfzDpnWYD9KHotAfXKR8MbOf360/V/Y84Xu3ze/WoJShYPGN2m3fQQKDGCCusO3uP8Fbnr
WV1cOzaNuT7YlXT3lK84W0lEURlJtJmmXYor5rbOJK7mkozFuuHG6l0sANh107r29qyaxJQcTdOs
ZOVU++NlNpLWBRkZSkVqDcR9EgU+ZMQPjjJc7HE1GFuJ0wsON+2i67RaXNa3lM8uVVpSl+d5PBG+
SN8B0s7iVSBAPvFXu9AawkFA1FSv8eW2bFWfenmis6+t4/D0PJPxtnnZR0fCCcMDngyhVON+t0DH
dBjoYJOnwjbcIc9UbD5SmeruT3eE3d9FBYhjMgR4yd4uOxk72Xw3WQL4n3di8SFo5NLCeLhmwT9W
CFvis2nqtV4CJgk7ffZAxr7OWMLYGWhpLclti95VPaqJqli2m+NEjo1H4zPj902IpuR4ar17hgwq
NdZ2ZOscZkjAb7wmudBQiPqWQ2iTS07J1qOGAAKQEzMFYaAzhtPRdl878EMufI1WhPCrKLcvaaEa
GCrSNDuj1EGGzNff0ef0wkpbhV4LQkM9nbqToKgKBRcBTVbZ2Okh+y3nAiFSfLV3d9jZmHCu+eIE
qDXzLzYYc2jCSg/I+hFeT7IS146AbG6Hir4ufyM8aJnHMNsJ5GECuPAH01WMbl5OoX303CSzNjkz
S0owVa/vy8Un/lSfCx/rJiICwSDc99I/RtH2WMCht3StjdGi7GUM08oNcMGLvHqIIPhIZ9JfGbJ+
FiFgMqa2OYF4wqvIQC2LSn63ME6zxNEeBOBhF/bFvVhhFHPOCPg3Ogx7SLt1d5sL0XeHbbDjbT0T
mX13FV7LiArb4w32fJbi+GxBR8OTCKB1cbDmqWjjTFo2gHGyYIt9q23NO+avyN11hFmnPiRUZ+fM
TCc+LEBRSWWiyybmupVQCIfaqqPlynxcqeLIR81O11WqN5NxKxK+T/VHPhuQalWNrXvRgb0yRZh/
LGmruFJpb9UFAqh5qaqvl5eLeW1y1bSaKjivTAWJG6eVT1g2Dmc1DDyzjoQMR01TOSRSuNFKPJyP
GKJ7V3W0sJeyqiAAYYlR+QUrPptBXGVmDVB1kgVAEbRUkXTSZKIF4yWgvSD4mjgFeEhMcoGevCFm
RZInDlmfy/ZrUxOggz9d6AUcWTZGsB8+C6BlPIXSQoBXfQZC2zQvvSUpO+6mG+fEscf/sEXG9Icj
LJ3HuZtbj97JrVfJgyz8EYM57XhL95EHGAxyCMvYqNrRElQ4tqCLwZj94ASyqheO30wgnAgXuFxX
6o9MfBzMo/ov/080CClJEjzbHiO6GgfRr1E/XZ7gKwNX1QUCH/LvrrWxBnnwhenyxK5Jcs3ol26z
fuvp9CP5xF7BVsbxxDhCStzhn+yetncG4AQ8+x/f5AOzihq4YPkSsHSVyHj7cck3dnlu457VnGxh
zSzQ+l3ZlOSl6THzkUNm2D5EZg4isPEozzWnBcs44YMDli2BunlvytZFZFfmG1ZvYdhEdJcrEBMc
ktFZC1W1zfVr5Vc3+qjAk4XSeVdZmzIrhMSjMrtpj6s5l+8DiwmPfQSOc20ldAyjkjypjHdhnmPJ
LtbI896wuaEbvg//xXUwglX1CobeRKsCTnE6A4Jvas+x3c7kEGncY0AVflwpfBiP2kLm2uXKBBZY
JqnOJIw9iOhXIxq6UFpwDzGNLfSTjtdVgWDHbMtws7M51rTzoCUbd85i1PuNPgkgCpNdY9TTFPgk
rmxNBXZ3EP5YK7i5+ZOfGBl2mVE3Ky9Q4Bx95A3vlX3blZi91Nlm7eEEJJY9UC56yV5EJ7sKFvrz
ZncbBwAlAZifhzX3xKRconL7PhtskSNk56YuZSmplfmNtDZViF0+74sECs66mFfTRfZWkNdvGclN
byCaO8ZcVp4Arht41RwMgXQa+WbOORjU3r8eH/Kfv76QNIhs+P3NMH/K8H6256AGTKW4Y3C94qLD
BOsf2uh8WCsDTDmpv2jWGos+sEXy8OVGSxxlAhaz7d8OWETSsv4mWGesOD5nhchlsZAFvGKChTEs
t8QGCSh7+pgcaSs7zJkav8SHfuWOL/pkLpvOkmI1ZkdnmFOZtu0+FekyD3Sn6j4BQB+UZV/ry9Eq
ukJzb4Qr+AwWYFX70B302QUN6fuQPnHa8EgtuW/K9NVL30OcvOZCKPdP60C1TiAcZ20YX/vYP5NX
cYtP+EqLhWVjneOXt9bPo2TVvF9dyDx7+my5MGbNxkxX94RQmDj0kk4yQ6IPFCUaJgDTdjviFfTm
O+SGEWhXVIW44qqeNZXMiYF7pPDwVAesHlt7W9pIIqUWTmJj1yfFqnLwZPv4iXSajJ94GtgZ0r3Q
JlqL097iJ6nXriq8oqM5Dkovs0NjzGSZCDgvJC/bzwlereSHav2/btl4GxVFyUWsAoJCVmuD1Cpg
9Dm4Iy4N+72oYHAVknbq2w5+iGD+Ux2vJnAmMETDXp9JIytO9IlGw9oJnKgufqDKV+8/cvbPI/4H
MkGSLvYJjVvUl3kRhSbJhLdHgdYRg9U34nb4MnxznUfXPmZvCz3r/k30rjueiqoX9sZTK5ls+OO6
rxBsRhJAqGxD432Sanxfm8alFisWKwL4lMGtyMW8Garyfgyk3+VgDQHx4q/S58yjNhAeSTvRclvJ
4qZkPocQITOMgvAJOEhNg4PurU2LtH9nPXclKvYypW6vS3DxOTch43uz9qHOTBwXSb3RYj9jyQkt
ejPhcf68xfug1GgA6iZ6tFtsRxgQFqM7aUPhKvN5fixb1R/L6N977JHmrl6fI3hfhHcacqjxdTHv
GgEYnBQ5L7Fxan3p/Ypb8li4kU0nC28HJQb71b8P3qy1uLgjJsAtbgxNxPdnrZvforTmFkivRokz
+JlBzi+AKhRzquXBsCgzgF/oHqKf+pDN7VjrPHRDHGTOaLcBDh/HUex6iahBL/SY7RB9jv/K7EIV
OM/6ulheEu/cw55btB7SgEff81wn+Bo+XKrxKCkRPyvJzeRsyCzVkztmdPnM86F53OMOqzVEDKLp
ZFDS3E7E0p+ylwW5hgYYNxYTxOovT9efWZkcQ6NCmYz2eUb3c7VW0tOODO/jW506guVF2PVHzkAm
etIPOzSdmawJ3EWC8DKovvQlvLwL8cdPtHZ6orOr18GrcobDz4ibYWWnvgruYVkMsmv6ibYL5bBa
bExaTHAfAQdWuoO+u4s+J+O7p9+nVgVPX5KJ55a/hKwzYRfobkrwvcHw6hCNfLg/CEwrDNMD1d7n
hLvflCQKUx2UgNxuwzhHT2KGMYf6aVb2wPYJ2Y7TXvgPCjCMGrxVaL/RHVdxPRCviFMdx2t7Q8Ws
J9ouOtJt/mLiUY1PTSATj4VrPVXbXsr2F9xxJU1757UPmi6skw5Jc5nXACLiH7afUbyeLKxZD6r1
idM1Lixoa+PzuPu7/pREHedxYPztA6lmV51yYJdrfc+Wklz3CDlkInxbRUwPzr5qJYGNh5WEF2ob
aWKTPNYA1DWY2UIO2a/ORSEwh91ejbdGjQ6YAah9yLhqFIhnmAnxUEWr+qUlwck3mFoJd49Kr3FS
PR+rtgmWC/fOoxuUZkvYOduWq70CCRCOXN4qwl+XrUxane+syrdg7Sjwc0KXyY7dNXvnWclwMLRY
WaZBTOXTKIHI35Bv89i+BQRn4TnVrWKZyT3wnv4Ev6kRriQlSDkWiRBq5nl7AzU1aDTQQuAXUr8f
mv2qNm2Lmb5RtpHtoJ30akisxwXOVUqBbYAl8BbAIk3A6SVvwHi35wNl/xbvMR3VDqf/EiPFNbrh
PBX7OYbe2TuF3qWcqlmOpKBECwaGubfIen3u7MAfUnCtYMuwa1FisyOu4k9sf2KTvKLO48kzR2LV
XPGMEsOqFHPP45mZ4Wy/aPiJxLD+TkobxSgKCnaHpUgb2lKnoinsceIdu/7jyRv7yjJqGnV8exPX
kvXg/XFkHjlXA+XVL9st0Ej3azTa6/mV1wgM7EYwhYuXtehJ3WhICYjXnPEkgBgV9eSz7ebOgxSi
SmxQLR/b074/ntu/Iu0RVxvqV0QwEH1TJQx02n/056HNjILW//1+2JGhkNNXHPsI/7AjaGtOC413
axvsapxu3/lqQMRz83JOhPH2rtKi7uWuhExjAnmEQlh3v/njY/AzSxfj1TaaxhN2AaXe5kaYFEtU
5n3pXZ78CZmn9YscMWx5SlW39NUpTk51rYhnk56AS5F0H0+1jFbw8/b3ztmj/4zoo708s7WR0qTT
XIqbl0OgqrtfMVDAZg5NEXtWNoAnyALrJduD/1Wf5VFkV7ytcMrzC00h8Y/UwW+cCNIpo5ZIjpay
vVI3oSNGSfq1Dky3oc8xrvJWR7PoiXc9oEmty+o52kTh28JNeJw9/qvTlBntOfOXW35HnzsZ+WE2
PphlgVNEiB/6XAzw6mrrwBUL1be/OjTtdlp7naS56Lkl8MiAXo71CKQID6RJnERJ4qIKFWzrQnLs
MKhapIHo3S0HI6praHe02EDXvN2Bf5kG4JyrhhAHnMEcpt41LdHm9DBdBiDg2v2PzfpoogfYo+zc
j2qH22SOBWCwp/breaUhCgNPizjVXN1/nxcQi0JdXrBIEw9j17bdWjI7Zcydxl9yoE2I2wRpOjQO
ymIUGWwhXQT4DUfVVZpIFNuLvS7oNTVRj2h2LMRk5+QpQAJIGxjWeIiY4cTEi8LuqD0HmQk7CaWq
NA29Wii7/aC6eDLZpmL0/Dft2IHoxGI82Jqve81YICBYtdsN3esAp6FAc+vY8aFXK/YJYtpEfhs3
oxn5KTyGZq0YKdTeVp4te1ZCCYgxvtlpka8Zh6xsyA1b20X+RE4IZ0/ANt+6CQBE+yLkAevgN7+p
CNrB9jtmhXCBJmqyCKli89kOlU4QZK0dfv4e3udY3BiZ7CYS6xPDEl58QxEEIBXeCpD3DGoGiM5R
l04tNDLdlaQMCtVtv06qy6qxbzTe669Ll1KKk6cclp+aVV06d0IpUSxMdtASsDpiZdEOpnt49opv
IhXPFiCncfZTBo+9EXDZ3oZL2xeRNRTMxrhet+lQWaUv7snVh1duaX+XNwU1K+UoUjn5aM0PJV1t
eopqwmR7+lD9pP1F1pV852GZ73b3GYDU9eoJ8UQnAu4Nybeeiomby6RBG4DG2RjHpnTTKHfeH4W4
A4ElcqCh0AYnnnj6SQNUhc3pMWAxCiI6R5RcgstbpK7Y/eU6DPLWL+gKkk3drGDV2J4LcysC3X0t
xUFhT9ajSa9xKL/C3ERaKQTYCTNFHCUVSxS24pAFjCifcnCgLsP/5PZNLXGhOUJDV1YlAav+pNwF
CrRJeQKc52Zwp7bCtD0085O/oc5Cny7OFEWxHd27OrxRfGCxwsYOiLUcCrBsWMkREZZvgRkqizLY
CHG99P3Uy/suU4aDKsmuqAChhkek1e2PO2ShprD+FQWT1NbW4Yq66tYyJytWfS+51kGuj3CpjRp0
+g2V5yZgShxbvFvL5kC/lb8SAptvsKN7FwjVANs6/LYwk5nKJNJSp7BINmfaADtF3x5/D/9qY38O
QciyAznBFvic9MjtMpcoXOgs0WNSpVIOpcaqt8Ec7aTrcWdB/8q7zVtF7KJjKbNcQ9GZKFTqedkN
r7v5AWywCgarxeZMXYWgNbGJwAZurtbcssGmz4EsPC6dSDiecyMnfumY2cKeMb8qWxqlrjdhCjtd
wCrdRne0toI467PRz1Q6zIxXYoUN+YLGLepqPmcdIgc10Lz9LH/iSstBAhva3Jui9jCyOjOJofqt
LClQEpO1Kut8WvEtYydkhdzqIg66cTxxbs6C53/Z41Cs1FC5JGYDuc+H71rG9U13PWYqikYb/toM
R6AReQZyEjuZhJZmKGbLALHfJ5ZftbvZJu9W8CsHMMFbHsZ3GCF7NMmOFE7IpjS4iYbD9CMjy8PL
DR/0kB7RA53zEkzKJAgrCpmHK5367t2O7PxG6xK6q7TsDHeovsdvoIavS61rivq1nAhpYivMvLA1
7vEesE48TsdIoYAp5bmM8xu8L6u/clmOVZmOBuvGSB5vwFfdrBy1AvlAlxQtUp7XhYw1kW5dQLgH
SCxsC2SPO8IbZMVMIaJ4cTFbEdQkZ29jFw+oUVAdtUXSXJNFjj4oYQ5hAWlyUDmbrCdVzBgpBRWs
nZuNaTH9GZ6oK/Qld6HKKx48Y7eEHV3HG227OcgjaC1TeRLxPiV7fLFWfv8KP+bchv4wcpMPSkA6
9xOVJKWHJ3BDF4Gi5DudZiMqjGEpqX6hjSll6uo3nHHLYCGc6kBFDEumZ1eGQghx/R3/7aGK3DVy
4bYqu2d/OsfS3RJgm7WmPEOXAooHpuqT7NY0HRyzeNId92yLSLuCmv+XYvAYGX0mHZGJYo42T+FJ
yPgWLGNieti3zfinOZpyWwRF2Ez6p1hvsatwkbCMB6jngJS6Ni7TePvC2zZBXlFhycHgaIjbX/Md
IQbl5pm/o1o/Yy6IyGKcDwMRAzLziolqajO0U8a3jVDmyUn92t4bGof/xYh3IdJiDSbKYTUMoFkj
/j1b9aKpSAHZaB6d+XYvH2VY+v+2Hu+U5vBubTvaa3x7iBvIw4yYqaXjuUQppcaaolQkZRRhmdG7
1i0u1Wel44p+juPgV4yZTeZ0yEdZVgAncuDATVR8b5ddCI8IcHne4pu/emLYdYBafWMgqaZHOH/r
BbwkFV62IEM8dUn/qgTEkeXVxqj+P7yfzvh5laZuB8JGJVI71+SZLX9MzwHr+gbw11P1/N9IWwQL
v7n0T0AE4vjMz4OZQfUtfipvIrZ4MF8NDFvPFRomxtrokZm4mWskecVjHbusj3VX1VGEMWU/VWqE
rhFo1ZPqU2xyGkcb4AcUrW3x09Tk1qGynvD6baPdJ858QAVhow1tGFOJTFfgeUYoStNDTYoKw75f
XB6Cq4wa3fh01HK7otEUDYyOsCPitm1RlXuuSZ9SNIibBpxqUmbnAmKCjJiXt3J4wtkVJChLESTC
BSo9BwJQtM/gb0j0Sy88aaE2DpJ8EpaWMrhzXCeAr1axP1iZGRPOWUH7PvhoqCs68pM5OT/We7Ge
7x7QD0nWXsRG9a28zu9Li846GrepmOBDbE6PlGUtPxtaUGNm4dAXLW2W2dE6f3Oja9vNXLOjEeU6
gHtpAKolJ5skDTwov8gWn7j4lOzEfgZpOjT3VTcr/k1No07+SyL36yeOQXGxeuTETW5gK6jEvZSL
ZK/YHBfBM/0uD2JESrHv+fvarNgh2WzPuw4eX1v12KA1rM92HHAHipuLfrlWUd/4tcvJ8hEnIEHW
54JrFXCxWiqVofOv7wQcCvFiGZI7N5+Q+OmPnms0p74IbPbqAkNGrvRGmZRh03SIGxBvI3RxSfQj
Set7OcWF8QgWifI1pNoJlMNaIThPT4GU9LkJZiENEWkkcv4e/7eYLDInUruu9aU9Mgu5kqoGa2E6
hk9d5iy7wBA4Y78mc05K1ozcyTvuTsM/ybZPZAbUCY+Q0kBQ/e70DGQeEoqg2MlpNcqWDpl4MU+5
OZGGb59hOPF91r4jL08Bc2eYMe1TU1V+4uvj8eAi+FKD/yKhUm3zutxDHEunNzhDciahjnFAab26
5LoFLz7bHGfExQux7i0olvBX324cuNuCcVQ1LxbSJfkfUctnAS3SLsFUf9UwbDFmtgIg/ioybdJh
fzcqL9CFXVWgzuo+x26d2VI4FIB9fHKdVTIswxzc0XZ+7rCUt9G89R0Px7cvfpgb+50qsmZozcuH
FDAWVV2tjxJvxIusMWpFRTkswXQsVIk5GJOpsFpT4v1HyUtW0al1C909Hcu/Bl7q/1IHGVYWEYjV
CHabWKYY5xpSLqomg71TxGnShLJiPXSFs5uandh8M8j/jItmdj6qgZyXYrLcmDslwpEIxOPmGt5M
x1mPM5TWmQBRyRVU9iwzgj6HQVaAEqitZxKZ0vS03h4HmjfMFOMC9CgLgLw8/ZIg3S4ukz6hYtcq
+AQuK4+MUGNOlhdvVjV0Ned5ryiAunY7LigTJnZfkZ3pjBSLMG4h+U8J+U8R4W3tsMyxWsqTOSkP
AguaWY+imQoZQdAT8kaBzrlkGKcXDLKLDw4OAnfnhJ+CWVYbq3yYrrR+wjGj2bqKIXCgIrKyXAZq
ophndwOsiF6cYTnEhjqOL/b9RWzTmhJLO/okWF9Zc5N06pZ1fRGeSujx+3FL4WEPNe5M2iuXKXKQ
pBef1KQS1wnqks5oTgHOpG51j5zkIjF15F+LrKxj1/Frx8/6CgwRhRfa9okomtsAZZqgZ+ngoJyA
BHd43mgCKs0rwlB4eIpyWmc6Gw4KfbNpIN90VUliBetjKzwVdBHlR96dowPwjTCWD5Y5D6spf2XA
00uD530MtkGWPZZcMs9yMm9jn/EwkMBVZ1QhWEBeTgux+mvp/TgJj4IsRd38W6QgDS7ykcWUb1U9
ix6cWOXY7SiR8f9rn9DoaQjeghSHehAJyoG+WkCyI6HT4KAbLlnVJo6lOK6tTIxDWJ+ojoFk9M5i
3EaNg5TY34gTPNqSP+ttZ1L0Bn0behE81Zf6P2jbf2jJNtta+12ZjE0sXYHJBnY3S6PoP8HzpUL5
/iC9ja6gjgzgY+V6hEDviiq7BObElaRy341E4LBOsIxdhxm7j4WR/hfaG3zIPnO4wal6Fb98tvZS
VVmwnUejJt3+1J23OVPLgbv+XGbVkl/1lqdkTWFCnwapXiknW8Rz/395SWd0DksoyPWmoRhmUEbf
cX3ukQPnZqcS0AA/QNfcNV3eacfiV/tdWIZCN6hzR/8WecDJnGX2FJRmH7BzOLuhzr41YQxlrhZu
VJFGlMd2aVyZJwpcfqbkMcdGW4bBCJteIbXswmJe9EcV1P05w1KUPOYG3qAC3agM2KYn7+NfFV08
ylFmPCvoIElYRKpI+szLyORLOToW1S9RqVJ5RxD0nSq3wuYMDMri6kej4agBesSIKgT0CkfHLPiv
vyxWlh0JDLTRWpDwQ1QnNGgOjzQFVuHYMN5wlfYuYgVHoH/Hkki+iM/J+7UTHn5mF5L2jArrwOOU
yhVNggzkGpjyizTaXpe+1TlP86I8HSojDxE8f4xfzYcdoHR/YJ1aAti/PQmRMTKn1/TruknrNjms
29R8YzMxJLH1FLDFVIKdX1mPc6xLpDgUdKruZj18WaaHyk01f5K2zm1Piy2OoW1TbbYEW6yL6Spb
9Au/8qc15oM+QCTS5h6XUGc/mr7Gk7IsGCPrsYjv9LHqIHnIBiqDnCKfIiv8rdm8eecfJJHQkLZm
4fhjL/DyKG3lr00u1DKDWnwU00NxHd2bHCOW39jiVMGYLgGqGiY+ScG0CESHfcBJ8nvnUIfVa9NE
TiIMxQV8Rau0OVH8RqbkdG9jIv2Dbk1OUG1h9wmnGTQ/qM+iM8NMQA/UMErSBPo9cfb6FsbHkxsw
NSWf9yEc1h5ClzM8lCoFRluOTtNjCMjoALNNfni7AQFRVTPmQPpbWYyGfos4W1uzOKuF6/LgyUf3
w+rMv1MwCazFGmk0KdIiMW3JldObrs+LRlqzHj2W9T6JKPdcxz6H1Xf8rUVx/CvreyVJZpsOmAba
ab0t8EZHbu6lkpprKHBJm1b/2D0nsIU4dt+kUgQQcAs9uSnNuc9KuNhHsbiszqMFRM6ehYIzF4zv
MOPkjXg0cRtYgTMzoZWsF+Rbb6gFkxN5kI9ZmGbVH5Z+60P5CIimwmzjoyTQEKJDtJPbOwCIZWoY
S5rGo6GYP4/lk9QEZNOOh9zsXF99lXzma7SQRXn0qF2FWaVsaNlsSkqzml0cZAkSrRS1Rh/YvaoN
wRqQpOegUOT/9lKJc0LUXFgxyI02sgf6dkjGnilr6oizubIEO216Y8rbjf8oJhE28YUJnJmq6MJM
lEIcnKbNPvP+BNBgp+mG3k4pB9tPBfPBvgp1SNkfsrvWZZ47ZhUlU9xbYZSUiP26VQa3tss4z/sx
p2l5LzuEdA+snMDlLAfvK30Z6vq8BEUI9gn9MAIbwwip7V4hJ1qbvcJxB1fVdvLZhXORE2mjQQru
rMYfdZbGZS5Y6v6jX7fNzpySIOF18kKSFfhtur/Z7lKmaIqtwVL2BYDxU0GE0yYT0AQQmGuE4VJd
EZm1cOphbxe1mSognMwDvp8+51CR5J8s8OybSxXeifcCJbXO4OeqTnPEJyIjhRRjCYt+miCSN78Z
2BSqt6Cdb6YGzrf2St+iPWaU+u7n9d9pGJ9A41OJtOojfbjiIZkEOfjWS5pHqnL1nMppbu4wU6Am
1e9iNtxWILLVL3ZX9O1hqveijlyUsrtE5GoLKruJCuKQbMBsTX5O5l4PJo0PA2wwzFEIRj7Gt0r7
SuK20gveJn9pD+fg5dfvk3prqqPIMZB5rCLWHIh1crAjXWk6IYRZq7S4KCSJnqGx6Ir5xvCIXGz3
6N2PpSVUoiOl/7Q0FBbiOujjvZPphvv3o24S4FJ4iSF0rlZPIn62ONOnDkE3tZwtFwHSdSbRU/9N
S0CNpnuZJ5WH1SN6zYufLoZFa1ZbeIGQ9uf1UFVCwbkXlT1BdFqX4r3uFGf2FzCez4h9dGrbP6GD
9M//XRl2VouVcFCcWU32FOAPhnYyplEshFRaQcTQwjdgtYoaxQCEwejQMZUjBg7rQoARq0HO6xba
4CHQwvGQmSKjnZBB/zsUJd/uoYqEbzwbPGGjLPblIcbEzIPbDkBu8LOENkAUHI3SMhMGqMnM2Iih
4a/FuZB+xv5T56T/4gtW34zjKL7Xb4zqMP/NCAJTeKgS3slpHa9Y+z/CGOOVri1bs/cVo5S1YTww
HUTS+R3b/PFQQ0Z5M5NGKqhggwLEpIJZ4HpcBxaZL3rMJHvHqZTL4EsBGUSzPzHbYW1+sUsadNLg
c6IkNs5Tzzzpvqeojvv+RCohxpmBzcG244xGFu0grTrAKfxC/OVIfdneF4L8lqX7+qvGWGmbL8Pn
UO5u2UBZKmSV0Gj9iqs9oEuKnisbT2jj9DjONYFwhsdbdJiqM2LUgx7swgtgQa3I4DRV4mGu7H+J
Y6y2LI1I2wxUR3ekE1oStBJbKV0Eu2Wjcoo4Af2yfKj0D1g6r12pLTmbydMXyiyGZsk6kgSD99Ek
aJKVdzKIrVp+F9qMN5FBKjipBU60qjH1yZ67ksJ3sdWbtYF4qcxxiev7GxaCirahCV72Uhn0m5Zm
5cnmUjf0EpG9gLsqmUN1CWo3Bavtb8Bc3UTL+eG8CwI4UZ8bzcWuWjhzhMEKjXag8+fb6kUJBdgn
N4WEMPD3XxoyA7B+onEf50LsJwVKmCy6TNIbaLpmGQm7UQ/ADDm+8GmkQWjuOGAxBvspRnmzK4Lx
4z3XGYmhiwSG7yMXjb67cEHUlPD2FsJ2r6Op+G0hX0ab1+UjMl4LUtgDgI+6jNHsImT+YdeyNzfv
ejlXubyvxpqVZQ8+VEELruQQnUm4OD7Fm1MoKNAo39Z9mwQUDgZ64SFNouiNo1ifmK9x639+ehnD
7IHGvmG3JL4kWos8CO3pNmyeZVzsovKFQKggrO9j4uHFWH6QZ8QblG7vd6CTxhzUUFS+pF83rT+M
7d9yT2+WKrCxYWzk46XyaQdxxfVxHfrgURnnscr7t/Vj03u5R8zwYRLAbGfYwZ7pCDOVOYM3fKaY
KPC9vccCkOWCL2ltf/jSWL1s0TtfoOMGkBZYqyBy5pf5XhuyHTmuPW2nuaOQPuwSGeiToCnsS99Y
JItjK4OpcOEUb2WCS4K/KvOA/9oTKFOb+P3Wv2enDvcRAS6+u5sSTs8nkEW4PeyUW90d9M7ONw2D
NXt4rq+AIfjBWJ+WDzjtlf63nbesi075Drk0IuUoDck3Qo/dbn3NKyWH0PfouBhFWuHf2h3YlE4k
cGt4BTnlP4CdLVPvjqHX932XeCEXKVfXG9OuCIgRujrXCIh5gM3nxPa3u1EhsZfyKQua4GpSDnsK
pvsiGzY7HBzeU7WYEfdW1yXmexS227f8h7P76pIQ3LSWwjxG6vGQd2I2HCFLXsUAbBfkdiQ3Mwcq
QfE/nO9XSDpKPntf47xgwTnTHxDYK1lnI6nYI1GyXqW6kirLptPI6MQTmAjhtEnv6SNmP0oFnffP
Rq3HkkyaDlFTR2C4rvpY3GVsdKtBqIHON3pbY3zuXIzJwCLmmHKt8gTKvlGZbrZXZO/Gj5hOucSQ
Iq2XBxIjS0DRwTlc+XnfYcc/SLIBvsfmAYf0/hdSWPvZO4kfxRMvOKYWaf9GqMpP+w0T+m7qJlOV
X2dwruJL91gBq1JPmx0vTNMrGHaUmtmfHw01+OFJJOLnT30ErWJf2pMhqZNWhKvBrBaw22oJ/I0V
wlZAF7bGz2EvWiTOrMBpVxt7/cyv5bdsG7WdphCR2ysnycGoY7/sDE8Pjv+LF9enbToeTKJlLjnJ
IlZFzXNueylWF+dXf87/TbH6pK4m9ZIgVBGRYm7fNW1TkNmnFKC7rcZoVbq8A1VJmESZm0jDbxgi
JQVqo1nRbduUEPpmpg4Fi3cnQLlpV9lzrYc961Wb17fccMTT7APwCIGi7R9YdbNfuqjtwtWXqfdU
J+EDDASGhOgbKVWasyAGgioKLnrqAbGZ6W6YnYWVyd/mgCtM6/SGafVDhnpV/nBcdxiejS8bRHdD
lzdu6GI+FJE6NyTc9fKlI/laWtT0ZDDcVajPzH9x9tDgWE8izT/J4fNhxureUIZiIKRYBzvmr1+Q
g9kkZ2mfTiIlb3W7VihFHJxw46JOTMGbIB3Po+1N3W7KBPg/FBS2HlvuErDSJZ/sOA8eRO/kfK6a
+RGwKC/cka5lExW737hoQVhPIsXeu3pdgO6rERLkBpBpga8I1a8EfxNcLvBKqVlYCD6o28/p4a0R
iiJlUT8xDS7UPkXkwUIr+SivGBqQ4KnZTF3lk9VQVCWRh6qEISde0ofQie3vTA/3C3OkiM8GULE+
BDNzJqHrdVyEJI7jZMaMrR1nnJp41mxkZLTsvz+diTneD1nvEX7SBEq1GmFxEzS/0zdp6Je8tPvj
oT2QGsqTjrQbFySczUjZiSXll6rH0tATLCRsL5DAOS5y09CJl+gMDdqJaJGpno4BKVsu59XGrHRE
mzC52oIr8MJ8AjjKU2/E1wvpvGKrpbfds5+rc2lld2Bi+2A4cvgK6S+MFbaUzYrI1esewchC0eoe
DBoUTXhbEj5oOfgcFfmex+h7v9txHGFvofmW852CUUMw9mkTPk2KR4tSGhHD7wL8SqkLOjC1QpN+
ZMsn/gG4Di+f9liTPYnGK3yw77DT+p/g3MZJatZ0IU0by5zO7l6GIfM4zVArY8eLa1U6lNxSxK3x
W2WkaLfkY+AuTyAUC8RF06Nr5EZidS75NZTi7LrVZgyhteoxyswtqHQtcngwbDukDlj5pQUT5Db5
ABwuw3/gko2DnkB8D/jAe02XunSQVAHXYY1fXSaJnAke+kZMXDZt7pnch2ZGVy4sXhtpbcih00fT
x7pKe0YO6bBfyc4T8mdX2zP87Q6TVmMHw+hYXzRNxpEOjjcdct2AtTVOcZigNMipfpG5fCjehgWQ
qGiIKgMh7gV5uxZR2Q6ICyEAr9gcxJIFmz7GIGc6w/BlIEOTo1S8wx7oSu2JRzFPFofoBZkeU+eW
nWpaGIl+iaLO2+IL+h5gMD88NbM4RO0G5f9KGFKX5AhIxBQBjd4NF0bFuiRfHX79IpyJNX+AU6z1
YnsCnCURrq+cJbI6VV472tmt77rfNwlKuYz94zDVpAV4kDyAcGcTZ/+hjdvE+XL+FuF/pbtMbuY8
Zf2cOPztcRFuyy96fnKgwN8v3Xw7PEjAcKLJPDihYk6R3qZA16uSEpDM/eBzQXYqadSgAayqMusu
a4NpwEZnEJo1QeqQuN4RCeOHqDPtIuQwvC/3kvsxYmDxh6aHx75en5pr/vleqBU8HeSucbLht1hf
Bl8s/PCsSQjLUike3jJ5vITvE4fGKakRI4kHcFpgb1m9lIyXMMUSHlDvVyZy3wobVBe6woRrPQ2H
U01C5vnLgVwwfmwUftLOvwBWKU9R9rsg22ya/89TwsUX77U+IMp3DjbaFjdzOUWKb+qQ/kUoffwH
WiiyPhnAdb1FmwWGFQVfu0EWQtWNwr8LU2RhK3YSLHbSQ+5ba1+iPRbPxE1/mHOrNTFZNiX8QJPh
KbWXC8Im7ctr7VWdYyQ0SU34AsiMbROYJoc+L+q/1AvQp7E5EbNLBQTuRXrYQ1QB8Duv5Cz5wOVO
zYb4lCU5u3K9Ixm8F6S1azsUnY2Q6CEPbOvQQv2pV01BnL/q+FYD65VfXe+kYmfjwORaAs5MQPpW
4+XbpCszhFwGQio9J6MwfJ/P0ySUhj56Jymfk1ttN5ET+o9LgqHZyVY54RxuDXcxLfzdxgDZ32WY
5gNWhIrIZj9vwhJ9pDTOBcuJPRFsPU+pxc3XlObUH1XTij4nI6IQ7l7V/C/K1HFINFKCFkI1c0q5
FJDyKriebmBy/zGPcOBsKw7U0vXH+sBkZxEIKmTvmzM34UKuP89hCipuupcoDBW44WXyGPY7mBnz
sx4pypwobTUMxnkzZyCmT/sUa/taMQiBAjaM7zY5zTf8BL94fwm9fgj+7PCouFbMrevM3NPuzqSa
UL5mZbqX2YywFi3zADJG+eRNw/zr24yGrd4MS7sHqZV7gMvFYnN8rXiuKokbWGiSSfieUae8Q7Mb
qbBQsofUNXUqfWgG1crgPneNoUWjr27J6URXalQSO4uTP/17vJMMmObUVwnyIFisKBbqi1lhNy6H
KWloliMU/76EDkgZ2eJWuz+ZPlEeZJMJZ4zsXeEc1kkHBQhxSYeIYowg2Qipu1bpTpmzM8eXfSvC
GaMyz8kPFzaHyBEqaWbyZ7uW69qc0XizPV0zEbsFaDIl6sbHU+gqr/401gpSsFS/jXYndI4Ll9l0
fdtM+xSiA4/ut1qlOvGsMyZXTKRoMUT4sdTpbWlvct7ilxTwumSnoQ+2qdegMULh7ojNO4UYcC/S
LACFbz4UYl7a764ttDTeOnOS62jeb0eI6MEM4c2ynIG7uvRfs71BGtsTOgApGLYcFedog+kF6gDM
KMbm0IhFlUsiG/HR0n1F5vGhr0XMR9S24qrBafbdPvaKXRHc8pxlenKAvvns32k7cgeD68cN97pm
YrXEqLmdjxGkTcgW3I8JKjJruXYOwhuE6AaK4rjfGSy3w/juejC3MgxtNvfbxI1rxaSfxpRVOZa3
m32ImV9TWNtQ68IEdeTEmTBcE0K0+lj2lkEBVJ441r5uQSTgx97XK0BnMTxXOacjWqZMFifgeo/W
qQ9lN2PEj50CU0c1FKgtkwViGj0S1STsFDHjltjgLpDdlUs6qBtb3Dw8tvkp0wwWfpcPgoUfuX72
t0eRXGosSd+5+UFRtNDmUlwTHhYHfvHV9yazhzD5VAAuBgc44tPIa652J5QK/+tx7ykgBK+GOu6H
KZCXL8/9F/3f44liHfEDlDUfT3RXbfzYuUckM2F2HDiowRcFupLDtDLpCJBHw1pYlalYF2tVUOmW
scpTtJ2/t8ZbVPctRXhGMf/oCItJLr9ODyE0KnmAKEfLql0+6FlPdcesW94N9+TYEFNcFXnzgt74
DSG4NgrDZZjWq5D1eAtwQzIG0QE+lx+dmU1rZzSwP7Jcbawf9lrAKeO+Wldk5ya6KsChVXLIcKPP
qpUusy4VisOQs41GzOX/rGPWNRFFemaXis2dRGt7NowpiYL8Iz2iGdodPkFhijEB6kcsgFrKVFu9
lGdKsWUhr+c6WL1P65LnwIMWO//oWMPYJWF7nkVMns20mR/3SbH7oMB+BTn6iaVnNlaeZ+mZ/jBg
9aaEljH5Bpt/R2gPJbgREp8l1SUO3c7k0dvUHiEjg4FneKaOSE+XdZgw+fxEuDBJw+8FTg7aAIPR
FOfSD6jc+KCxf9MwP2VIhHw0xjQE7dE05LshDC19vxZSHTVSnn+67JiF7zEiEQEoyFCE4gtAuugh
tgKPwtNmIAjH5PhbkbtMZ+o1IbXX463vtmCrXUoiZiVAK6SKbdIGrVyEO+fjyVpgQIasPj9uQ2BF
qUbzAnnstukNpked4yUkgk45FKPU3iwwuxX9JB94ePRXXNKq1EaEBfgCdvYNOKPvAYYt6DYZDr5H
pmd6S05igm65JnGMptLhqS/hg+ZDCVRjUoOBlxflHOJnmisQMEnTwpybdRUhFYdzGorEHuIWkJ0Y
I0bOdxdmdWRmBTwelEdE3PotQyMZb2iiOur54253CjaeoMRprJbk3SquWOwH9nuCm2WcSmezLJL1
5Q2wENHm9VJlvVSpMt9bMCobee1F3ET6QS0txT1XeLg7H5j5KIHAHUmplXihFixfprADqtY5qdaQ
/rxT/+ygncMHhCG1eJzBxEdIRGCqvKtK5eU+xk81az1MT4Tc0a6fZS+X0xb1o01IHrNHL7GmFBeC
Uo8gYa1AHZKMzHX+74NG1WImGxjioad818FIjO6bFQzTTeMLeG+Q3IRjeRZ3cuMIZ5POOL9ND4lb
V07bMhIWUT/oLPx1O5i3kHSSVEVVTybJrdB2qjA/MQrC1pV3v0JGkBu841dIPpZGNyAveqX8AOG9
7V69MmhqapH8ndZPCNiDz9UMT7FL47IvfMCHWhxH8vllCWkJ/Cde6tqGGNORKr3ub0RmYTzDpUVI
VNsAMmcd2O+DY6lGUzKE+U8Wq6mxDz+p94GX+UUC9i62bpmHC3AnLCARVobaInFrNCsU/xcs9aDz
6FNFeYksln36anGeadyYxA3ActHaNLTUdBX4T6GidZjcLwFoN7O9vXNwcIvF7GZIgZN4mPw5tYq7
AeaaEfs3lyTW7xeZPpU2SDYNKudtZe4cF83gE2ildWV7HDv+NdHfh/dwCZYdDFpalKF4TjVzfGFF
N9ixlJ1No3jido40dpqkY9/Fb/iTsWtUZL9CXhT3Q0axHhkaZ50IyKzGreJtBw6OBisyMxchtOvQ
PRZmZN7FqUFqEIuXF/46xoC25tklXiw4unOrNpt+8CHK0Xk4BF2ZxHdSFrwVnGMHx1+iLz+qtATg
aQUArPS43hcmcnW0V49PBRfTwryfqtuiWRMEF+qZjxN/t4ilqJc2PFoxngnLBEgUyQCOccRzOJZY
eTgaQQJ4NjqrE5NKxbC3p62IR41vWg5PukPKjTRdSTzKbtclGmmhuJSAGTT4xL1VlUw4W3bgEtFX
iyXd1Jnlvw5uQ/zH/nd9P+R2S88SI2pUUmaMbwiheDEH5ufY1s6oms7vR7E5j+u+0G+Fo9oGq6kR
wI7k1mW23di0TtPuROGcnjaJlOZM8pPtohgF8QNca/CiP3QIqwb0I0fhCXhFmS57p2X3yTXBpyay
ZNZJ7LegyQ+vxuUHAncAJXOjZyHhWB69gsc762N9nDYzqIOr332NFX+CKYbid9cFgMlhv1xieucA
rfyQDpK90JnZxiYVzCD+fAqbFqYmyLY301tONRhqI/fF8/ps3XkGqlh0XCFXgiIuBlMI9ulG9iWH
vHfrgxWBdgLW21RTMjdGE09g7FRZQxzs8TIfYr8dq08KqtmRrcqNgeGynANzVbGVINoQoHNZka7Q
gafKmgjgNdl+MIIGuooV1oSXMMCnY6XK0gvLGn5DjYQoP+TKwEdJiofkC2xzb1LrnkIQr7ZITj5F
Zbv+RXrX7ILY1YsdWmqNmxsMG+bp9DSCQFAe5WGLXOCex8Fzyz8Rz9/PaaBiJg6SlkQ39CYYZJ0o
wVmvMkp213BxbdTR2W4mxiFN5Q+4sBSaGbilh+M2VKZZYXuR2pOvXNPrUc/rd4b56tf5P92lFgOn
hFyPetzIIu/3NK0pEVSFJL9i+caWmrEZxxj880XHa2JUhFHhkQEb7Ti6b7MPOo26eREJ7rycbIOJ
CVGiCYSxw5CcV4HdCfk05qO8MrcevAVBbIx7ARbZh2a/ISNmqpQ0rX8u5oh/evSCMlUlhhF9HYpN
15Bwum5/6hdXZoCXwrCmVBwBub3JoCMfalDgpo9w+71a231ochrHPJmxR32dR+x6UkKN9Yl53gg4
os2/G9H8Eu1P5h0RLRIIsCTx52LemTn/ovfR2kWzBh0IxobQ8lYXD+bu0XVQlROYgl8PnXq4HeP+
haXqdXoshunqB29ACbIH13No3lZG/PG1lvwadPFd6LcqerRnyzNJav/iVSBtFEW4ucw2TLGAnlM4
VzEb5IHAdL/RlaUwOtPeJySm9xjzJwbaOgr0CsKAGHsJ8Ld1qouQXlFxlasxKTB3ktdoHKd8kGnL
mzxcSOe33+hGCWG7CseYFLmg8aniwVjh2yqAK2R6MyT9tUiKiWDDavfkuK82nQVRHfl/jYsXDDi0
sMEVa1iAwrqJ3QvGwTZhCGHfxEUhpqpfJkmp6+7jDIptgFUzKSV/fGcDmI56WbWX8KmRSRvaLCKD
QSp9cGbFJU52sSQlKkytrE5cKraE93V3CMLoHjl7LFKNJZDQdjkAgEQl3Gr5lH8x5l9Cvx/Ld7xj
JpruAaYMXdOiKpWBseOeABHBr2hCit6XuNwSOIPxhFH6ygkPHZSiOIAblADBfzU1oQ1/d1vLMYhS
oTM3OFvX0sJxRFs/wyUMk/j6tbWn6TK/V5k5jLBdDaF6R6ka71ezzGJLv3ttMMD00Dm1R3BfODTg
kni9q43G3WKKYBbnh5ZD5mcTPlKjyv+yCJwWFDAO3+pKkykcHQ9mTeYrPoOPyUxYWgRU1XRfw1sz
uB3+W9EdHZ0192l3dLdo657LPtObJ4dBs+pTLpdEkNf9GX2oliB+br40aMYE1jzafEx4f6V9nnVG
aOX+db3NcBdDLLzCT/+c7XZlOD3qdyqNLAQTka3Sqo8utscqSZ1f2XcbwjY0BMS0AaleQ795GTmB
Zk0Gvz15mkxfEyXg2hnGymg2eaXjPhLGB6s77K6+1MQ7vFXqiLORzxU1RLdbe8lJFkAlTHMckkoj
1zO8suwF+BcJffP1z7J04yfgNRUPl6iitTIG6yzxOago6DTt3ykqvmBv6nIwEcfJz6caGLduoc8O
G9rlSjc3hlJ4wTYKq22hMhYBZmWrZRjcnlALdAEWjREer+E94oYNVmt6HT5GRZWOssiZjfsUr/Xx
96kB0BuaEd8cfbWvaZVcPBt/xL9r8F7ozXdMr1f5StOXlB7/x5TJMA7tghzU9LPHT+XGYGaW4PeD
IsiigqcAh8ZuvULgHO0BEL0LBXrTyDEQt2GI1HF40Y/yGM4IvHSh4S3MqwbYOwCv5fBP9Lqj/wkt
7uPNJVUVIGdW3/Aux+6bNEBt4u06hoTN4NnAZRJlKO7tXWzEgKn+Exx64aLzerhXH+EWa0MQXdE9
XavkyHeZ+xIkwsj9+S14n4gkkpFDo8Coc/tn6NBlMxYw8IJb61ybXVEOp3pUrjI6NnEQ3Lzoe0n3
lb5P4DG0zwoC/YPl0P3AcaqO+mYvQ7TMmj0Lbe0INCLxQbS3MaQkt2A+Yvw0NEkeFSq42OpTn18k
RFPqxHr7K9ZndV+JsFcsF/ir6MIdrQm5bIZYg6Xh3BV6No74I4vK4HHTYH8w8pz9EqM0QIDiKUGx
xyxq80ayMhil+P+A3KVieIJV1AytMWuJdnzMi5riqIKgj51i4jVokWCYjUSGu7n6jRulhTtoslwR
3zJ741nun1/IDvbBuLfqdgQqJCxv4uZcFJNoRUFN1zCuNnLTWcHRmK7tskurN02lT0X7O7oAQhcJ
B9hl5ti7vJG3h3sl/jA+n0ksR+QwKtJ3SLQAqWxGGMPHe3SP5N55irYl2QyGIcKENgLDZnXWdhoU
kJFhvi6JFRnpcBmhE94bEoPsJfQYu9UCUHbLhE/qfF9vYAwoE1NJAqavGJ/Id33E2I1iZ6RKBYSY
/Hkjdjz1G5RXuT46J207z+pHIRTBjmjbmOQ7pTHAqsAwzlkV+weef3C3Ikr2nbcNEJIp5szeyJA1
+0K9w2Ay9HX0ImaE+ThR/CdVQt6hZnQSDZN8aCqbo2PvXlfL8gRw90Q7FsJSNf567Vtkxs20KvnQ
46c68z/OcvJ6lM/e24D5MMtwBXVzwVLi0kXgfyaAg9BBBFDtx+m7H40E1itMHNebduTn+PckkcbB
K+DPd48H15qQSUNpNssDt9PBevfTt33HJ0ZJ1vLuI52Kwz3igcec8JwfpLegBGBs8o4pUNwCutul
nP0FttXEjh0TwgistXm5uyO1JyHOEhkDUMZslmDI0BMUGQvk43SyY5D9AhemCzCZgG9DZf5DhCpo
VZ6x9kaxL0tpVxbjVBBBcLo+kqK1qjjC3KpbUQjRg+1mZSOIwIuHaYKIvORhZhZ9dBuuKEGZfyi8
2Ktv1XJXrfWUd69gDGh4ARk/gWXdDVcLkWb0GiscfrlXsUObIzwhTp9yOOSz59giRs2OqdZl1Afe
I5CE0NVWtuOkd1BefkfvzRomvas1Jx6Ow7DoSru6kZqkl6mKiwrxdSBFFbNqhuwH1KP6QW7mTEDh
ns2NRWEotaRPgZBsDLCLNWdijOZ9+u0vpvoddmJcicbGpfyaLQlFkx0u5vWD3qzjH7hjBZLrVAHs
YogN6V04Swt1dUSUSb+LP38Q4TT+5Ln3VQauzugagF2+9bbZAqNBpzh6BFq05zJQi2efgswUrKCx
9jhfJO84yyGXzV8tPZtuTJNkUL/of3BzEJ8MSlWXc7Fe5/h9may5llccBiMZKPexNPL19kJ4xT0Y
SGq5Glo74w9F1vORloUK78slI2yDCG5RILKqqq2Q8bO0xL2MOsl2LTCxlidZWbYEiSFdzYwgobE2
G53Shahm0MdF8LaboXnSqyr1jRkzGc3/MeHT8J3EFBdQQpwLb1EZQT+ZwRl8l1cFp8TUwyAQN9A6
uf0ldsX4LGiZratrlI/tJ1G6rvuQwKkhqUp/DM9hIxyKKT1JJYLXwsPz9WERyhxxcARNdZ4Jaz/d
sa+wbYPausfZ4CWd9U2u5/Lp+2NIVtjbqGKoBCRzyEloWp3JkqLe6TbPbN+AeNDdCs5FtaPxFVWU
dHglEtSx1QJtGZ1QstuB+yoSKn/TzIxWnXrYjZSXAIDWGeEENZV9LrNi4bq6C1puYXltlMKfRqTf
DXdptvyt+q0gHZ1bRhwndXc5P9Hb9W86y8dXJ4KHs7jTALLTlxW5zQAfwLNAsRn13Mc03cLHoEoD
FWa/ETTTtk1yjQ7Oqt9FK4Khu0XmZMxPkOopnv5uiImtdQBrQ27vJUIZB0tXR8pZrOAnZVYmxzYj
hci4CJNUicdHzXExu3OGt0Pm0oEdK8sa9uplbzB8fZChlLzBiw01b0OdX++ODKnt155t67gId31C
OSVjRe2watollOlovSnVoJVdgmNfEmjnesfT7zrodT51ySn+uqgvmdNQmKw67swPAEBe+XNw2Ae7
/rAXX8+WxZS80H1ruxPI0gFykTKTffJgYNcLMJqZzx0Ps96wLWtjToa/toj0lthoeQOiaD133kqQ
zSJ/DxYlOr+KMzvw8iTM2IsIi8ByAnWvJY/AVy3+84sxdL0OqsfKBZLxzrN2McFSuN5RHRcTR6jH
07Tm65bM3rPlaeAvO/NuILbljb8gbceNrnWVKJeYt6FUm3hZr0u+Asc3lnggpUWGHStA2QkxymyS
RLoUF+caUEYIv2Z8WXm7ncFPI0VvnxbKvGRNfHjUeaVajpFpc+wNucspTdIyrWgUWcmqzVhdX3PO
K1ehlIPb3fkU+/kf4i0AhK0DrSEt8RPuiin05an2W9Dx6DCnFHI7fvG0JYKdz+qGGXaucUDG6aU6
3fQ7cZ+bKc/R3n80bAaW0q/JYxMXx9VYrWggLLonrs/n2cnmSupFjhW6rDAoU+wyeg9OXC72NPz7
FRgoqjwQNZHp8Or1iZpgSV3NwHsj3xVdwJmRn3ku0OjUCHBONAOUFUMPG7vnkWPDFiYIL7sVBPmb
hTTl5INeZqRT7NBJeAGqFc0ZNaj73ECPyQwoOeNGk/0/dMk8yeE8TDM+7/xqMm0cRTn2dvLkhdS7
2o6rminab7IMFSiqn0apySx0VpqpNDaLedjm1NVgURu5/F+V0T2sGHUnzS/Qt3FhQYqpSYEIdYvb
/EiNsWbg/gmX8Js63ZSSFEFtodWdOsOR3D1tOs2mSGzzkhNIGwF+k24L9QFF5ffGo71J2pJoQ8hz
vXxOCm28ck+x1wieMNDJntMkY4na1LIAMo4pElrGYzZWitpzHtUqiWLi3hjarFCwVp7cpBzt09oa
ZDm+IGyAc3/aEImAgSfYonRVWWa9ZAkLTeW6Bl7dT9k4mb858oRSYSemPKCslX6R27SKEfWiBw2j
eUIQxi33RMpm9c2r6AHPgYHqB3NVGKnHr+bduxx/MdPfZpQqv/Xr16SEVkcNseWG0/E7amWHx2xq
iuLSa0O57PjyavA43SCXAskL+Y5YUQqvAv3F/U+fBHSYLErwTWkKeq0bJd8qgmswIIKJg9n7QMPr
4ItxvToPGsl++m8ZRMdp9icc8nxsNKJo7o1ItxokyS0Zr2E5jTI1KkbBXPYWiURS+5+T9bAwdHE3
LB0YLDJvwIq7WUX7fevmQ3NFvTwCxSiXKMgJQv9zIA/Vy/g31bZSWGTvvP3Yvc3KUz1IfIH+WZ2l
us0DvKLKb2VWbrOXrwti171HEOk6BKN6i8kp4Yyejh69uFRJtPtA9Xg2D42Db+1r7ZVQ84v/zmfD
Qgi+p43PcAGF2hyUVdv5a18VqTFyTxQkl0xZdWFaQh7PiI1IDDzi/WN/p+kZaK9ysrorr53xlhtQ
SFHq+XjUFqydDT4DO3DHBC9zOhWi8b81ixzlvucTruRiilVPO96s5hk4stHMEJFLPCxLwj8jdK1u
J4+3OzbuXTXE6KRrvG3PSHL151hPkxuMr+PJiwEh8/UIBaFYmDXzFz2jOPwtqoIQvehiJMpGB+bl
1RJ1O13zQKTiL7Y2NuuTwdVoNtUApPKKBPLRnk7UxF2rJQQObYpg2kbdCmiczNmZrSAh+oq02ZuH
FMdsh6+E8NKQT3tsUKNA7wdaJc6s26RO0v1/9R2z4HJtldFEjO19ej6+5OHp7xSZhR+hgikLGtLy
qXU9x5AaoGaTsrUa1LBiTZCshSX+2dsFwPi92wpU/SSWWRsJxJLWeY8x7W/vO5+C34JzIxjwiSOs
1kvb9Qkvzj+6iB08577qAjZz6RI2hhcz78C4LjOJA6r/+fYY+6uIboDJYkMhjSlIR8cI6JCyvxem
jlcSnIqRLN94KpvlSsIAaUIJ8/46QvvW2MvTIotNJfg5LypDVS8jBIlOkw2NS2PTR1actIeEM5QX
Vz7TEu2vvRqal5gqQ205cVovUh1E+zA0oM0uc9M1nY24VNu2D2eDu/sQVMDoyY8+RsHYcag66o8L
/nlSvKpV3tuBDVlkr3zsNfxUvfY5+W0rkqYwWmFsu9J/gVeti/likol2IcoGuv+J+b8beJ245nmB
k2aqxN/ZgIVbr5u4fwGXd8Y6DXmyBloIaW36hV1SF8Q1SckCvfXhjinyIUuCvWgTGvkxWM0zs2dL
00MetuZgoFvgTsYriVVRksVXb+hXs4Fi3MlDReHtL1w2SzHvD9NCDZgAA7Mf2wQb9IFbsAGb3dw6
EQvomUCtlx5yyhbxbgcayasqEO067CM6w2IA6/emPjkcgTG0ouiI4Yag1b3Utu60yRBUb88Hxbr1
ogecLtEwLIGyN/T38LlYJ6grxOLq9QqL0Ll9PrTj7MSAN/ms521JfHlnBJb4m8FtskZo12KNVPdL
WLQTy7EG+izBeb5qyw8/mUh/x/yM3fjndDho4Td/4M7S8HOW7yikAsv8BBcXIrjmbZlm6e3/1n7G
tEeNcAyYKDyQkoVqCLmYf6N1qrZwaPltt9rj7oW72lVTYT4w0uHuuEQmvj3iENLa1C8Ept66x4pn
T/gjFGcOK50xt9s9RqaIWr59gT/Q4xaL9F8Yx9sXkye78pzyNApfOXVVxJIrNbJ7Gm120nMwTybI
JXOYtLaCdlfAgO2/ia+dut2p+mrgdayA8RFnVCF+h75jGBYfpTbMtU60G0IH/A9+y+1LxcF3hCC0
j9XBaAI27dPdGc8d/2/B2Z2WHHsbI1zQ1IvoV2qOUN6ntZ3GJ3r4Sl2IzHLeQR6BFhB1JO6Ane1N
oy2FNsSVTu+MQmtyetwrId6K7+j35L54FkiK12mdvTpZM4M2vU6Un06wjo9NkkyGDYeLUh+sKGqb
/gbCsuo4Wu0R/8El2cRfiCTHBJDttKqMo1q43dazJxpZTyyrjZ9TmNEv82nAomSmKjGk3N7x++KT
9wOl4pe22wsf62KBjuguA+J4ioiyBJMvzIs2q5lO1qIVCM7D/UQ4aaKGqaFFFWvaugf8X3Q7s7Ao
Z2jRQJ4CGIll7OghEObhFmq9OmtCpIfSzUfNvNhAaJrER2f+PVbv4D7LI34EnwlSDENXAOQj6Dvr
uRDK3cekEX27Vww9lcEVKlIBUueVOV9D04PKtDBXJ5EsMzVWBzMPA8tjD5rP5Lsg/03gqkZzi6jL
/Fp7EimrPV+9VKFT3nQT8ohJMQTOM4xnKq12yr0+mKHjMwV6VFW9aCs7D5UsgAy94fiaENkI/QdM
E0vYnzrkb8wujylcS1GPYOXHzFM0dom3iRvk9jIGj484jcegAZr+yyyIxrGbAQAYolknVaI+Bt5R
DF82PbCCpOqql+hK1WaUNESjm2tL7I19FpNeyasGLb0JZuPIJ5dVB6VC87t+waUoBQIXIaoLXczI
LcOAZ2zFRzyqQlkDBzmjStvjmQGoNYyUHmUewoe9HuanafMZ2rilCLTYomAtDsU1WW8nTxVToUIy
Loy+NGmcWxx5o0DXU5GdU8Q7p7ygg1rVnTcQA2+6SJDzoK6By7pKPmpgyXXXbJ6VbsngcAGZDtoz
5CKb52cnLErHYstctGoL38yWzAh/dH2265po3wWhxmq67pzvO5MlQccKOtUmoHrNfyiydKeWkew9
X86jvbt9gQXwI4z5dsr5bt2VJ2suTTFsHFvcOb4oXnZH2OcVfyI2SXLBx5ouKOe/dBvXaiYVomta
FkDHhvuy8va3qH1pdlDjXPd1XLWX+C4f1nPRk8bBCRR214+5ml9GgyU0dyqEreGGcT8BaCM9AZP6
HqhBlGFPeKVk50XRe2N8qLFtnd4jcC770+uee96kfW+G8NvW4CGKMPtofW3ZUWPWjBNnISMPE7NO
8wdnPMxvRiku9rNLDavIdlf5D62e7tnOX6qXj5KipKOT+nXOCVcKoT6Olqiq8txLluFnKLe23tob
dgQI/s2Y0D8xC1+tvBb+uIXd3aihTy9UmhiroW43t9EUgwptz3SIPwBbPZDI+mpTG0kk2JPh01+E
A+ESIGek0dvLq8ID/S2/2ZdWPWDR2BC/OQp6sgUyVmRTdcbx/M9EUbw9LPFYQNd97KXnRQkGdrkH
Y1wzmQ9IKOMF64aEDbfulBFZL1QXcWR987r84b67snjblMj5johWOXCnOLLyBDh7iH8/l6pPRhqS
/eAfXLIADrHXfywVzD1EHqyepWODOTPJWJRbc4fThSUJ40Hc1Ao0Swh76lpVVljGmZkplrpaqXbe
nvNhfecIGDXO+4/4QGGWme7YYYYfvNtWnNveZf962A4+GWsXWXUZ0+bk1EvCiyefK1R0uXYT941B
ciOH7yhPMStxstdR48Vomy8+hbxxySruLDp1keWrv7N+1rkER8hZnzQ5EtdueQ+eqTzGbHire4vk
r+HkvwpkM1qDTJWiXhO58uXvdK16pEkIEekJHUMgXu9W9y6WnpwONkNogl26q4xJ9k3KbVhZuWgS
spaOXqWrbu7EyxvEg/raNxC8QUuOrDosMv3SnLSpDWdQ7WYt+YTvpIAHKT0RzxJWItYQdxZNtGHu
PpxHH9Lp8O3yx4aknTnXEEjw4xUlcs2TkiQvZi+9d0ZCiALwDJG7MLWELEEeWuh3tLDWfWtOITd9
N/fFES3p/y7694DpN7cR25m1MBbinu40MXkS3ZR4J/Cc8QQ8RTIk/MU6Tjf2Ds2kAvpBQ5X2Ml2M
M4+Oxj7yHddKldYPUdqxLm4mJnYql92sfCsy0a4LKfJpIU4g4Q8CHE9jbO7PAvZGLnZuHGH+5muL
N5oDLWejxNIIzceDlnQUJJW6/AUJMObLwNdANLs0j8FQDancwuPVfITfnu7E3gGJ4+q0kLtwgSAG
Q/TQ9fEkCb7W/TXAi04WyQBy/B2J3x7Ovsh7Omuicg2Ad2m5na6kqH42x40KVSk6wpu1pxOK9HBi
6y+H5F7scFrmH+2dNQ5AVKSVctQYLy9MfFwFlaJY0FBhLe7TH6RGWpjiimXWa8fuGQcDcjG5ZCC/
3RCCmMEyB9gDYHhAIl5jh01Z+gwIVyzkR+pcg6qXfzfxdQJUtJY+Ln8rQCjLWpQaraU0lye82u7x
OU6NyLrdI1lHoA3nxIa1PpJAjCVMBX+H+qy/2yYnFbuEvpvECzL2ZiCJI0Rj9n3TNx6EKEEd+tqg
p0qQagVmDxR7PycApa+wEAZzbW4JVhjnYVYhojw5sRu4VGd43SrO/vNFAArtr49UZp6bNgmZbtJ4
8oJy3qkftARjPXuhSmOMUQ99s4GCOEa+KS6CXRWQbtkKyt0Io8kGkZnn5MrD4VsfygBGc3ju6WDA
u9Z4Zd0qScC8cBWJbaKXf4Dwt9BZIjn4xOxOO6w/iQkY29SptcrspnYct6La6J7Vf+hljAe4dVeq
d0il7BK58wXZcb/BrqPMO0nz7ipht6RxnAkTGa3IO1Jz9XM955foJzKGyrYPDZ3ogINGv9LoJ/eL
/4UGXL60XYaVjKDb4kEwNRjbkGrVaqB/vq0fryyRA20KgGXOlyInVc7bsr5QX5eV6wR90G33bSTP
4SSXcQ9LjpOkT68HlJ/bJ2wVDtS+ljhHSi4E9lOuGa7VwJbiJiLm4nzl2BULlg1u5g0/WMNAbiSr
8myxEr6tWob5raDl16DENGDvUR94c7mkbL6LCUrH0B4bHwqULutnUEsGCJ8jJfCPDCkORCCiLq0h
1Z+sfbnxPA7VDTHELv6vsy+JPqTxTfZYuloiRqYKCsjyUjuyGahPTrajigrRb+HM9kkHN9JzrcIT
ShWHIhc7KJViNxgK33yCDqL8uc7HytXqTe+uj8p9hSOMEYRGURaPpjqoSBfmxG/nhVsJccuvpRh7
LeNTDIFo1hZv9JrKYZzNZB18nUhifAK75CDw7eeGd8NJepREYHpm7hxx8FLMV9eYNYljr9dyPlBy
aneMANdCTNqQ07tTc5mp2DJwi9XKhuqPMusEjNXelFkMc8tjdjcoop2Xcp+QSM4SBn02utqf4vTK
la5yXQ8U9f7xiFsa76+ofe0xxnKcskI5Po8f7mhC8FJyjPcx3qVoUwTwhsbAXI76aohfw9yFBm1i
U4Sc+ADFzJouSuuvvhQQKWvwC874RnqoHsNSQ4bwQ2J3XmI7OEnB3j0GFYhd56Db1cNcLDTnKuOM
A/0ZqZqpw7XWurRTD4jf7knzKFlwAdwvpxalWkfBjnKRrJuhXCXw0AI0YE9YLHQUAc9gD7lomyvi
By6nLfM2Rk7WFhOfU9k8EOLcNJavFBNCpNsbU94+n7Uz834uXLc9vX8vLC121wNvtKYWtI1ZUfXS
sCGWOtM6Z5W4rnXoJzthg/+kYhNM2aCkzbYwaK+gU4yMjEO0mbl4RJPJ9YCEdcqr3RbxZhT05rXc
3u1GYMH3AxXJffiLYk6cMorRQ8/w5pmr6US4EuRTDOkeahq7ji4VV0x4We2j1D62U4D/WHDwPHlG
96p0YuU6jKNFsf+MJg+l7rDOdvOhNM1SSRO6gvczt4ne+lNvTSgxl+7D1TK/YKdQsiWAYe50T0hA
yIPOLRpwmowwYvRAUPBTtgflWDqN2g32+H8xjl0VV7ZPwNxpYsQJuDcSAxPb3uqkU0x8U1w4Jax/
PgpPUhkAX5BafKja5Wauohm67+1N47sHA2Vjt/ze+Fs3cQU6lDOTEzGCDqcFpc/oz/KalrsC+ugJ
A0U2WIow1GnNfzTeAnhLc9S6ylFv6Wo8RHVFnG41AVZZ70WvHkyKDMGuMLiIaigCNLpdHKVw6hH2
ZPGJy+1kHs10Nf6AZmmr6JkaBYqX8giBBV4kV1nCFDkNtBgX9wG57NhQwjt8sg4eu3cT0pI1kYM2
d7e/oL17zYCUtgizWuqivozH38YXDycvWZWjTyyhgulima+uEZ/s/tR9VU1liloymtF8RmyJ9G57
Y1Epi2oJNluLP0MNrpKuDjXxbTpJjaYsxhB6PJT8o1hZHkwB0gBbtU71KPBYpxlsucqeefrlt4E9
AAh3W2BEdhPmGhwFe8kPwlykvHaJ7YHlEi2MoAWTMCZVUksUWOmwzSoBC5Hbh0DElNnFXnxr2G15
8sOIwXuYDOoU7ENwQ57QgI4KCG+UvnPBUni6jBO7Sz7gmhG2gdEiLecFHPLIZ0kUgk0ri5iR66jj
XHt29W/+wlSDg5d1oYkXXsh95b74BaQDecK7emWMQSaoTDwU2L7OY2tViVRNKweN93BNjXxpPWZ7
bjbmxQveh4qzqb3U6aU+/w6attG1aRnfVhBZG2CrVF6HB6uHH+m5Kdb05gAZpiGAPKdxWv8nByjk
1FqoyQIvgbebdVzM4vK8QCF1vvXdDt7gmGDhFUApBfC+3stT/9DEurpKhZcRaE9HDNXVet3WyNDy
XQCY/dXCMHdXZZrqtKooeWAE73b2d5+O1TfC9hQ7D+SXqO6OaumA2upN1Uvs2vd/tuys3UkZdCs8
Rzqlcjn36fTvYt4QkvPqnEwbt7Mrmae1PR84oR3NuNqpsOlttyM0ZOJxqHSx7Qrn1UbXbYAitgQH
sV2IKbmsvj4M8nzbyC/Kt40AIHM/aHvl4AouqQYubFVsSbJA61jKfGQhVNuLyqkV2NxbuwmZASiF
lTJ7cSYTanLU+caqqr/xDBZC/y6NjGAuG3bxuHnaoeFwoFIghvQyhk74FXWYd6p80EUY3rQBlq4n
Jw2qBAhK/CGL8IDsofiduhbqYbyArUCX1A9XdZMU/RtFoGXViy7f1fmZlymntB3qI6OOWrara89w
YynRvcnleMNaa6YveFshmmkEJ5RjxTM+NNi08J0WLvwaIo0xx6++U7ZkDf0UbaF4EuH7Fm6+53e+
siGPplZL5OuzCvHkCyZFn9eSim6h+UAVA//liKhexiNTF0ajbSLqaI8vKISl4to/E+5u3F50XgqX
FqDXibQPHF91nONqFrjs3AEu2qg6cqLggb69uzm4MdOY8I6NJNxxQLqUYzGrUBF+6v7NqXj5pODn
+Q1fYdbWptKiHtK7JWWjQO5b0rLRme+vOGzYokG555bw4kCOQHYkKbgjsssGJwAZ2C14IV2qczbt
OY0wOq+ys1/7rjRJTmYRtXUzwRs+cbS+mPTytmvc+R5wdMjJFunPfCHpCw9D3/9OeXFLUzkRciYx
BclQA9P/ArNuNU2xG3T8Mw7334voDfMX37GayVxu4A9sHFpAGAYVhqWBBar5N05R/sAV+hVOd3oY
7uaXYq7f6oLuAALrBB8weGrmC0X+5svGh6obDQuB8WuVOmlEy0rY83WnmnQQICY24+jm3Ptp+cyf
Dr6gnz6IBGCziB500lVFCAbdNZVGE3+iCIgww2L4baD3qnmnarxxtmMldOIglJcGKQ6LzHVQCWC4
FeUQZUMp5umkucz6g1DEraPCGXd1bR9qj0cOH8mXZkK7yTmba8uD5SLUTf/5JQtT95m0uJHFBKl0
DTdtyOxdhjaT7pbfintjZkl4nfexTSyS6qf0q7iQtNYGvAtazVxJ7aBAguSdJcylm2+ex4KjqfeT
lwjx+zVAl1lG65RiKqHDQ5gPRYOXCr7qkc4iGzeKXnmd87SlK0QrA9B0B6UoiLHImsWpNSH7/E7Z
aOH9LqBsePA8cJNBpZ6561rd4iMQWTndWlKx+a2cMhgSft6KrlGu///srQtwywWqfGYHq40kDso7
HqujRnOLQJJoYXObmJ6IvufLMSIiPj0b+oYu0eflo61l5S5p8w6u2SnV/33ONTpjXUAA7rTfeqgV
eJ70NdK2ObF57epXw9wN1Jq8KZ4wo7UM1xwWDwO8UYyP6YbtbuzhmSJmNucemb4LgMM44ys+Lxpd
Ltb72WkIuc2kEVgdRuPqKGFjxXpGiu8ljrKJEqx2Tdo2qJXtjLXtvS6rlxmF5PT1QtG6POOF8gn+
Cm7qMdVs4sxIix6qStBh822/esq8eUQx11tlzuh0hVo2JMHxZJi26SKJnje9TRR+9RnLUrII25SP
ru4nRFV7EtW08/HleroWk/3hAviowHnfz8b3dFliFcHzqse65Al8qMMIOU7K5RNDRgA0MjoqKgmp
TF5T9tY1lk3LGHcU+SBCrUpoPDXRwOJwSbpZXWCPU1Im8drD/feGoDcMt77le9L2COL06uHPBV/C
41F+mAIqjV1tDqpJN0f5oXubhm8xAnTf7oQWRE1DU+4SrqRDxWaI7x4NgKKUg5K+1cS9cDMesFMN
CvteEAkH8EjCwRhiuBAoBNVAe228t0GpqrP18rbnpiPubZKbsoWWooX/rfb+4w9afr3mYvVZwCZd
UGp0VQM1xyhLyHIyGa1z93oF+Vxi2Mz4vyX8emB9gPlT6VfSH2OhMWoTPJZf8bbCjX68hl0LhhFU
t5iILs8o93oDVisR2bjqvw1mII9VW1iX7/95k+vaGSzUOYhE7esnJ2qxwByQXi3rVqObhkFOu4lc
mfLBJcaAV1ltVvheX3k1ceu8Iu7fOEB+wDg1tkUF0/64K/rovGH83zpOJ3eLhQUUHX574aq6sLtH
cBn0v4j5Fn1ZQkgc5Nx2rJ3e8MF+0wIduUb0zn0DwFwbujCtRTpcHzqov/qv76BK5edAcXio7HUC
CUvWHCeNF5KVwAFHuH2zpWtrXBHvppgx9VGwR7uZZ0AJQ+txxUtKeDtx3ZrSLIE+rXWRATtEPiPs
A6sugSb/krRwAmEx60lBcZYScIcEPojvv/tslJYUNbk4/wH9/4CeGxPy4bVIbjMwUrlrLVWOTDxa
QQDhBSGnxaU3hOMdaKZr2se9cXdJa/tkiC0Ko5nrK/uF584pUO5SIB8TMXn2bJ/Sr4t6IbQkRJBS
KKX1M8SkrAoSCyUujmYEOkNsrbib2Jj6boMY3JkSklLD12Wol9LnTTrjhCAIZepVMjFaJLeSKPSo
b+zS2CbUiH7oyETlfMzMrCfbTCihv20S3kwkqrXvRv5jDzrA+RC3zq6tWYkRwHpEs3cgp4BGpKrw
QEmsv2cUJ39hm0sEW2uURl/42QDgLSDW7ghkkldVeiEiVZVVSpV76zfdh4BnhpTczqPxEFmVnJ6G
xEFItJIcHYTlpt+JnqmsO9J4ki9Gqj5xc7BjCvTg5Lzqtx2zXWRGrEsK7/jLWX4nDXU7ZVkMJ2rB
rW1YVley1kV4VNZHsU6rNnlhTtx4h++2G8M71QSgNPElU8MIzAhqDxIHZuv8LXC8spArYSyLdJhm
JS65mRrKayYG+xhlSjSQt2DK0HpSwDYJom77FGw+CA97jWQ0TqISQGH15pxf8JwLjmTXaHEb53Pd
gnoFZzu3h5oc5OpPMfNj9pJ3vUREP5Q137Aso5eaqU4gF8pEnXhWiUVTdf72pK6FdntobEpMnhKA
U1k8zBDCJzdFNrwmLUydrgcKW42Sh56kDEn/j/EN7OukAaJ2Pvd6KGZ2Xy4lb7/K4oZpxABA+6FO
hb1qjFc0f3Xj6ZW5bn1IboByCAmZA8lwiepmTJ6tbsdVFlseYWql+aMPIkrc1HbYTfry++zThZak
fhp+j/i5pVDHZu7SVN3I6/vwAg53ORzNe2gkjPpfWmcL/IU+mzYH3cU53IKtbMIWPEfJORQ0vbnq
djnLDYWo8K3dBdxNDYAVhbwhlTXZ9yZlx5l/v1Ixf9CXUVktWCCIb6YXOcJkTJ6/PztD7C3xRhXG
mkYzrRq5k894hblPKsoaPAQ1gxvy2ng8tW4WVQ/la5yWC7RaS9CsaJ0CYZCLCiw0a013S9VnQBC+
Yegq5XTr7GcIy1OjFggzQtBiWKfSyYhMcTGAYSGTcr5bgj2AFxPrHYr3qcy/FanEON8A7k0TR7iU
QIm9yud8nVLW+fku/Vk7gRR2KGAt+eFL0lE626qPDzKGdKCpP0YoAYzlqyWUyIzObvwXSqMeEVHq
0lBOCjnHLhRjKL+cNPNFDgJfupDRlHx0JYnxI72qWJN9oNddwgHXA3WwSXefgP3i96puZAb5PoYa
cORqHO14/SWGNlBAXd4QTnbSK0ybtDL/rb80dzLgIBw6LtCnHxoiXcb1qI5WynL/ruD75fSiJ2j2
IPpzGGDPR6ABcqGENoNMzkhVpjDYzVBBY13/2IEdtFKf0INKbbPVXWMfLgwqUc3oW71uctGRfG/G
uTAoXmbkbRx9sJ0KNVdu5E1sNW5M1b+Xn/iJd+SjUH1XenmuywiIlpl2TCifQN1v0IKhMATAAMj0
Ujp3H5Mt9cXiQtij8ah3jFKhyxqQqe9A7DCVhMynsMShdfLlUCUsNCMln8Twm2swFV3R3VYFsdUn
wTGHpEsAMCBikHlYBAyFfTyUWP5kgI2uaB0rFsxch8oN5pCkdBX3KrXp72JrsG5eZ42Rhd3qqWA5
LE5QY0pbiraVIngFl59Ffi2WNyU2+mscP9CNbCcaJT+6nvcITZ/SqZeahLGe0DYT53IZnA6uT8cQ
Nr7DmXUgIEbnXgcfrYzF6GmRQlQhUYooAtG3WuP3+6eppP+Rrqr9Ie6OvoahXbKpTGLWD5rrmpLP
XFdqvhf3WFhl7JHWBrF0eEjiWukr/gb6CgMSusfH22Vf7XAqmdIapManYdNIHq6HMZbCNv+LaSts
k64z6L0Rvfajz+K1m00WiUq82chgZ9KNl62SLtIXrXuhl3BwnIQ2B7t6Zk9e4bW2z6mKZt+/sPtm
VwaQjcfIpN39Mi/diFv3fk0t499iWAy188E8lAmYb2AYYzecrbH9T3dlWUgwIwXp90YvDYx7ZHtn
bsOFiGVKcD3nN58zD9rmpA7wJe3Zxx6XI6RV90X6bDKtoX4qdyr6n6opAXiAGrRU1ogjAbDo6tEf
9KnuQ+ZBQhblTVVY1Ue0OV5lMUpmHFo4ySaNdR5rBDiCSJH4bpeUVhiFhEyXw9gFX6yTQww7fxmo
aAvE9++xi2WuNfvLgtF4AIoJS/L6gpucPDgg/tbRF3fbCBeCdt2IK1Fi+nxsMVYYce43lyhaylf+
j0E3w/9JjlsxT91Vqk4bm2bDyBpIGSKQ1QYaABErP2CmA7bEDaErvLV5iwDz+5ZbkOR/u/vVWbKd
DgC/fUpNRwLcWPwiXnoFGZE9VuEU5j0ldZAflKDv8BPQfYAIi3ZKjk2FWsZh+eBwSRBVGE5FKUrF
WDLip1ztVBwXLCUHOP5gxCPEh9XpfIAPiI9N7gBiFbYzLrSdca2x2HS0nrvkSG/g5Aow8zCZlBHq
4UHsTsOp3yWILAEDUAf8jtPiZtfcNDv383u/ol0HydsvxZxKeiYT46/J5FTl3q2wJ+8sJZHsDPcV
4Vuq0AAyMeaB23ZfUtKffh41+x97b6aZsP0bUmpOMO89ib+gFuhPuH28GIicjrIFU0PU2ccsAiCr
kfuWzEDFICFYaDK7itFkpr5OH5bAg+j3cxg/1PSDq4xEfTjGz/wKeuhbYDU9F8aktTsZdmalwL8a
4yzIP6SM5AoHSnKnDJrIwsSHO53WZsn/dRqyBFKnI6pejJw8ov62fSGyhHtMHJRjZdCFAYzdaBYN
TDHocnGZw/weiYUYRCSelGg7YwEJF8qdmZHoD8R9BVNiLUWZsgskAMXgqcD8oVtiexrDRtsxWPwF
BWWG29UEloMZAvPhruYmGL+R1MOILXsaiQfH9Q4m9koF+7L87YkA8dS295TUx8n+ohSUaiGxZXMb
IRyzHqCjYY3nOARHIksHA8h7u1ouIxOBnG2afISYz9mEsqy26zuvitiHxVOj2KzxtNzL2DQfuRGz
sq5DxnGzvet1OGCLu7mZM7l1gcVCV+RTvWKPZPfcFZWroHIoVGTPSdc9Ng6kf7XsMNLnRZdnAD+3
qA3r0yqGy9WdRtGZLB/442Y3TXhum5z68qACqZ1yty+4awG2vlvM2AV4K+26BcEAcVUegtnhjo7G
SN1zV2QzsS+h/kiR1YsUSZy+rGjd5+YXYINQa/ipkjxJe9FalRciueQ4OAmkV4gNFiwwZGqiST9G
xT88LO9AIcPrsYb6xgJOEo0IJ9Ex8NZilniiw50TzEtDDbUhwsbZq1KDJsCI3Q/PKp9iXkseXS5T
c5UBC8qz0KsRfQpJ7A+LoOYl1kJvcIDTmKWY0ZEcfdX4yGCJV502AX3aeLSK0COU0b77ouzzAHvE
OjTJngsy+h5D3D0dB5u+e6k5GapdvbeAF/FAlZa1nUiE1hF82Meurzy4T9cHrelyNKu9+46kucmT
c1UT4lZlFjetqEjJjk36FsDKZYtXZ06h1zJwOiQHEevJ6+FztB0j0XtR5A5Ytv4Zl038BL2w9y0V
GpqqYd9qWZK+yT0eFGk5porzCfzpcR63i9+S3VaP/MLpixjPavWYWlH1sVXG6g1M2IkFTKtcfIT7
1dwO17bAIjY+YcoIX51QJ2Fl0+yOdXGSBkH3TlXLkglvP8ok+kT3/UpoZ6HqFn8/AcX13T0vo19l
JuW/FHw9y1oLGGe4DobxM3mCW/qlG9HnYhhvtGt+UUkK3SCHpC8hwV+veuLX21aXNXO63y6YTlD3
Kve8L7nhS1CI0LEqAy8Lmz4sofqwV7f0WrLAV/E6necRKrPJu2wMMIRqYupmrJRTMII/1vKpVx+Y
7/oKgR5lOznB05nMTWzfnUDNIF7GsA6xFHjoFzZ/veq9n7Zb6eGjkCP6cEBCkP59cht7Pq/Q5pcz
q2qZvT4Z4mCS1d/MPqyKsuU7PM+T3U4hCDi14+xz+HojSZ5k2FJgakk5lakuNqwp7DXRvODGFutw
Gf5Z8Jpt7PTvEmIE/3MPF9z1+5nRniqa8doef0VCFDI6uNybLq76EPyk5tvEz7t5k3msLcq/4Wny
OUyYSAUxeP7Yb5Zv4q6pJZy6Qz/GpdW2NNP2eZ/Keia6HKhQx8ufJDv9SPZwNcPPch4q+1gVVgeD
xjyVGS1vyPwheX6xFd4H8Q1nrwXF6IE8fgy5w8g/vi9/fiLWE9GGIi8GWQSK72c2EqcriSVdam9X
lEGsqNs8Y3+Q1XpYKgVeeC8JGJ8TLGN+ehVNw6wcJJzYRKy5xuytXBLv/74L6I4KI5f3l9At3GLQ
tRlZZuccMiYXv1eCRqnbpQLcVmo4VaRHgeLuMU/cPeRIUBCm+GGteBWv9pk/u/kYMszKRdaMiu3Z
HrF8AEL4Be3eNJUMn7mkr6LiQ7WYlmlRnR8Dh5Xg6HKtuY17vmj9m7kzBjiUEeTEXMsJHJ7OyGhZ
HEu5XuHINAxHJRTOiueH7S6RG3G31o+BP+1rrnIdgbhfMhumFPbB9g1upsxHAl1Xbp1CE4HC+SRO
TRRpA3KgQ7fZDB4jf7+eTm6c7JeuaWtdUzKpEkiMIASQRvgpn1+zZ4hJGKwAgZmNfgx5IKTzyoZ6
aJ/2/4DoiuuAv9aeR3xyfHSs0Z7+li61K2Nsu9yeSR0TalSWVbp+RWvYz2KWrPM611JTcFh7hYSh
uWqqdV5IvO7nIXpuGPEz+Tmg7Ten2Zm4hKnumQiG71MgrZ25Ald8SjmK6Ssq9NHiDJPC6Fe2HO3L
3ned8oFGxAuSKITfnT1yR2PcWU9MmU5+9sJfoF1CYkcinxLpcCNFfDbw64kf/W2mX6oijGPq+/TC
NfudQM54Ql5xNue9hi3WplFReMm72V/EXXAz6OQySlhAkynYCra/wZ389B7/D/c62xGuP6q3sZNq
VgkSVJeRrHEk0+6LMfSGXjPLnHGuO+h2057Px5z9IdjZ4yAfSgXdxPLpXOXI7p/ZWPGPealHjk1l
APHEWE1+NAZXboHASHICMDZ2W3GfzLFCUshjXsTalsnUE9d8gebBtL+G/JFEryXoJRYeMVXNN75f
vyA9S1d3xCgakfoSgItkKHFDO/cZWYFSSrVBKcGINhkYPBNVqfjtmJqIMxV7JClc6viCIx0IGI3Q
m+3HwzM0qFFCeOAVCCk9jJlVn53+r/VCxYkH0dNv+XlITv+RYCwhcToMOE86hWDPr7i+VTUHEanb
GXR2/k0JtVdPDiaBsySxm0s3ZRjfIDYp0pv2cvk+q3iMd8Mo/UiGHfkZZQNm8y9DIoXEqtKTkpgz
aUS8zA8xo8ELSrddpMwBnjL+fUrJzOYNxeIhiq1D6WEe5XmtRZIJFqtndlhPYvwKYHIY70ol09Cj
MpOPg7FMDIEgYc5ZMZ1SgydmVLy6Zy0ap8XjBIIsjizQuDRnlOKpeS6JVzHjKvG9ZYPo/SelOHvB
o4siLEwNQFGDRDQCNURL+oHbL48susHbhxduYIU807iLyD1EgOh1L+UJYoEzsvFeY5hQxPToodC8
P0pi/epCjDQHYhfMmJr5d9WFHIGMRta09pjqYXzypSG8w/odrMMbO6FUCmcuZRkL449znJxdxvx5
kmMltg5xvaVj36wqGwCIqLXEmQEY4539cQgFP8e/P2u3rJDB691EZ4cR03hABUmYrY8CdWxFPMoi
SEfgaDDZHi1UXdu+UKwpRkU1HrjAA/bQBbFk8TqGgKXx4ZnVud643OD6k5GuoitMW61ogRCHgiVb
bsZh+n7xkCz7GVHizPEItzMwWmXJIoxgkkk4DMnASZoZze1G3x3XeEXJrjcmCwd8In+YAKPqaC4d
iSoRFIOA0u08ue07Idsq2Sad7am4aqxU2KPMnkvEqARm2G4r0p4Yw6QZ4B7ouuA/EBcz3ehBgKfw
z9t6jVGkPgorpUEJkUIBsPRwfsLddyZRJudD8gM6FZRKqW//RP3F0f2DN5fHNakRctfvTKeMJ5Hw
8MNnTJ9JLJ/G3mi4s9Y4ulcbBa2qRniIS9wm7Ubebd1nyz0Vly1d/HO6QQLo6uX+oYjlWip6fZ58
M1vg3CPneM1+C4R/Sl3CeuGjCsodOIA0yei9ykai2UBSi9PxCwxoDwHR5yPjC8UwXfugjKJ8kYrA
TB4qzfI40BZOP/08UM1yTAieqAL1ohJwzkrV/bW/ZxhW+uCGIuBW5rmYHsr8OXC1XP03X/Z8yDMO
rRJWYgRyslDP60XUQIYaK9xfiJHjnicxIykYGsvASiOOc6HGb4rOOP5VrEbT72KvXsOQx6LWlwvx
oF3j+a/H8B3HAnNIjX+fC44qDF4NWL0+EBj6C1p1fsFPceowT2VuCdIYdlbHZZBfAN9WYH83XscR
ZIH/E8mbFUmP7MccUsjmW5KYsJLE+yd4Sq0C7q6Ob3k4mOJHHn5tAfYek4R/7P3cnGeuDzLqHmHH
bK7NjsOoBn7u0Oyysn669JI0rezLQtMqoqNy+1aN6bWCF0WspixurzqbUpzU+lo38AoM2z9+5ziM
ozw748UUvST8tq62tO3u9+mTniXTxSHij0Z4KXG+HsqKPQobbNFWK2/sFcWowhcH/eLe971NtRZv
GWFJ+HDD66E5GrEakywHg/EpxG7DxMSbX/KDkS0ufnHnjKA1AR65bJpFJER3b2ZgU4pid9RNKaUl
poYuP2Jrehk6s/wts5Y7y1NJYoSW6TMCTYx21cOKqymyEP/dIB5F69+BPCYll8kukG7cKjOijjTF
pnrNHrtwFxtjLxVYKBjcNMxrvDSyifyaBwt99haboB0vQuLaCZ/yxV9GLssJF0s8/s1ITyJ4ywCY
PMQJ+z4Ezn044WUdMjb03yoRRvD9DvVzzTCpwnovEQOMTZ3grHrn3rEn2GfS5OE0N/Q9uSvgARa8
cIaIWkH2uiYNaxSghkIsaHKBkZCtfojKlzqC2PTTO39tj79SeCi7L+ellaVVHrGe0WTXxV6FzT5N
vT9bMGl/Nxk7U01QKzm7dkkUJTuBVo6R5C4u84eHVjqPdM/p6785lnVcbD6xRMsLm6jXuv8LeTWV
3DvJYlXFKGLhYQzdNd8ytQJ4cqHCn/yqoExQBuVKF1nsp0ope9pNS6PlRC2aN1L+QZlILMwYoZ8e
Ed5VVJg0IVZCNt6iS2kiIw9Un3LWwfjxqAiMiTX/WnUlEYVrHSoqefgsF8HiiaO1DEnLp+nH2nqk
oCdB/5l/Y6mb/LRkqNkJS9TNskpVSK6uLvih9+BPeAGScQEZtRoxceTyNe7oy3SunHo48X8n5Oun
P2SzxlJ/QHHNwv0KsDPgPFsdOSnnrQOPgaeY1zGad+LkX8z4K97azNVHY8RuKn7LJZumYrbnwFP5
JTb8ImXBVoqRAWQ7jrx0ZyGqU6mdN6Ct0Cy3v7fUAV5NuXwbnHm0gPObKzJoUKm5xU7Gdi9f7Onk
McRBnGKMAk8l7lpF327ikEPHY7t96Uj7a8t4J1aI9TDKott16F8MZPRoFXM8XsTg7/fHsGYI0mMb
JzM7cDMkG7ttZPfRyYVhzS8EmpE2qAn/ZX/fDBCn7Oe9+XUWshJiSZCTmXqCrmajhpLyZsCNLVkf
wzaapmvQVhEwteyq9twCejh632E9KyO4z2WXaWX1uoeHSfQAm4n0xu6M9W3vI8I36Jv59cxGD+Z4
KPSjYSqA6qlk/pBr8w05j/XLcOrwi3bj/u1N1Wqt2s7lASOf5u+ldw/if4gMWtNj0RGhjps85X/Z
8KwmCFpaU/IwHCf4gBBI5ey7dTcUD9kXNiO3ummGqxZ7hNfvpShbNZBIgR++/Ck4jUefpJh+JqbI
I0YBQkyHUx861bd8rz3n625Edd+G8u0CdmYJ5GfMUq/SsmtWec06YZiZWzsHibCm3To0p4yn8SfL
kzi/6+3DkkxSHzBTIERiU+doUTXiOtx5HiQEuf2zFnQdOaavNEZBrxhqhDdgdMBX5QNHQ54YfsY+
1I7n7wkprJlLI1n6oRJtJoh6drY9LS3oqIPiN361cH5Bnjncgv9qxNIQeHXksaRML71+iGwSdpta
/FQdiKQQRpt4Tzlp0Y2GT9zukKWwbLUaJpue3PnR6aVmZO0p8MtWi6L2HvgddyzpmrQRkfyzF+ve
R60T15ycVzIX/86RUyfIzlcxW31KQxbfoopztvBpkn3QO0loZkc4ovTBH+Cfx95Jynk+rfIczmn7
mse64E7NcvdvTdSnXwGl5mtto3F/N1fu1QS//8tMKQDWw0gsVbFJ4fcGm6Z3/cS7PgAnS+0xSHIc
5hjLKlokS3oqYgjrUJSfGuMhxrActegz/EO+N/4ZOqKI99F2cnfU+k8wCgeZZx2EW+NHtK/wl1NI
VJvp4JVKyx7ME7nPnApl1sG8/OHAbtbG+VRNR/n8uZMRdNuIY1Vki3C3sHpDedbKzPh9hXVrO1H5
2QZBRs4D/2j4+dGXekKNQmclxZUAgft+vL6cKXnGWJdrf/vswCeAkglhy6lSfwNM4smYBz08ZhXj
gqSLf51akgvnE/FNspOgef99Q5CGg+Cxw/rgVo7UezCCgtrgmH47wKO/aI57YrEvlBlBwPhPCk+4
zRis5y32/nzG/4XXbPBRdZSqTYXyhoi88qLSDjO1h+681Qy2JHNt0OOSMy/9GPeslDAlnlLPAKCm
vssMuofPuDZwkDV/JFuj4ddRuo+CT+mqi/K183ZJGwF7EeFQ/GLu9wCLpw+jMH/9kIn7VMzB8Lut
HWZYH0XLLlcBCQTOkVgzrnHqlZlGnRQ+wv+mXZ8k8wFXC988umHBim0B3Tsx/c3iCwqdEXRbSnXF
OpxBm76SPgMA2C5678RhpTVsJyReXgA/Bc7IdW71odXj2nY375LNy5CYqU+NKTMHNbygNVTGa+WB
XVSOy8ShiN+nBvQMLTrPcq8VL0e9+I0h/nB1aLAZWdL9Ci7wOIGwPYTl8JE4bQlYopSPsq1RHTtC
U7dZwniIHDUhcEtRjeSm/WmaNKeSHppnpKmDzHl4hmbCvHKdM7zw1g/MQUeYR0MkoutAgt0RJjTO
x8giX1o614PEDdB2bFmpBOkLs4uSfz8BmHXGmsSgJIquJEd4yjT5dp7ikpwZ0PB3j9HREsBzT5JO
RBEtV3JXk5Lw+oj5FfZ/rVBZc3QCTkumMy0AL7DpDB621ohjegkc6igT7Fp1PKfz2xEOGvm7a1qG
f/JvLMWfWOkIyoixlZXAMqEK91SpuT21kEH1eef+3rjzDUrNKx9YE61ZBVTWGTqL5Xv5LTdWRMwj
IdjtjrQ9AOh5debZvRVo1jyvs72L5FgtqwkMCR9HxxSDGdRxAYNOS4MAffobCx+bB0FxkoH802Yn
vCds7abUqbrg7+2yvO8Xbf14Jt/sEt21CRKRUjotTMRsL1FP/jcjzA1poNe1l+0q7mXaNmBFeZx0
AU/MOFmZSABpEFynSSp8pSwof0LdImgcwOKv6VKUIv/kCXZOxwE1PrKmpo0LpH8vGl0jgBZ1CjpO
QaW594wQDyjin7TgOFl/S3MdhhoAzdXodwdMg166bj5E+HqhX65ropEOr6iovz+OpN3mAZAIobRz
4y5FCKme39Q5NLPxptUVKEc0bLjuCKSXruWqSsrhqoDWlV4fHuGdY0PcqzMcyCrkacN45eGSsOgu
UxzAFwPzjdDNPbFWfdSvCQ0JucFoyJzyoRXuXej0K+2dRRPYq3clMVvfrN741YJd3r3FvwZLSkj7
a+/ZWcM2E16/MgG4fnRcUjeJbKBYono8kGD5bK3ZreJnZ6hMOA/Js3x3T29PEwFmSgNsfeOXsLPu
ipjc9Cd87iY4dNz8OpS40pxtv39n/6t4SXoQzfgdIFi4plfAcKOx/3pk9VEZ2cSi2SSfNroqMwwS
jUmC4UurpEN8lUv1s9sdxFglk7V19K2j0w/dIW5dPiGnVzVjGbuZEyNEaH9DG3U7Mivuf+Nq2U3S
OlVKrCzBF4d6ocVWGLjYHdxN91+qHnLwSZfe/9J4Nnrmf5Kzj7U856w6MpA2rgP8dsuvi94GaxL3
E1hYxrUoSOFZj/1tPTtMH2X5g3LNslHpmmJl8mZrrOoZQ6ySA0/a9+FRLUB0qGntEkYcmmmO53lq
uZuTraNFCGC8YnNWkPUEjDwTla7tG4i1QzSSKKJxQ6mDMf3yxAx8R1p4JZDRNUcxheQCJ+2Ab2Cm
FU5tgzijpF1IckUu5X/tGTJ/PQI0KPjQKKmyBENdMLsBxj6V38kd5fMA72kvbHOBu0aUg0XJEsKk
nr17nHbpkbOZf/lqRrxpthRMHUD2eXFLUadtZi5rZQ/eSN8lqR4mmmQgqLFNjtzntmAPFf7zaoXj
igsJkH1xHQQqEPcHuDhQ8+dNyB2FaKlnf96ohj3cWXtUjYt90B5ZPaA22B6sBBKca9qSo22GnoSe
oVwlspTaQ7q//sjqyw0wwXA/wWRDGUhDG5X0CYqHt9/ZIa3lzwGB1oJc12G/18MG1JVi8ugON7V0
v75QHkB1lspCNZBU2SRwpFOHtN6zs3UXD128aOYOG+LYHLcWAdlismDUJ/opUzmgnZsNV//AmxvO
d9FC93RricL5LUbJbPURRuhC1YWCfuYcuSW3e28bFs8z08aIxQ0U9g8jz3Uf6Su6zohKzDLxxKT6
03Yiyy6QW6j3/CVfsHgWWiJ2WlzAbZ8BAT1sz3lhS/Ap2iVl/FqS2Z+7zhzLfs5MGbnFHlD9QpJd
GTgInWyE1wfhTO/EBukU9IYb7hpC7KqPrZW3BpUdJ+ZrH+EpZcEFN7e9rvd6b3lixegnZsX9z+2L
14p4tpc+7NjzKyzHxqXNy+jJp+V5ktJbft+7D4XC7iJfX2KV1rXd660BZ7ReMLq/NXKabRGHf5gp
LzjfgoBJcK5RFPI9+fPixg220y3Hxmtjm6u0R6HkPT55sPgB8mNWMwGn+tQOnFkw7KiiTlPIb1Sq
szYP6K5dztj9nRHs6CNzbwkY+JkbDPO9WgF01wjRjQU87SJ+pXYNqCbo4vIGQosd92uytPTQ6rFF
rv/1hqyCV82rwMteZdV95l8sAqytRsVANWUWwtOoBLuxIXvz0mfXEoMOtE7qpxzcUXuqOLFzibaa
L32ueXsugQykKIiZ/je5226ZRt6rXssQtmY8dbrpT6JE1tTyLe6J9o8KN2zQNYGSCq0pew1LtkBc
1X2a1RsY5mIbdMKlSxVE+jdhtW7bNeOGUUyJcV06UakR5HnxejhshY3Rm+ePMsUJswOladZWXisr
8AZwFcq1kQJzeqE/pkWpuhHK40w5MvCKfoKFVmOMg6HgO1Z+o9tUhmUjtePLjaLW62pwp7hM38fE
dD5240nnumL+FJjop/e5KQlGOLO7wrej7c1sHiVoBQ6vhv4YgrM6nBCbhDi/m2jfQ1JC+wwN98r4
7rzLeUdjkbmTgB9avCEUD5lribTPi7/zHUZ46wFZGnjePfI2yQp5pGdqA9Tk554vNaIKDXC1SXNC
Orc7C4rTtH4JWGClZPx32d97tZkNL6QdTLSdLMwBrsjtU7Xvf3ojYUojbpjZtHtzT+jbK5njFbpw
GJCYJuyk7MH6sDCQY+aEveNfU1xbI6htNx3GyVsvQBUJpDYdbQUJqVBP+HTEtDlEhowXOXGVCcoN
tU2oqdgJykyBwvJWuD/2oAlji9M7L2e7+yzQmRB9k4H6rrbO/5m4AKBGkP1Ecmp+iJu+xsQLmOS5
cIrT/wI4W66xlQnfgp7D5L2tlQI2IAApOEK4a7w5GlOXMA/+FxIPtDKozEZ6uASw68lPo7gmfS3i
77fWyEn4aobtMgJ3ktKysGAm5qnTRUvpEwteLuQNeGAnfQd152gl/ZRc5PAn0MfH397uSpLMjQYa
8TAPQ/nHCwbmxDH+i1KJuH6Iukxls0mEDuXj3d3jK25ty7tCR7tCofdV/KxpKPFx+uCvD0ywm1nk
RkmBfWxnOSqTJRkVbebQsYJPZPyEYIxnH5RBDdMwsndOrAicjO5oHviBunPY4JkY7gt03z4Dm/Iv
oky+AE3qHNK2orIOgRMVxqMHwIPOTYq5k/tRfPXSDhNuOu1GuJElzqCpvEClYmnTNnIegvioQoZH
JkjBNWPR8qykEwqWCCTe0pcAJqEwowFofOwJhulFBpFR7fQ40kyq5BstdrSuCOkEvcXSWPmsFRBB
fDeOT9yk9WDVYTSdiyXH8vqC343zAcBdaoiMLtpCuc7v5ar0Urq2h0DL+ZaU1VJjXir0qydTrDqv
uQqKmKu5Pr3w/VKKKES1+oHk76IpjTWi/MjyHqM4iTd2MbE5gAjwOjqfweEq85g+1S05k15eIFHc
dbt0QL1t5svzJ8Urv6Clj/VXur3tMy8RTQjH/ptxuIHUzl6oxqvj4LJZAdsh6aJJAC/q1GUMPLgL
iq42TSs8sVfsdqJDAB6IVXhLjIeV9/0AOfBWg7O7PesP31h96k/iQEaMyTUdt7YNMTU/CEbejBPr
/EC0fEwmeB0JyLo7N/IhYWeMm0P8T2Ou70tLyRmhYliBxmgiVzhsznJy2sh//QqiSO3jKOb2Ejyz
IabDA7JaJdUb9c01adxS3a1H7zD58jNPumyZcL4JBbpbgpx9qnnn9yCAXUU7Hwj8uT74Z+BTnfRc
H72njKOAKx4IixNNtJvq24QUKm+Zy9VJR3/USXjsKwPBjsFUKNUV0Wzi9224mQWi9uWVx8D6IJQO
glygs9QSuKzR1aw+mOQkQUeJEzep0g94KHp8Ur6G2zlTe2J93cHIDD4n199DvPPSSj19pzPTNrvo
GrZLXfsG0ZQK7yvwtdf1zB3mXL7adV8lvPOHtKVhY7nliDyUdic9pA08XRRk2QynFBKUztuGdefV
iuK7MDM95NRUuPlUXB13oNVGNJ/7Wtj6Hq+GUU4H+tgRaodGcMCOFUmPzF9k/NmiIHADy59TLm0W
uh0qAxohjK7gB3E6UGp+Za1mPixbScOWHrRxStbwHxjaaYevBVYDKUunyrJ75jiMT6B0Jagi8Ask
8eoGydwk2rsH6blaGr5j2TiTQvlQjZtbaGQE4DtjvkgxyW5oebS4SX7nBR27/NOe1YHbhQRaS0fI
QlWG0wdE6nhOMPEOIKm5i4WtSHPp58Iz9zRCk8YWN5B7mm9wbzUqWpy3797fkf1uAfRoXWe4FYAd
4sNiyv704iCRuu/a2bpzCtkrfo73jtgD4KEKhIS34p/pJ66UOaNjrnUPVdnWtaPAFcdiWIFugXcK
4Kcm/DFY4ASw8wd9rsuY3rZfLxsLj6iIcoC/dfFT8qqK7WvQ0vfk7RwnT6xY+oeA4No03uOaGRsa
0AisCKuq2Qa6144ARxYLRojvTUPx4sIo0SCLzy7GCeav+2VtD+Y3OlAXH4YQii4XrsAlkZ18mGLR
ScFiwq0bxJ62BfrwxvOjL3DDTx8KbTa7E1xvnfXBC8ZslA7ooi3d4q2eyQC0afifNT/CXkafbhdt
Md7rzuZGhraD1UFh16l28jfu1GeUZWm+pCuCteSBb/PfOFY5pyrKgfJjXtz00tZAPCQFjoxsJSIA
NMWIgyFNlYDLl/Dm+aV+MpQM0tWRY8CNYhOTJMuLNVEjKqjmQZrMQPVXChNSe2WJpcjLdg4LhujU
Eh4FByzCs1bIFP39YhgDL59f6JZG8lL6jdJdcUxXATuUeO9+hsRNpQ8MOAX1l8J7HaWlDLRUQ//Q
QQlCa8qQXMpvkWMKZdLkT1JGdbDqO5FEVwg6E9u2AtMSx6XuuIrDSlynP8HP0gzS4dWohUj2yXSY
5f7rd+wrjJwVmhLaJbt6rbApV3scVI9ROD8T4MJNQlqvzszmIn2P4VV5dGMR5DEDSGI57sUiNmGZ
Ap+5Y7FJ84qONu86pqdffDdBKZ7d6VGHWmfQcqzT/isRXWn8R01Iw7tTi58V6ji7mugw1JE+4Fn5
tpLpJKzzqf5q+auY7LyBXkOK2P6Y0cjaIPxlWLYTW8Eilf8MTStKpwH0dSwaBPj/qvbW/NGmY+Az
FNVJoOM+zT0SNqKZaXCKwPo027JoAtVK0gov6G3uZHm/2AvtbXqiWLaJfLDVrY8MfE/fNkAEEP4Y
VgxzCb8CaIqlQLWnTkvzGdbMaH3168y3O9ZuULn/wP76blELAeiRLuWDPj1d6P8CRmDT7ioCrY6A
acabc6Bh+eT8Hk6x1ffsroF1vxU52gxdRO4HgGU1iFZij0urq/fTUuyFHzlGD0iOJTPf7bZ1U0I2
9+1bJvJ+Mz/XnZf5ADCtqQ+SE5PP6/ZegzNTnokONuJeHUW5D/UvyalTmWaEv532vBW0RjSgoPk6
45XRKilMaZc2Zj4rCf035FXNZQy15Q87lusmG2J4j1b0PrworSxfRsq143QHDkEU72wYSfKcFeao
rZK1Vp+pEklWQb57jO2DWj5akbHNL8/oM5OvIAqkaezImuUtgvoz3bXNIoaRK3G6bux6m43bcvhL
X6JRs0W47LfHGqTuqaMGwIddhAC5+Bjz7E72KC5q0E+2jMCBO/Fjh5ICLsf3OSvoVbvi12p/cfvS
F4w8fmUU0xDS6jJ8OqVYC4H2JIRXq2OfEw2gPgsH3EAtLQJCYgk/nM6vV5SbYlXahmaR8tYAmqvV
cMvAJfkSP7hC7s5+AVfQ+y7OVkDY9PvnHKziBmkbXdUoVz0DLQmdAqr7rsnnQr2c1M13a0S1PAZV
Ui/lVM03XcNqfVWalbG6t1cgO4z7CvrZPIqACDORDWAc4RW27caEzUeNlqSKamCZGMlVnk1a8prb
s6C0AZ49X6jcB13zEMkjp6I0Vw8CGkjS1sI4v4pmnyKSsPIhE5j9eDxSPpEIDQcVLiSO8Mmsgf4S
nxBX/YM3qxS8178wiaW0inCBikuIqeqQz/591Jm6YUm6Zk4LjyQSFY5nZ8FQdfPg/RA8+t+qOFsD
HbUByVnyEmIsbLwqpMZeYkuBE7Jy6NrduG+FcuPcScpbCYoGb2IFW2mEF3e3NQE3q8p+lnO7ScxJ
WnqQq0xaqynEWdBbYd1ypvdl+SVGWJK5cd0JRtAMJj74STngGunYM8Z173Tp3/qHi1reaWM3J1fu
TxhwasSaluSBqJlMFuPID7eQw1SO3+8FbXMgwPOnWwPAr8h/TefSDHjr7vki9F+1F0obKYw8bA/O
8MdKmHv2JhUnnIUyI9Ktk71ca/0GNzl1qmxyYtp3jcOxc+qMGOf7yjF5UcqCTS1WeeUXQO6YUUSL
TyT5v/MXvO69DYNbsdCsjE/qZ+GKkWcdCJVWVI8Z3MCZtcNcRSQfTIfSeYpG6FSg+KezdaG+ZwpH
jCRtYZ5Q1D+66mJlJ+wKD3LWqh1/7YNNTSKBraoR8O+mTSyhkwliZPQwlyWnxxunMP131xIXxJ/Q
lt0HntXBfE5r86hVSTjQHTPSmLgOdZtE1RUsHBFm30vku3bmIuTbadqE3mSmxKS6uWkLTX4pnRNF
bsGrKyi5XTQKlpf9Wvd1JJFQ3F5gEEyNVvCErYgMIA82zA4WCWXCWwy9IrkXyD071YVkhOSoCkkV
xlAHSJoBZJGMDSsq9o5VKnCq5HIAeiwPPsWr0UUClTl8G2jfO4DyKE6y+P30W2pRnlUvNC7ylYDm
8caIQ/xINlnxM/ExtsRZmP5O1XPQHoV6oCXYxji0rIPKcKXo446y+ZvJYTPf/qLe8Xlp3DRMA+Zj
ERwIKX2SR6pw4OAYDsT290F56aomPnKpm4raTTw6yC39ztYnpwZdkp2vEcNogYwXQsTsvK3ef1mF
tfNxQY7sD6XF/Lkpp202eflH42sekGuHoPfQRaWk9Yx7upYvIdu6Tx8VURRKF6ZxUaOmzd+OfJIr
z4N7zpnMB7oulbgqeoUvaoppicXhfrGkKNRzMNcs589x5keEcJbF9KyCix3OBFwti0b6vviIaiDO
AmD4u819QqUA94jBFTb7CKF/IbLtQO0hgZZvUsB0lhzJ/tMU2tek0irH4v5EWoGCfFqfle4kwl9V
cUrSOUpjL54ORF6w2GfSW8s1nARDuIZ4W6lJQ1a4tQhczQmLXTPjAGoVeXdyNwRe1/pFxg5w96IV
pke5EeOzdCF2YsYXtTsFRcBnrKcM2FnnR6hbJQ+RTWY7228KyM2f+ZmfO7Hro+U6MGLrUBPkrDx6
3JO6qZt038hCECRfrXcojJIL/IO4581TbIrKDBpEkcLmyjSNeq5HrPJOJVELu7IdygkHMBp26HLl
ePFH5dk8HVGYmQMnunvVjLIaD9xAr4wSOyEvGfg7REvs9kDWsQTGlE45fL4uo9DvexQ/n2Yj0g4+
+2oaXSSzXFF1OWKytmnq+gQBKANFxdc/ZOhIOEkYizF1L9ecml/3BGZghu+lWFy/g9Kzmsfcpxed
hXC6pwcpl4BfuqgLfDehPqRxRhrgJ1Sg+0xuA9MKdXFDSp/OCYvKUa93Lv/ZGl5BCdMsBGRk14UO
VV6l2Yp3Uto2e4udb6CGKYbCFk5LpcuKgM8ku0wL5sfgt2lVxpfad8mooJjh27GPtBBQe8UQp+u5
Va894Anc6muL95iZ3xAGS3/Hbvehlx+QrOVWMEnBoD+LshzXlK11ov1xZ6MbrKxf7+OAFoZwwaGD
MAZ54xrS9wv81qARDLq7mPo3UaOlLa5lNIVK+bRxYPGiGbInViyKhX7VNHzWPnj+NdYjSyxZ8n7a
pS3r51s4IaI/L4aVAnHL46G1fXp3g+EU5e+cXa56lO3r37rNNMBe2r184TsC9vnc5miH4A/cRsn+
x7bBF40nMjfhUQwYfmNk8A+meixu1R9vwSNGr9n/aCWdk94mjbuUW2s5jIGiNktjmtiYRjE1Xjdt
i55hE0s0rwyompkaOiP7oYZibOwEtnX9pP2MeTj21sAOR42FoS+s5vO6u5FBgJdKEQ9q219GYOfw
8Ld1pOVKF2AGl5/+scCfa5ekaqQsENVp8kEMJiwRVBEjW4j5CEiQACEhgmUMaSmsak04O6yrb6Zi
5pLR5bSoTHa3QxWvKmu0gGRCGiiu7dOTmpnYkuP2SAdIc61Vo254KCg/OZ1gnCW7FPv/KbhktFN3
qWs8oRktD4lU0jyVHxKAWJ7DCDn4jJItfQVjh9Ip0sxOuJl2vJg2hjB3DsMWQpeS8GvXasSjeody
HY2vUCJASUmy+/xSqUN/DWfJAfmtheaaXd+wDc3cK8st7Q6p+Vfmiolhcf7wvcfSWYHxGAJeHSLF
P1AIaf64KpPm5k+pmWul1KIw3Ys1GUsBGvfmR4GMVLmbpjXcYow2A1Nbuk3WPJVgLiXur4yLNc1a
8BSQB+jNkFjrhTsVAn3avx10WGow/2ZH2PcDQhk6fvmbiMkyjARAep5xG4BfpNCfDYoR8DLBg8+m
4q8OGR/An/JqCRX/F6uZLnMKopKDLpad/Xlo5dLcVHf1Pth+/u/sBe8WSRBIMSaQQM0+NbtqshgI
K4UTUAX8hf4MRCda7Wuz12F4grYsLOYCpeAzbfTsC+gtjl1OSIVouUbe+JJ85ClylFKBI7OYjlnN
lfAX2zDOgB8Y1oZ/FQ6iPzm0exmavogX3giICTNVwsISZ1kvjJG7iFciIi1JWYfGQVJcTc0V5ZEY
t2UE0vPLJQABA3P+ABKab3MklXygPeU/iNYM2eJzrCLW/8FXBm5rTVvu/0A5kAxaG1Vm55awCjz0
I0KjfyGg5S2QfpuXVLMtYeggJk+ueUCcsZ6pjCAmQtqOR7kqflrDSyLsiTsKc5LGWdzJRRkYE3ci
jBJZd0ssUaGWf6BU4cq4nYXunj2o0+mUlUEHdJ5CVc1HZuR6F/8EyfPYEid3hOVDjewnC//hXnKV
wnp6/fUlx18gkFfhvktsdQuULBi4Q3ypKie3h3QArEJSzwhg9626KMgk5TJkuZ6tfkrsgdgbdpsy
zVOseSY2gniCf7pYwALywCic9oA++xGIBkXgxCYg24hJ/D1avpafiotb6RE1PWCysTa7ArbaMZ1e
puqGuvMA/s4eMk1Fp6A4sx86p4m8vZG39mXE8qVcYs1KnHVqnA3QJJlLUzGMjC8FywXZOe01tbr9
DgK3s+kWoeCgJGY/xwaoTYLaTnNu+T6mOteN5+ZWOjQ8OxmPOLAmAWW/20aIMX5pYFBVLki+eBoX
ld9zyGgfnup1a30xR7EaF0L8V+bnjf1PQjPH8s+FLdJmepnlroP2w7kSBZVjcMnPrnC3/GEQuGEU
3odOgSUVuFFiN1Q5kgoy9Qbj1X/ikXjvLCeO9/dRWIupBTAZdvr5elfzZf7ENmUrl+OiseA3EAr9
Xy9FDe5yg0nNxvH/WCqmKzjmoyKelaQAU6IXO+fj2niF7CMAjkddl+61G4+jX2YVZn9XtMAu1ly7
CaZTmezl7iQtup5IIwH4u0Vz0MrqxWSDvRgpnQQMR254H15Qk0SV+cz/0kXY5Q4LZRv9+aCr1AIp
cGshz7AvgiIkFJC3R0BF4B0HrfQ4lQZY8BkOC7jjQqTHQ7Qlc/Bv/Fji9Oa8RNV6XQf4XiNK5rYk
qMSSYZbeiyXUcXbUShssSlBVLh+vNGOUFn2QXqhbmai+LZKMz04VCLLFmko9dLsCiaTYHlFyExXD
U//JS3woA1PaOArOGzErxXU0fESk2aPiKT4mUgUhELtb9Xf2bHiJfrQWOupC2YO44jxyy4q/zA2T
0+UFFDYn6ZzWdvMGWKyRsR5w89RmRN4uWiRGKElSbvFfA5LyEqONvPDgqlZUWtRVKbimPcPgInAy
gY3RKcdb851DwAHO2eav1a46Ob+0w7XiWQqolp2YHpA+mi08J/P6sjHThX1EjnkomvJSG1s7LOnX
RQ+GZyZekCgL9luOULhz9WjT/Wxq1SHo2BiDyDx5JRh43YtJpH2G4iesTZGpeElpfl3YIQezhuR7
7CoqiHxKAFRmt5NEnRxxm33VXVNn5RVvmNpF/clLycl+m01FAE6XSawHWLyfm5ssoxGoFhd30VZ+
9SCKFLCNn1KAhq5wL1s/DV2mnzjCQeigWZy2OjsXulSclRirS+HCd8qDHrL25lwu3Um6vX30r0Km
xqieFzLrcKXd/4lQKVuCybw0DrlvrBId3W2H8tDCsZEyqrh19YHqD4NZjonZDMK8mgl1jJR7+Ybh
z8gx/Jpv5uAEM2sXtn8rPkJOsVhurk6Ssi2u1k2sSgZTm/z2eXXmNIjzdR5Q4izndSe1wemuktxT
Q623lzFCipSCUAXDls7jRR+0/Lh3ksXYalY+1PbyaHieEevn75lQ54nLc+ddwM0AvMqzxZ0VtWuX
Vtg0gnAETR+L+tHC7ISnTAS3j4UNnPwCgtNqB5+DdmQrtnU6Wfz2qf9nzQS/dFU4sCP1td5oebDj
bY60BWjCIf8b8FTIzAS6IVMRBuBuRejY/LOMplsG15U8REDg4ZO/XbHZymCZooYAFANRhF+dl7ay
PcamzJDlHwZZntE3L4wh3tnfDD5adDQO/rlExB9W/TV1aL3AE+LN755CW4dFhuG1idBPTz9qtSsl
swjiMtKFY1A7h1IxpTMPSJuPdNLzjHTtNk+MA5A5XaorTmn3RmeebXAa/4MWl5nHIUFCkftJ8H6c
2sfXBfOg60f16HZRvW0Ve0vh2UG3L7yos0rSlOa4TVdRtQUt8KVkrLzQofHcfLB5dy9ZhvptPjSF
4tyoKLS1wPzQTXA7srhWNwllbQOZ1E/Lo9uU76fA3+NxRRNBFUTQ37n9lEkxkmPkPCJLxezcDTe2
AdS5i7Y87lxIl9d/f2rE5wwQA6b6T4ZHMnVll3wIzxROjAvoFODYoMb02+EJJEdHD5qhxXGCg+Iq
qfRnV0jnmJrsUSP1qtwjxvGqZ3lPcKIe9csPS4/DBgZDJl1h6dmbrYrvHe1n5Z+ynCaXOl5j8ik9
RYw3neymmBjUqSjkhVVY3HAndIrinEmGlDmJsiHF7FQzMulUjMk44z6NrqvJtJ6ZJropzFfNdWVz
kS8wmyOsKk45515cRCFn7zl6C23FJvZAZdAAJr04RD8BCWZT7kdWwPk89GryCGq+DjaUblRuXQpj
QZrNH05oKHsYVrpgoW6c22p8hQ+RQ1BYZ7NbQs6/dNYg8KtlCpUULGDfVlrLtNLukkog00AJu5bU
Y9rOerXeiKtG7s0dxQZ/mAP+LFVgAFZD+mDI9iiUjgEF0P6gwn6nEYaIi643e2jH0mdXYjXB5aD6
Fmehuc21bB/VgY4SwGTQ2BckbS1SvW8ftm1lEvzvwWVWTXvlH1XsRYXkQSdJ3Vxc5K3N+q6UIDsT
kwljZEIGzPiBjaScK2VIwui85W30CZcLj/J9C1YUhvAeOxSZbM+w/9ddmiWU6J8WxgDPjIY8BXcm
IEvuZkIXYuxojj6XmUzT5I+rexL7HKLUxRvhGDhSkJE5Uftj2Lf+J4w6auXWyprcZJtgYFLQo8UT
S6YsxnrF8acczQK/Zgfw6JRcTKgYf14vb95w2E6yUzkIgJUPBw1Qzw18T/eJChKh0ke+BsgXjRLC
3LPWh0NfFe1lMzUYyNs9vFB27N0bvTcNFyvnMGhR0BLxloLUqdF8BMkx/N/JD4fmefh9ecKt8RKz
xNdo4n8ZSfqApUe5mcoBMtJueQRqVkLoQsx1WFeMrwJ1WhfmaOkC78XbY5GPrMECR6AoH+Kj0Ac3
74mQkDx9jWV0aNDQV+103a01cLZdMBwAElCA+tf1p2DcEiEZg1IndEjHBFDp39KTJZiNwb4ykGhf
3QPnFMsLSFwHgmcKZvzI9kECynH/ti1retCr3QHsHTm8DKFe+4LfVdzi2mZb2CSnwDkdEO7f+cnL
J01HXZ5JKU62vBJkkcHO1XY8NenKOTcnrZg/oC/WlMXg4mWjnHF9AdRfXDqS0IdHXnmO+TuqiBsE
XyYJZVWBKexUwnudX9doN9z3rRo7pUrvbQemRXZQQg0OzgegzupWfBGFdlJ+0/+/5j7PuQ+8bgO+
M3LlRvOiq1sizfxZN65d6j1bA+DRmeCmYkkt7qlB5kI3CA4Dsrtzju16XMzzQxsWJHtnstT2Blj2
lhbQuGtojoXhDlVwlE5OzWpbWIrhrOVB853a5nNVO0ipzQrRoEcmgs2YIN3gUaeUmJDIXr4OtJR/
dlGxlpQ+C4SwgdlyqvpYD+LRNjlQkSlE1wv8p8Y13zGnkzXA2cgq/4NC/z1OIG+SFwgRq7a6J4fq
DXdgEhY2V7+7GvMcxMgq/TIVtszjEdBqN3kdhPVNkb15b5Za8l+eafwLHYr7XA/GGai7kLVD2wAP
JZCI4qf/V8s8No2oKWu/KgfW1y2GJu8yFIw5u3/JsLAO7a9PklCunh2V2LIfcdynC8QBtb0+CPnw
ecp3qfOcRGThUCRoST9bZePiW4vk6lYqEB1k1gXtbQyCsQ9/EvWkRi9z27TPeepDMHj8qWY1FYDS
BN1qUMd8zIumy1AwQs0RLAQ6T46qJHtRdA2yqWLdDQhb6iNgSY4DRSrC6CQIQfUoHDSypMKgl1Oi
dUgBTz1LEF3rmeJ0/nn9u2jdqFgHD5P8g8O1UDojTzeXveSZgzujIvej2rrt22zPmYtgtmvGNj3V
DZMvakomzNtIp5+FA3+Jp3Vof5T7s13LcIk/j2pLf37sTdNa/78TS8jyQo0GZf3WWSDkCQ44djU5
SukeOFCFfaO2KL7qcuajPgN2pjgsN5uUKu0AOdUfxACdpxXCud3Qn9SVrKUf9Nt5X3iLJN5wHEXc
0wj+rn28B9C3+p9VGPpJIGjjwH17edX4pd6RCESqOCc9To24F7CxSKeMxrNOdP19uZ993i75BCfz
0mzOSp4YjQ54dllNDsDXWgXllYyE+PyvCVqsQRksMFhMIIMjRgEWezwc8TWE+ChPKFDyvC5wjcKe
zouNJaiBI27+UmDkL3NMy3zpsQdFh7xyO6rWVINr1GNk7kq32MRUYY8VHwSVBDXPZS//QmLNys35
zUfeiWdl7e38KYcNIi8iRx6qy4RpVQ2blTcyD5BQb/L/u+jtlujv58DHWMv5CIFWYrXu7lY9fX4Z
OHbWN42Tj5IWwrhT8MJa0weAfhlEk5kU6a1Uoz2e6MBtmazXzkyqUELXKA450lslcyy6SEOx62f0
TAB1W08thlty4CBLUVqMphbvy9UqLUdw0K9Jw7fE3QEtM27i5UmOJbM2O6vuNo+p/9RwmgtEtYlB
biIfGWYrDARXEIYIp2fuW/nvxvbq6E7iLqttBNzBazWisXWcYzG03xrsywWSR4YontUrRi2YwICS
43Vu9KZCw4ilRtPGYNt7MLixgf1rj8QxhBH3nJqs8mw7mrtgb/cb/4c89Eerv7Zud3tb0AEHKCCu
+goezLGYHMvqx3KSh2KWro/czt9iQRYbRMguUCjdseAZBcluDwbULiRlmt1dc4rJcfjKfJ/iHhV/
y7m5e7U1HjSmtNEahHWXpkmZDkNKoKyebS+SXDHr1OObiMgJFoEBg4FE3JmECm6Cvf3jxgzRnKin
Ww9mUAI70KiAG+MTt5eP2ZLXO9ocNveCvszZbxRdwrvMX85YSr4Ue3RG4z5VhG3Dx2VX9AEnY/8h
17EZhN7lBKo8utX2dxGJWEo3J5rZ5VgT3OIyA6nuZxdEo9lKDSrc82CiRLbtdVsV2Jcur60GSoVD
qD5i5sMfBZBfbn9ACZTEVlIrBGREiwCqWeaI6P97NA+yOh03ejSGm8jACFb43MnsBqc4B9bPyNKO
08xGGsLTIQ3rWoAuv5BWx8uLLK0jgMJknOjTrqWRaHjPm0I/HYzFiiq0tues37xILckPcZm4b9tk
FR0OfaW5Q/Xh4hP2T4wfYIPbVMDeFE5NEjTga3xz91RYibpO6KhZNHyNVnXYZ8xIcX7DxGN/VsOa
UokjKqulCxD6cvoh9PcDMj/Tv2SilM7RdYxdILLeYRHchxtS//iWFmnicsaeSsxsugw82VEjs675
dFEWGeyYtNCztE1+a3rPFuvmsE46fLHEZORd+Hp3e73qtBeH/+bwjleCY1A3AktbgoS8fBRN0cj5
mJ/aJBd0/icgTg1QVIKH9s+xIqnABmxSprs4lslRFqrVLqD/QpLghfjeXb6uXeGi61HdlsOnNfOH
y72P6GR8MBWR7TQpU5GLVT1PMRNv4CVMo7hYmCCxIDvn+z6jrLP2O6JbB8jU9dDFadGodsEnrxbp
ZIEeHnDHIIveBTJNf6Os7q5XW+D1UFMwsrrOdHiWZQOWYi3AloyZSL+M5GIPhfbQBgW83OgGL2m6
oUZDDqO4c03at6a08FHhIKtzcE71SBt5mBsv3LhefX7lxaStWxYBqQOvPvApbvxnj5KsGcMzoeY1
9gYNfCwFEFw57+raySgLTGHoH/YZJTNc5pqEh0hqSx5zJ176iBGdPVezGWx5N48GEdjmbPHwr/24
l+RYwqQHu5747hVNblJdaW3MAnC5qy72JaMECPcqGmLVANViQ3NtgRAKCs/GS+Iv+4s1BtDgaoTO
gfXN1bmnHO9hBDpjSclZhwfZ79SQ3klPRAQEeRZ9vRsYKwKwh7DZPM7BZFfQAYQq6eABCIRyxjmg
mtY8R22CRAGv6CP/IH7n3fZGYTTmyZ6kdROjc1X0W+3E9pSyKVDQ31n5uo6rUs1vB8HZMqA71o0Y
NC8ydApCXOpOjqntOU7mgGLXTwYXjxjpweZMZ6b2XrnOtKPdUjPcCzvTWVPfim++fHMqk6SCyc0q
tzRkIPdsdHbX3Th2vK1BtOZQi4cR3NBlfZkqCccX9s1pE3T1/agQZ+Uj+w06aB3No4HacHD8aSW7
eFV/UC7cpWrEvRfo49qrOnv9bJ1xLBCruahdZDtdi3Pzfrsmu8inaBuRsb5da9bwV/hze9hJmEKf
Si4AnUDgixLiZDB1AiweAkBtrDOfADEC/z+ptnch4UDGRkUoxb6GifZAdmLkaEVI8Ki9eYJ1hz0l
yQMc0xCy8/r3e2d4gFbgQDzAgpn9ulH0IAAD+f6Hgh5PyPNrXhyCRa3en+kG31uaNHZ4EWfbLRh7
z4DfFjADb3WT16YZRY3bKPWrlKIRIyI3oNnEZZzv0HH4Kl9rwGcbOy2oXDIekycxut4ZFdEOax3z
QLhKGNWEX1lEn7pH1wE2Xwgk2bJ3mekEDyADb9qb+rcYwywW6eXJDW/x9ftkXBeQaRqpVt9WYplp
bmCZGjRLyIa8glpQufgKoB/GHMnqCGZf6ee+Kd6GsJVEJGkyrP6nRPV6vhd+SY2ahVRM2jHbNKHZ
wLrkqNSi4YnotzzS/0+LtbhRtVpi7eA0/1EX6Uo1JdJklZlfWzfN6Wvbuxt7UTDvrcmyiuMGCV+V
o4vPbRZZ/GL3k03KfA8POFHnKm9Y3fa+FUIz3v7/DOQjO5rny7FJTwQysw5USS98Zh9YyAIgESbW
IiBvAbFkoXolLLc2AQv+d3JL8zTHwuWGXNDsT7ZIE6OXZ6q1619QacSxr3mK7BcBSi6B/DjI0OTc
BnldsTS9BsTAEvIXSLQiyYhsl1DcrZZkMCeDTmq4yVvMWwFu3y+tkIs1NuBZG/xj+z6jcRYYa4J4
JGwzrAP/y+sAFpOLLZPsCsQ8LGdawP9aOo48gbX9r5PjkoN+P9RqvVXqyC/tmdPq5jdlaTuZb6gu
bQyENiwiwQNb8BroCiaqEFivK1Uz4wXr70VZF7CLXbSaD0ibZdxDIkVVsUC1/Gjviw9+sjKMONk8
W7qkMZZ6/RfUWgngYMF1N+4XRxgkZvIVRzkhoYajEEEb6UfnxQXhoyFRzXScDth07+cOkBN7Czdn
8Xx52d4poUjclm+RvNlg/SaJiZZjRs9HX1lSFCa5otSAllckiwlvZaPvuDEYOawASHdOEJ48EEI6
NnNpqraXsofX7EycVMduO7/JG5yYFf6ChpkZH8k3jka12/Kfx2F2F03NJuaKEMwPDoM2H/iNsRvv
S0M78eUk309vMGf3YWxxV2v4dK8ZsVIgPZBG0T7Z5RpqmpDdP5Elq3RNNGlEni7/zyW6w668S9pf
rgWaQI6Otce5PVW0jy5F6SYWgzrnZzVvtsZYGJ0MWCQmurmmVOjDntNNQMpv99/pbgHClKSyQINq
50Tyrrh7AIgOP+Ha/RJBcVv316BnSIS3DmpprDcwe5IvIMvlRAZr9lTp5XMABzcXvkWFHO+EKCgW
ESPMqlXk91ijlFoi5OkCVJ9hUAnIetvF7Z3nHHhKEY2haCf4qlNNAZiZcW77CGS/cLD/AniUziuD
pvFZ9EPPDSZau0WTmYbHjmXvZ9497mBV6XPJYrA8IiO6sfzQV42uaB+ob7JjbXHpdGIfUz4+hIbt
wikt5WOEbKczqbiiyaekutKM1fyIWXMXsO+EYI19ndUxZhOmRpLtR3qBz0iczeW5KY5nMyK7scip
xk3XHhXOLkGrIWA0BhujuUPPNwqRB4HguBPi8DU2JsU8iVKygtiVQ4Ahx2b9dqGUAE0Mc70U4FYY
VEB2uKZO51DWoBO5Ux082ZHvkXnM3/Em+2TVSFEqVt/y3UHTZJg+FjPegejm6WAIvdULftE8kcNo
stmJLXQVb2T5I/TKgTzNJniQSsfp1P9sL8y556bhcnJrN4JzY35c3Hj8Ix+0SW3xlFuHyNMuWRG6
4kTg8nV6j/+QEsubphBojMmH2xrs/D4uZyx7THSSCyFCoPXwJ/Dsu78QROpXOxi597aSHv9dlCbk
Wu4zjza5CJIW+GBfvDZM1UWt8sH4eTuEdyYy4/cUdYRGftzQLFreato/24iByNQM+BvIGG8vdvLH
sy64i2E5XlubZyGstkgagdsb0VJTyJncocm+6a4BOpoGw4s6/OD+xsWivgNe1Ov5k+drwaWcjgbD
DN6pv1CXeO6bv63h26Ld0deiYAcDQFuvAkwWOFaj+NFekqGa/c0n599RAm6XJ0dTdYA28fK09Smc
vhLcsLo6sFaPG4cRzlbLf3ZYcYWpdEIask9g2djR9vVrZ9eCoXhSSHK1LKDfD5GN2k+vy3XbU9jg
3iRrAlIPlS00xLku2oJ9CXtDW8S+Exu1jSYUc/SE5pZgmbaHJ/Yma7HN8xSRy90sntgU/BT1RflB
XDdLlCroszdDCsPD97nPIKUfdpa1029P+67OsMTpWnxANx/RRE3c6f1sOCGzkKho/ezucDfy/jMK
8I5Qd8UW/QpGNWJvKVXEc3udh62MFtSn5V6zGr6gwxVaJaDA291ZRW4dMuu33u+hJjFYcqzuRAZ3
o3lIA8e7mDlvoQ88RT/F73DUKnYCAl2awC/gM+h01h4ddjLkUlFNxII27Ab2KCvmtObfaQZCVIwN
Qz4NbgVFJYM0VgXQDrJc6gYz8aepbfMAD9hw1/0CVj4P8ST+3emMe0enAd6qZkWJfVTV+bsgbQlQ
0RW/CdLKyq+QslQYRakVXgjUfNs3iFftf/uP5khGwseHoc3mYE+OdVr/9hRawvvWAzAC5t00jZEz
w1wRaOF30rHDNdvue+UpaFUO5tqOzRuattL+5wDDjauCqo2vGTkUJ0dTZO9MObaCs3z3ood562Gc
sD9gswaq0Bjto5Hc0tjyeH6sh9pBCO2yvg9Os/LB3+3J4Vjun+cMJavy5Cxgtsw6lKGRkZCnznap
ceXmKgQUc8BpuRpCF23XbcYjqRusR9RNab7YZt+y24BrSdmNI+1YWw+bBAIbNJ3vLXeKY8+cfbrA
MYl6JFU2TS0fkfP4tSzwkE7JmzGMetUP/3BwfqHMYcpjjkJFXECO6Ec3lboNOg/Wc4nB79G/w5zF
J3zxms517oc+gkk8V2xHXO+4QiagQtXGE5Am4PvsEXB89wMAzMWnxx55OhU0Q1z2/C3EuR0tB6b1
GLb2QTJB650jiI9NatwlXsj52b/bT266illnYxczD4HaA/yaDx4tiSPwsJ32kdsy2ZxBS6jHAxSG
Z/7vWpfMDs1wzvu8GjPoxqh/6EweconKupiFY5ok7fdqmCkuT/PsCUp8BYwokl5uUV84EKr/0U+0
5viF6UAAyka2H4NYU0WsCXv+lzgPpuJP+6k1anmuSUfRR2st2OZHFoF6Le3XnO/JQfGDlsS9JfWb
ZRX48Vbm1do5xGoBrXtFi1hUaxHivb2ma1SCxAuGKwKP9E5lItV4gy+9IC7Vgm30uZ7IkxCiF+Ya
g/9wi+aIkFj6s3zVVPq5jMBEpk4M46+rsFq6aMh/QUu87NpwveVuNdQWaXAg+dyfnP6mpPlsBOpB
I6SkboS40qDi952iqwnk80E4xq1agIRJUTvKLOjQwrY2/hYH8JCcBrnz20x4PNwnIbh1SvhbDFBR
49w9TcZBnB72hfI9XMvxFtWIKQrdG0GiimkCW1WT9Sffe6TBiBOqoLK3puAd8XjWJoZlBDVmy1cs
UbxfAZN6V/6mQ3E9UjKJgOIlfZ0EdeLbGIKUrotAS23wJ3PNzC2k2EJV03/yGq6bO+ZmBaRGbXAS
rExpVaM4gFa/r/tFBNs2T0iWOKKv4hUrhCPizqjOvHE3/np8RLk2vBGgjOFOpeDxYpDFO1nw2yhs
QGn63cOmdaaSOFvVTbjaAGV8gEQZ95RBZrACRdmXUPK2sfcVBJp0BdiPpdXj5sVFu1+mG3eXAAR4
HgYdnhqTQT1fwmZNklUN7a6G4g9n2zLkXroG7Ez3onb4EuOle74u+pG5EzKaMt+3HDqccVJXOhnN
X4apm6rCqhJP1FbeDKSm3ti2Y+vHNQCyYtnDdpmCd1ucouXp80UgFUifZRdz4oRlb9fS3JsD0ZeV
QG4mv4QjrDj2LmtiWiBz1L4zCGCjLnayrR8/9kMrIJtxjb4R3OMO95H8Io9WB/1wjPBznGy3jlce
JdfvOzleuCvwANXhCmv1/pCqdb85Im4pf52Im0S5HyDKTthOHvW4673T4ll6GMMLlL44Jewx310f
W3HCzOyQQFQciW1jAUqUjPyLWuMCRL8e4AVovdrJ2Gzj/0mrrUmU2/MS2HsCoQOE6Ye3l/D2G9zJ
BDlaoiq52lLwgf5FH8KpCoPuTo1BLxkBO/uz2MHcavfqJMqVCwSsolH/Lh5HAGv6dPTdGAiZNsc1
wxDhDaUDdN0d0MxN1ow7ihDptrBzUynZhJvXFhgsm1krrG6bpgB7H9fguW8SCA/kKsNX6bNmx3ej
qMc+eywuIMCqKAhBx985vgzh+wQqjJQXlCBCRBm0eQM5LrsKspydR25AyrZhC6SeZtYtF5n8CdDd
GMtsLal7NMJF1dQzMrZIOB+kAOGZl23xqh5GdtQBX8PIKLf+sMEXcM9fseE1mCFG9l9JhvT+nD19
xWv2Fie2PBqjsFuYx7GIbY/sjs9vy//4ZVLzFAIY1b1ubna9HZMeJN26TqHGqWDjFXOlQzPzz/19
3CkhdxK6VMKHtQQjRW0l2NXkGoMuD1uCGb9fIOmxZErfBufV04vh1IFBgytLssIl+/myDVxI3hVL
wEE0UOAtIo+mIZpo+5eU/EC0P7XTdRwIZzOxHD8ONC0kp05Mge72NgKVajk0fmu6awjl5dUg1oxD
XEE6fdjxGfCKgXtMQ6g/aAb9xFzOF6iuAulR8rfNCLwSKJlkqgsBu3mWlCL8M+ScvxDQtn4NS7d8
FRWFFG9UcZxKqfxdDIRr/zH4XAfUfHtgNvwXL7JtUI+kLE/IhMAekxKZPKoEM2NexKSFv6jhudzo
UF+v5FLZjn1fj/VSviLxzyG/DQFGDTXTjre2NyHpmEehAqwzLobZu5kfVBPzM7C7xEM1tH330ZHU
UqFz2F8b9vsHEkrS4bKPP+3Iu1H/sispUPHysGUf/ux8P8AThVCVe2jnXmpu9k310KTOghztwRtI
IsgYJ7CQcScLbvOQbroyZ5c4ZtMV9zLsLAbP1g6rM+ft0PcNR/zN4jxo7zIBIUGznao4XfTedqll
AcRHkr6XkXgdWsa6QSGUGlqT7x4k6d2Z8Mzr8xdlBUNHeq0O4gOi9tsMZdl1hKqgNnK8qT3ZLboA
pCUQEE3EXtfSjrbl9XriHZWzffxtX/XOjYh0x9Dnaa4BqB1dKMHQT8COqotT66DdWyYr+7cw4Uj/
9wN1YU+IktL1dbF3sO9kRVyhjcgNXuuDdhITmge74mwoOVAVHBQcgJMYtkjUq7H+LJPNYFH4OhvV
mB9EFewGVXprxlnk7PByU0JRmEsHiqlVkQUWB64PQ+ANojc+XHcEo2mQNMlU0H4gowPqefHV6A5Y
LkOCJ28xdgeqIRKKsCl404J0f7EN3jM8+TimG+E8flzLGH12B7SlAI6Cx5GZEfKFyvh6gA9jthIv
BB/NyQsMF8KI/gM8LTj9cMbMqdITk9y77vYkheUp1dCvxHGuID6PeKrcEHaMe9eBuu5DMRUJnG6a
c1n8d74is4nDAQKQKtIk5KXKxFD1QWj0cRnSA7k+OypF1KRK34/CrFjoobk80CI/tSouXeKefe2g
XV5un1E3O51jP0Qa4sqCfcO88e9I8c2lfiP+0t5FRVBEDnlcy2WLjYWh3+R/GQ6sgfpyZdMn9kiD
8Aze7r7pRclw0W6NLghIt1LsjzVKqsBqwwhHvAjSfs3HpuD0mTq18TvxDu9VtSMsrxtR6ELZFY0+
tevP+Bm91smUtRqXvOsDMc5rcvBoeOf9kT3SICs6/LW+3xm7eL+AJmFQct9LO2tqPMSEq2pk6APw
CnyVIln0kYxe2D1S+OlyyH+ljY6v/0cr3NNxjTCgRKJNQqWmh5iNLonFgsnoV98QQvIYtVkbssrG
GxtvDMnw/M7tzxnLhMp5NUGN98s6K2E0Blk5YMxcdhRZJJCGnYEqf3mImTQ4yZNqV0N2SOSgMpif
5TbpIgdoPnD98SQoTErPDv0dz51Ba3G4qXD10+Tj3+A0nl4LTM8F3p6fWMNCavKQ6wvpO0k9Qrb6
NG6sKaZX8Kh+MTw5IN+UlX/U23r53dk4squwKAtpxKe6+pjnCTDeWiumgGD6VIQA0LZDCnTY8eyS
WBrdxo8ux8MHwFopZ4VEPwaCNv2QSPuTj09BTVk69mFkT4qyRQZ1NTGjMV87hl6lIks8TJqz27GB
jPZNK1tVz5/kFE/O5AbyZcePnrCNpaeez6kiLuU+udhwTLHWjWjSERknXmBjXdAsAJIZK0XB7pr8
ViMXpHE6NUHG3r6a06h5cw/d+TnaiWYd4rxZg96sBy91lpm7WQMDmeGsZWVqXw0LzluD3Ft1bPGW
NSsKse+FlRogo2MLhP2RGYnpQsT6pFfClxLlaftVEjwUnYHN8qq68WmzkIEQMepDLcWV8l4raEX1
uyE/hcYZZSDCU/oom0J9G93vrRmkaG3/hzCHwZUT0gLahB3Xr0yOuScyMfqJuHS/SM1JI8FDxGYj
HZC0hItqqvSA7GsirFS4VxM9ABUrDv4VmPuq6IgpjPFA+rkrh3MMM75r7oUfZ/hVpwbz0TjRsjzE
B0nt5yNh+H/cFBLeBfw5zUpUhq6TFEbftBDgJW0ouA2OKBY+xp6od1sj0lp6s/jDPoGElXuBwC25
zq6QWUwrVofdBzHyrnwduehan1guHzS1jHDeqRB+X3sWczNxKgubXJtsej1uR+CvFdv2BZMHKkz7
jzg8qMnrfQ7W0v8kHGGWMdfpDcSSKrwIKjcE+OoGmD+O3CVAj/Cr8O8uN5qJ8AyA14y9hy6d5y+p
un21+nmLHGh4ZLDv7ec3eR1RM7ooetB3g3jZTjqeyJSxLUkFF2YYIYrgOlUdSIuHB5hhhDPU9Liv
YmOWujHqiQ9v3JbcOeYnrngsUTkQsbyRa7SMc0phDFZ+7sIiWQYWQ9d1hgcQVDbdi8kdGyVCvP7/
w+j0xlV4nYJApdQO5xwKBps2aMo78MxmJJBmLLmrgdUix+8mZYHGgjokYWFRWnTsBatfL9jxtReE
D1ryP/z9DbRdeWY+8Px8HEIdnPuMbwhaz0O8TpSlk3UxVO9Cf/UunFth+DttFEhSKkvhz8LfvbGb
WlvBgC6FnvPeZ34pkCO2uAWul45SJPm7vcg/OgTzTLYaibHtjrW4R9ztlWJHKfYJqsLSR8zez2lf
sqO0vB4alNk4HbKcwsvnHxHFrJoiKoh22JBvtc2FMPbQIEEhihGMrGq4XEtmWKFmfrNxbvPhICaI
9Kf9YpVn3uG/b0+mp5hcNNjt7rQLZCWGGUYYK7obVusg7KaKDN55SoQb0g4kCHPXe3sly5QZBcH8
Hg2tCt7Vm7pPmtP6+20KSKw7ExrmiygXz8mI5PI+kxxy/u9KlsD80UmZdbWIWWbr6gD5nOcSiCpD
/DTpjHNu1TnGbJNMVPaPTAYwElFxwIbOW20LGtW+zyU+HXGbTnTB6abru+pJs4KuPwzEKQ6Q29bi
5cr9sKe5xy7bGYQzVsYwK0KtMC3rfWUwAawa0wHrMBKUVuXDI/O5usLUp9mWQPoJU+19TZuQX952
+BIlgxc4VbezvMp/2Y+P392vZXg5cFGyBqVfjOe8DFNBKMVVll985gvEUUicjD25kHtYQOgX974j
QaRpzffD9AK2tILH6OYXtdkCQ6ZrIY2zz65L7j8NJiowBhotNsVoTsaCWVzKm/2O/+wRoQkURqb1
xo6pVC9LlidKravuWqrROhhNLxlcDFkbmwk7J8LEK1LOtsAtEgHoiyzu0uLjt3Qg+iL4XHx8F/ww
EB09ARLsDrCu/jBFKh07ClMnfKbgCWMK1HK8Q2LREsokcl1gHLm4HGTW1pNLd7MyDmM5aTwRDcYr
vbm6VrHSkeRfcRmfHqcW8exOqTXo+1j7uPy2kr/pGRY7W3lUjMUZMiy0OkGVN/mgDGOyutyWYkeX
NhvCuPrQZ1r1IiPWWGhDAE4FX0+6x5iy589RiA/mdgzYJzdZTmTVDdBsElDS7+WfYkR2h9D+hi0h
Eox536q/R2p4aNlEKxlOILFFHuF1p2PfHWYNwkfxPuHHen2yEpCyA93aje4z+OaIALvafiKmIozv
NXJ4zo9YPeF/b8K+X+bSwL7YDGIk3tf/RUK4GEYDeiojeLsZ7zqogZyMZsL27j62/Bus7s8F/h8C
0jWGzb4U77g/2liKVzUH3KZ/Z4MvV0LV7YJHAyeVc/9ZgJ01lnWS5D3xDM7WycyoZmKf86XM3eeB
qYLFRLMYgt00PCjwfnX2KmQeEWpOhbgrHWHeKe0RZrWaZf7YckQ1sTpm+2B2HhJ8sb8y3Uq4GBRg
fGBBcTyp8PlRZHcqVvxEKRPBLmwcBUR8wFqcU6gRmhloce47P0BdubXgU1un2ks7pY4yebOzP0Jw
54MhXztAvgthsyJhXggliozKmaWc7/c3N6bG1tMww6ih2i9PDQdEWy8UspYfRQc3HsJ0vlamLD9q
kMYrHmE9voCwMAeFxyi2utAqHQY3xuWYvLBb9Nrubsa+Gv7Pl4gtsXDnAuLKFs+OwEJ5YiUcnFXg
iZN/PLgQ++GeODHavP+6AE/qthD649b6akU00btTOe6a20tobhq0y0h3dEZDcrlHfVFHFmI8Lz2Y
xPV4pja4r5T7zKH0d14DgZ0h7HdOxY3w+X65yGbtFBbKy0xKD0ZIBjzvoKc8DXtqowV3Dol7QOFd
UQFVWxdL3uSvIQ1aplyN9TPf3F4q9ATd9NSamBOUJUtUlc60DxaW8emaDMij2RNKzjMLo21TPywh
nmzq2wMmLrVJn8eKBXfkJw/DnHUT6u4beSt4fyOyPNOXK4r8zVXK3r2S+9iVZx+M4LqT+P4nmYdA
eTmZE8puKwiI9GECFliZQ7WgWiXLmk4ERYtgonsg8ADfT+plwS19S3T5CZAS8UyVN76MAl1A+syi
VEGxdKDKPfEj7f4eBgEJh/59E3gXQmJVahTWYIGtuVNra7e4dI4lEVTRK3njPOc85qWxFgffRAla
C03FBmKr9S/4iVatXzWsKmTh08Pa90ACBEIo1EgaYh4t/2eYPI/fsVkaqVmmZKxdBElPW9in2I69
mNYwweauJMHuf1z1PDRN5NUw8irjwupS2iHkEiJf4RXjlWcHioDITFE9fWuulls3HWHX+7nZMqUc
0WFSSncCFqqTc76pbrWnA5nwC3/Bq3XmsyHlmOpvVhkKexEcTLBgwL1sm7PC7kLed9oCwiRt+ZFS
ofUie1+mSQtRfP9RWFgmyVT6BxztadGX7oe/07ZG+U4C37jFc/7baxXNtijcNE3EWeURIktnIcmr
0FcBsr/w1lS8+5Pw/SjcJNoOm04UVpzyRL/lrMXMsGg8++qASzNFynd779gx1lZ34ETHk5wFdOfB
Rj/97VnX5Kf4O1knv0Ao2EgDnST0+DBq3IMwBPRDvPVMypyNlkCyzmOcx/gzNgBTV4cMgaDviWch
3mM2qWqqRlDWFWXSN+OuYkWvMtkjhaQHvMJeQ3JoAxpLTRZFuTvOnmGJl5jtEgiyrK3k/LRbU7Mf
lExBPb1Hlv/pcqnAXG0OZPmyLQ0zt5wwzDZMTWq8S2F0CgDny68rXAiGha7y45ZYyQEPlpsHu9qc
htgckhMo/mErSo5oCgXUzkl0YCEjYRKa2HJLY1PrnP58izI0J9rADwjNd1o3yHLjDVZuHiK0WlOj
LWMxeYbrCE+AJMt2MciE2MfCsOk4NhjdYMI4j6voUDiwRf3h85H6olRBl0iGQnfaNg0vKQz/9sz6
7LvuwbOw9SraViPIonZ68HhJ/OEEJNSh8qQlawXwHERcix7VAobR6RsmzfwcKg71fBEP/Z+Cegcv
E9azB1osfQUQ2LEhYIH+Pa9qzvJf+MCrFHDoX/dlJprLj/2jsQghoibfkBEAoQ/JJrTAb08N7/lV
hIyLaRjMbHaHuCYCEeTTlby2IRlFZdDq+q3YIuiQDCUVRin2rrymiiF1vYBfKsWZD/icppePGEmZ
ok+fm6Y2smVHniZM7953AwtcRCSfLvsCoCAsgeWDJIxKSCbU5ivSWBvEs9uF5tYzU9zhM8aqZivV
8GNgDeG/yxW8n95T4DRfgothRwhg0MCzNIKKhJoIompjKUZZAH1GAztD5x8cu7ma4nTDYNTODpI9
yjskyF8N4K97ossIWQ4+8lBACYDeUpgCe1YO/zJCcEr2dm5E9rw0J4ANEPt0rI3JgTI5QuLKlyr/
3MR2h72PMkf8UWdTjyG8JKIeV8b1yQRZ8n+G+D7udO13utNG1gmqMVVdygrJ0IvFVFxi3cmk790q
0+0wdwWPmT0zA+zb0USUJpzGuSBCd8Aum2PCqKYmv9KN1yV5O4oRXVJc8jse/D/sqXL781VyP4vA
OysqqJPFh27pDuvhAmDMPjwYSmSSoSMDCTi0Xoluu+6qMhbwUjjZ9pjQZ17v0fXbbo7dE6QV96dI
L+z4gamu+CUWSL43oZqG/OqZJpGsRYs/23FKyIZM8RUxTOrcKH4YCl6FsmgaawxfXwy90xR9v4On
Jo3mKA9BBGaVOlHbiDMXaq36cWcpgI6M3HJBHHYsIfCAAY2LyavnnM5+ydSup6L/esxOJmh/ktPM
RCKdirNNOSO9hZUX9EI8+k72HMO7eLfbhFkH8OZLMe2THzTj9w5TdH+CHIwZr0B0uOdgdXdGD7j6
88J9DIUGChryfXNIwTsZLPS3yhXyC3qRvlpkvUm+S7d5OhUZrnKzYLQxOl9u8CId2gX2HaBEN1eO
f9s9z4hKEuukMpylMZBL8WA9n4meTH39/0I++l92neuNS+9eJUHPE9JhRMPWyMPDD9dpWIMjfkzO
p4TP168prnb5ymq9n7x5RsqGFs4g7p/FDnRJsXV+h7XhatMfbHrY/WAvZAUx2A0b4cShV3JLoC1B
uzn1OKjAiv9nS32QT673OatUrzK19E/XSVZvsftwglI54aG7nW3X53+p4Kcc2r30HRTiFoFKITGV
50xDC/HILmG2/vfSAU3cYmoTAW4DVLtMnO+HUIwI8PsrZmOi8crw6CRn1z9XZnW6rlTI8qLD99GY
L8Grd603pwIyqv6tG2EdMGe0/TJWwHnBipvLGK53hD0MwBifNbmSczdu3pOaBQ/TuIhy6oDjqCci
a2n0eBK3Tpogcln1+A2o4xS/pK7glYKjLTJFleAv7/z5Zaq2OhkyS2XZsOfjIR1L64jCP35CLSSH
PLyXqg5cA062AHG4z71T1Ia1Da4RkwIepeISwt+lI7DfgBnpxMiXT64Or5lKQST02QzYrr8uiXoK
WaqF49yQfgrFum/jNs948vkTN4+gtfv39ZSqPm2MhWEv60F6c9SJEbKSIFEiV03xQVcSei9fRT/S
7XCB23AlsjaoNIq2BM9DODyxkqpqh5q5MQmRql7M1hUfCWj1QDhLAWmUKXudunukazC1m6PmF794
3gsFvcVwL0wTYFb9g2+V5n6tiqYFOuvNzGauWCDnFscc8NFo4jCfsbs7fy32ZyJAj3G6tnP34FsV
68kxvhcu5CYVBWWrYoPljDFPQJtjKxhLzMItHhr0VnNWcw4yo+qz4sbxZC6ub0NQi9fXMD48tNXp
T4sxSxD2EmIFGlsJYOWxHcaVTlP6LwP3XBjer5vecJo+Za1s1MU9GDaq6sK5stga15J44WXkLDPA
ATf1jTE9OE0plyvEiT7i7QdO9meB0kO0QzVJY2scv+teYlxHecnULTXnTb6u7lf7J0H/dGZwDBKD
ra3/SzFKrtxoEppuGulq1yxvewQguKG0t1wrprQ93jqMMtvycjR8E5ex7mPhKBvYASsG4uxtske8
QdEo1jgyxihUiBgh+KriVkrtbEyVTtH+QR6M+jYVSfz3U/VDFdkpoKhKICK2YHjn7IFz5LMckJUT
ljMBsWHLhqBtrqj37unW0QsBmxoPGGogJ/F74H8SX+FOAa7clM7HpNvMx0RCN6HgzrZeMjx+Y7b5
vJNvsNm96nDhXWhW9MRSSuhFGhR+BN8JKN3XMOug6dL6atXnS+N2GZvoYAGwnmNnFxhHEZUtlgvf
Tr1IOb3+8YGm4ZnsGrYZbKKYbdI6Z4x9gBmdbii4/su5ZGjGWRbRnSK3M9canyLeiU2eQoRUI403
LSPqI4ua1LI2bXAdF0bUVa41Fj1n+l4yWhcmrgovW2yXA+mxnkCuoDBHgjEBQePUcl7IYFV3oFwv
D0rCcYwd0kftLARBepXsj9RjEe7heiRIbWEuiZc5OIcbuwTBRh9wLVV20ijao0adYqav+gxYdwcf
DNiueCwcJ8zev/is1IRUp9vYD8aaSds4TLYA51b5W2G+9FKrWF6kiWUagb24Q1QFFobJb5glV7VJ
uzjjMji1qrMFMJDd0JNg0nzJY4RTHc0lxeOB/0p521M+iy/7sXO4MIEW72E0nggQYqM5Y9Zx+u75
3TnHg8Ts0Cu1CSVWJrYz76Wy3e1RbuuyXVb0mj0il9WCMmva0f7UQsbMBQVPFcQrvBnpNucM6Byg
opTSmH+2PtjSeULVy8w6B5gCnYBF4Ju536R4Vv9YsL42QTbUaGU2zC7HAzOHvpoKA1DYVzr0CR57
nCBsWVaf9SajqMfjV2pS1K+Lt8yv3pzkFEzYPZJfH6v/GZDVtV4PHNyztBLphznQKC6PVonNexcr
Q/FAYRZQ/z1lFiUSspIAbmjDa7NQgsuT+svynAOwBgv2ktUPvni0II+bPYB0kjtXpZb7Z9/LbnD1
YO0qeNQrlDHJVrSumHar7qJKKC1nW7HpWmd75y2Z5+9L87VKaz4pPADe6c9DtxgqYaNB4HXI7F/o
4FRsUzk/GuwRXkDNjDdGcnGLYvcOT7TaCMBEJpFKrlzxJ9Fmx2kEWcWjHKjnkrAiWdMGYJx5XYhO
FsD5kRj7C1at96uX1aYti20PGOGDMAxvRZFlPLzxPbMg18q5O3k6opbNAklQuvRg5Y4jqvHnvU/L
DguD0RTsxAEclFlHRPv4DmFtG6xg9qEjuuyRSoBu6Ae9QX7YJZ5Hyv53+9ZQISaQMQ55eBND/Y/F
VYKOFKTcQIkvHHoDvSt0Wc9y0SSm1zfbClwUk/C4/D76nwrwjddm30GYmbAnrtKrr+ailsFR1/z3
Q+0+MUwsRABK+Tr9UGmJV2pl9Tg3ASH7pQNLEar56wK9KBVbm11cH9+QyLpCMAzfJZD9+UEuyFJ0
s4y8RbRQq+4/9YRNC0zn7LoWql3q54GjXQsmKm2/+niKrh4WgH2hcnDAZ6e59LAwI2mn2UlK3jHG
6pjJL5Bpcz03EaWJAiTi2nK9XrZKYsQpyY/3h4GaYFLh5Rsjonjl1hpGaSE1DqCdobHHsu2KmuLU
kI/VFhDEe6iVRfwrSkhLCHKnKMJKQF3Fl1WuI7GQZopYd0LnqIoi4Jqs/DaNCfoi49uMr+VAlWtC
KdDmVix4lMtSbSYvOhV77f5o3YmKRzR9oqjdC3sn/cXlcHniMVl1WwuxG5A7og7NlvdHcrrbnve1
SA7H08jCV6kcyrZmbbdsiqPibcDoXkEFYp5vKOBaMjzdS/orbTUJRLnz0W3yi0VU+WNCd0NPTsc3
PVwSyKAl7cjbdV37ArhwRDIR6/ET+PXYvZCw5Nvj0OX3jwbQf78xn5ZTlNaYIXrmf+kFu3rGq28f
jsAM33zxyXREDuOiHsgmwv7nNwyg8rayfXVikV4mHGZ6B9Pt49C1rFxzPLdjJiOKR/4JmacxbBu4
8oW5domiPMykGgUJZdSP0tOauIvLVzf7TEQ5ssGZcFqFEbx5CtxYiCPqGwG0pStFUP30fFBN6Quq
tVsXjwN+iKp2hxXI21OH6iqn6Km/oEEFH165OfHTzwrFAOTwfSXLyxD/2QX0jdskeacI6A2QWU9i
G8tPlw79U3kWUTHdrHlY3NeYSDNrXkOHIIVmMLZxG0U09SoQHypEKrconXo30bGGQA3l0UZbqoXY
Qkf8fZc4j6ttinE2B7BdP/DI+jR++hWzxLL8DBOOHKOl00VSL4xvoMFRsgJYsCQiWyAHg9A6BD0A
dG5CghkfSjQoqKQCWWn82xZgKbZBY8vAcpLo4gJEUSbTMRvVdU3ZwMQs/iud49l2MigCC66S9i0U
VPRH3bfzK68N3JrfxZI4nVLbfw1xNddGOmFLEzUYrN7lNACpd7iH1J1gug2gBrzROWUiFAwW54uZ
otPOiFPDGoDY6+jNtXv9LW5P6GucwL2h++orVh+t29hyyyHjeMjUtmJojhj+Dgb9fA3TKJf33gre
QhX6Ub5t3/8NbBw/6zVnCNBr4w18JByNUPW53rlJPtCrGBmrDaECSbfS7qbJLUrOxnR8vdYAJMj4
7TphekCWBZfqdCy2KxQg1hHX5l1cEBGLVMlj+CYPl7KSNH68siRt+Q5PRIfbcGEUZg65/7WFzX3c
R9kkCWvv1FlOYUQhIrrdEjesTRfEz7/JgU2BYtVMrWPFON0zUo3ILwvQI0pDKWW3U4TLN8bHZJtG
ux6X3wws341jvuXjev365/bgz6sodyDcfUtTGjWyBJfwBnLPrFW1OVblfO/dGGjkq0ULwtwdzNQt
jYeeGLKCwGv0Op8eyXdKLPvu7NxY/wnXPvjHMTJN1qDPThWnRRfYO8oi8bNjM5EdXWSopqqHLRET
k7772ggmJvaUIUbq9zMtm9XPjtifflmXAbbq/FKQGK+vIOpeaL6BHFwjDwpcB/BUSlkIYPx4UXKt
WQIBJSiPWddniC2haPBmnNCEczTt/OqZtkzUlL9LfiijbF1/X6uzk1QrQFAmel3oZgbGxnbTCGJX
T+YvnGzj0XlH+LcZ3ZsdQwupujY4NNpkiML6X2fiMURmMXjhoYRcNecLaJlpRwwHV6onz3H0zwUl
PfRR8hDW37Xn/Wo2OQXjoLe3QhFa4s590GedDtACOacrYSIxCaq6evD72DxN7lWP9lqSA6yxd5P6
Ok4oTPRKOXG4srAEMvOm5bjrWnKXpAnQnIYDOoVOavlj8HBU1SL1ts1qEmlv/VGlUrHZ8kXnL0Oc
Cup3/SE116m8j8IKaN7HtJZ3QD97AyzjCaHzjw1kfZFBguoV1Mgq+MJX2KP8cr0MY7vDZ9kuWnzy
iYB3Xlq5p7pdzn9IaKbN4GwRSmSKzijlSV0zl6xwxV20Z0b+8AlhUMnKvF03Px07qQwxT+mSOPJs
ysONQvx/M9KPVQe0LGFyT/t4rmuAJVbC9uN5wDZoSf6elk+PbJT1g6Xsl4cxbFqBTRxL7wOqhvCO
JdaqVpSDT8IVr5O+7rLu7inKt+XGKPDlL48GHLpZGTafJw2cCRRfYaL7Vq3O+RFuA/+FucdKCf2O
oX6He+R2Rx/HsDpEjnHEtCVVI53S8YzPXThEhbVLZ1dAkfb/cIYQ0iG1c4sIPSG8VbX/kTuhxZEn
Pelv47xLx/+Jo7CSM9Oja0tvrTrshFOloCGR/QH8bjbgvrFasLc264OV454YjtYBF9GIVjhvrZQ1
JGkM57vCDxxp/FT/j1QuKc05a/AxtSYR8jeT4Pok/dE+zL93ZtLofoY34Mfg3HKOlDi33dUetEN1
z1RTARyMpC65nHZyckvrdKTB+9lBqm9hVo8o7iZ4c97rIGb05rNFNZT1hLvtWgS/VH3jc4SaSWce
3ug+fSrJfyRSdqnoFwsNBLxrmVBHcD7G4BAD232spvX+nIGbRFvcD9mZn4FCFf4g7RklESMHbaPB
2mu2AtdXQjwonsITPWGnOal5L+z73re+AYPahafXKyCxRwNaPI4eROISInGB9eWWxFyTAOTUTPqq
et3fGeo1FLnCADs3fN0ZrqyLPtjg9FfOEgrXdWrlpPRIEGab2IKBOboIeEJkJHW/HRXlI8zP0W22
UCHV6BuRHA6MrtRsVpvbv5pzz7HmMVzWZ9kPGQhkmgvZ55CUtVsuvcH3H0dykoXcKEbz4mvXiWLX
vh4Dw2mukRIa2Ip1n7msP8cHTYam2BHlrCqFwmhyh32Wd0maNyF12epRcwqSxjAGZZD8WnX/0cLY
Fo5uvkGgQjpPaDJ0E58NfxUsS+XLqOwlk/FriLydAcB/KNVKm7weJRNB7tD8rUihJ+dVIsg3euJv
HCdARtVfcz98PEJfIr0p4TOYSHfPPY31yghq9FblQj2ntGyOUB6ju+qYz9wBPap5w1JwRptZde6q
TNQyJDO/iYZvtg7JPm57WN352Ua4qScf9F4ev13GAbTEqk0XUAL7OMXGhiJjN0+TpIdURMaErwFY
LcnHt266G72LF/o1EcYYPIUrAnsQc97X4YNcVssLl2yQA7gDT4/psgSgDY9Wuo3OJT3QIDgccxFU
P/IStPVkgoP2PVTu9btnefBsjR5t322kHGXW7JrwSveXXaaUs2Ra4Z3Na3K2mI963bZ1mlMTK/OI
uCdagb4N6fiFSAxbONWOcviiBEuOG9Ft8Tkj21MXQUTj3sCTspuGUNE0e8cvdycUd767otUNXm9q
SJaEsHgDIBR9lvq3rd6hq9VXvWOoaCcxwF4Cv1teEyQUDLgWUQ5k+j8Cdk7+gdlr6uusNT7pgt+z
u4lRH5WitcrQAca/yj1djd8r9QZgPpdgQM1qnJzw9dloyXEGtRBxXyOBXkhG7FMX0ZgrLHVD9ATf
H+WV0qaWNf3kuxvsuVwOgPrL0C1TwN2n/o25QQaS0Z+WTnjD00vtF0Pm660va56orHoXO56NvgkC
yPq0WHzDPejVJgF4HKvRpfHtRki56BfL9m8kMWmI1saunAoasTYzLTa/J7tHSk7dgMMNIE531df/
QMdIMzIrTEfWgVYJkzeqZyHegM735t0DrAp3PBx4P04qTxcGS3B0B0rka/XXScE33zvcnAMCk6rR
+fJsEIsABCl2znaKylhfSE6kAPeIL4xCBkzf/jCk+IfRGReaN7lgeqQZHzrpQsyQGiQYUkh+2cNj
oycNBbp840qpbG5/TrG9nAv3fpdSG4j0ym8uDEoTe2WB4bEszA3IvjuokFsQiqI2Fur/yCLLXQwW
k3n4AO+WRV7BpI1WzM3RCYJDc6A5Oyy818YjlOhA/0d1ke1OrrcVY3/XmK0ejVM/x0XSS22qsUw6
VpRX5YJWD+WJphr/PdqbpUvWbxD9maW51ThMyCPBnUuVmXTIShz3KQUOcOgopKZVOnYTtqshn0of
IqBOVmnTWdn5pPSvdM/prsdHMaPZA+xA4BiGosvQ6ndDmcqD1gZ39/AYRT6kvDvBYlGF61rGjXpR
7cf059/9fzvw5sNjLx42bDS8LBnIn+gjhTVukolE0SMvVg3IJv3vLn14P4xMh9m9YshsApfGuO4v
TmQDATG0/fpFK2K7EyqoKb2kpLkMBlHhACK31vtzAFA8I2+d3jkHWblCaa9RrAxRvhJ/xUEFBMpJ
khaAMMnRuF/PytlWW152jBkq7uJUNe0TRUr3DDC6iNIzhhbPH2jGmWkKREH/ALEU3J9WY+r1kqoF
C4pnFg3WfOQXq2RXz0PweeOlESk6meshKFU92on+nyKcI8+TUeTcFRNei0KLkNDI83z075ED2hce
6GHzyRDNPE+EN9rztErTh+iA0du21knkF9MsotYJYU3BpcfZt8kX3k2T0wljKEqXnbiiQNgBlsiK
lx3pkF77+HjFDaQl3jawH0+say5+JF+L2WHCnw0URRqfgmFxfCRnRShRBhxA027dQtI+C47fGPGo
Y4WMxcGS+rOqy00g12pmqX43UdcyvnbYdLgDF3dM13wbx/HWj3dUh/i038no+0a761aelYGJwzF2
DN/TpWcsMIQqOIlaQ29MXdqcEAm3N1zSmB0itfN/NhW9P+acw8CrRMkpRKR9e2+El3kwTxYT8Ppz
+xsuta/9EB6q1Rh+ZMYPVSYljDdaj3iYhjh9rabykEAgEJC1nrcQkaHOFWaVEyFjkr6z8SPpGr7p
j3T1QRTgCNPMdyXpqntaYJnPfvZQ74VhCSZHSuYErED7gmRfkyov+f1co2KHrdPi0gMOfxGk0M3d
ZB/LW9+SgXzPRexsBC2UVsCj/D3ImUmkuPnTOuIoM4rA+otMWWw5qUd3bwyHahy3KtH56unffIc3
Db+qeLy1dkj9zlzetxXWQjWRVIG/pIjLmjPbQRf7uUXIeFX5dA6bF2RkRN+FPSN4v78J89GfpbFF
P9u+JjBfDjzt9CurVBPuZVbzxu0NghYc0RLTfh+iUkPUNejwbMIosjfQS48tKAcd4yUyTA85nH7H
sALCbbyWlfarP0hz0qPZrWU2U16gScuQkuMOXOP6pK+rRAx521TeAlDve/MJf+ghgqq+wIJ0t+pn
itPAOQOD17qRIez0ObwulbXRcdBeEXp/NZekjwBSArv1Hw73VTEhFrWmw6M5G+8b/LNLxaT22Cfd
d9Jf0zprvgxnTmNOPDqvkbL6be49Kk/uD2VNInqNueMmMM6FMYO+i/kPyNeZkSEJpKA8ZwTvCSuz
+7PQh+CDgWrvQ/XHgJzabn8QoIkMyozkLRqpBBYpKaohYWtwNa9QuuQdjBBai09G2Rv5j5EYmBt/
+jxiQEwJO93nDf6JsFBEpb7VZ7tuMezca0fu0FV7AuD1y50qpyHApEPg7G+ES6bQEQjWLBjRMiNi
/SXyuA9PmjqaElm2issFSne9UYWtNFAQxp+1ZMPspzWttiQnWjuB1V4+38UMgRz3waL4Ji2APNKY
hBMcMlqTxkpcIZThV/rP9JM5UfRVN6mbxyGfBdCr3EpwjuoMX6hjU14bZFhhHVYDO5TAuhd7Uvg2
kJGjrcN/+uPqvwemJYfd/L01OFSPJQBJ3KtFDLI9QZPOS04piQS9aHzN+guuPdre6iaQjOoRStaz
puKYjtIJopEDlo912mOdPuXlMm739K9/qxeHInN4/3HW8ahaw5Ee/QfZenOqlTcdVEuidO3wM9QK
dynd/o4v1gOiIScrVnbekx3Cc/PNdseTeKIF4L7y+r9rNyLGcM/p1ctopyqPX0Toyy6XpI/gIIPd
iK7KCh4ILuPytuWBC7tgv4AT6c5K+RtPM8/uV5kP0Y4yofbEakP0FA/dZ43J7XnH7Q/1jomUJqfB
ug9eGEcdkWfQvqivyeuB5g0w3gJ+tAjvQ7U7v7xsacx3iTN4yyr4HR/UgV/VMCLh1uIXf0siSE3h
KHhNJBLBe9nIFH4L/AG7Erdr8eLrYO4YNWfvH0o3R4vuj94At0P6ijk+obXvjk5FWhcX6S4NrnFg
RZipVAlRp8tI9H3vRIRMv5U2yq7V9/AbTLf6rw3lbiE1N+N56dCe7PJJo2YtzdLnaV/w5lNDeMbU
AF2vEWmuOwFsu95FfBmzhIywcBs9laJW5ubcskRu7JYYrzlE4Gr6hVp6RoE6q7pF8/xs4dbOUPN7
w4aSMJZq0v30viZYsLmafGlyuaeLanCSV2lGQ8kqpbX5XimH89fM90kqSPOO8vmI2p+Axsz50dpu
6HkszbFsv5o5t8gSM0NMgQfa9+zvKCF7wOqBn02/8HPOoEWUE4ZN+ZzL8Qo3PaVn+J97bEPuYJCO
O5Uv1zBo0LHuD4PFeK97P2x4qvtxIosGNTuMyetNF/VUIOkV0Mavujg+VoKMaRbED9ofTDM0Hwke
wJn6FAoIJY/jJ1/MrHpfdwl1ysi9xMs5xl6uLqTkb0J6ebbRUGeMFs8AoqzYnxMj43cAQAGoGhb1
XX50qe4AqP1YKxjoAi1fuOuhlTQndYm9qlsw1xqw6fN3ECJsdz6OYtSXz4p/18HwjM3dzQFMWTAx
iB2nDJnsQnPHfYbPhOnj/ruCQKr9Q66z/5OEGJ0rRr2q8HlZ55frlmj4um0N+r/e5b2bBkhFR5Cs
4npJfsRtK4hmYwrKAEtAmQXnmgXCYoHwzh9344bQpBXq2NyofByIGbkCcjgLoiSyrJYocqYI3epd
jF0QLMxTkQ542XKGGO81vqjMQKVgnySwQFcFT6M8EOE2yd4MOFKuazJwGjXyBdjXLdGz1Dys71fh
PZ94Uvjnr7mkPLmTEeaH2r3vJgDLZOhw+jMMt/YeWxq9bdMgPR1PfxGoDApU15lkiZ0Eq7W1GuRN
5WdeExz+XVNOWcsPBi/07eA9C/uzVNxIxH1siVQZx7YOSYzJ6Eu19dQenKbxqJVyfiwn0h7dDPrw
3nq+S8YYIgAaNLNWXg+g3WuBupetn/FtzCuhQlpw6nxO37b02lKxfeT9ESsbsc566mSFyuzJKvCl
bqXo/ECjPBK0zZn5CzrXlNt0w+uvXsZdfPdEDpoTX0B1a8fECLXN85kV2Rf707lK8s9tuBuoqOft
mTlE0FsAT7eqxFdim3Dy7GaOtY00zTB95LjGLuEwJNJL69QDN7ANYMb9f6A0uorWicaD4CwgcbU+
nhd6Xak6RG4uukc8UeH22U1qz0Dyj7OkxQHZBUgeKBb6Kyn+qOyuphuXioaIato86o/0pA5R70QM
pfDfSaFe0OCHZkp4IDJDqUKEO2phmBdoEVG/8FsfZ7AHWkfBLdOqfumk0RWFzR4H0DqPk7Sq6uOP
mLgiXO6PewW4uclnEK5dQrLJIfx8z098xe7vrtjtkeJb0X0U9zc5MeOKvf88OfXJXtVIjYYvV+2Z
w+cZP5+e+lNS8GUoLEtSpp2gq0W+IjuMlC3exKJJ/E8kFEp8EYXrIJW9xwgpH4GulDfgeLIFS8S3
UdeOAdz+fvfaN/z5iWC/Fuzxo7wQBwuM1RzqI+3e6lZ90j0ALVh5egS6zne8rtBbFXHWXXmLpp9W
kijlFbVjP6GNrvuQ8zEl/gHPWt08yKGu10yTzh6iogBYqeSEFZgSqFbUTO0ZzYZ35wlVesukCD34
HSne7A/7odZdemeVo8TX8CwKVGug5+uVSZQYTj/sNu6jbVdvlxrWE6hho18IbIRAqZoedrS+ac5k
y8lYsetepb2ZK8/G3QH04AyF6r1h1nyoSrEnisTgcpHZna9yLlvAtcToypZVjDTcO2tASpazYv6E
b/WN/+q45ebDkd08aDY1GNxjHVUGJ6sYvpMAFRAYsa9KJSffnwe+3vEpcbR+IcD2Z2knEhbVw41+
gjrMbkhw1ZYzmJY2sUXVzW4Fnfhf8yvjlSVpDEsHDLHRRQ7XY8LBL47VnncysgrfJZN5Sv/EuCy+
3zW7anKRDKiX0tIPnbaUSR297fwIbzeLfzr+Ylk/FrUwkE+gwv6jm39IxLycsp/iMUBw+oy9qcW+
9jAeNMLcs1DrRVSYgWqJmaTSf1e0hBJj5KBQpjgJT6r7IwcYjhe1OFWRw21iJaJgG0h2SDhrMQGr
iyuRuAIXh6DaFTGYEyO2X6VwQ4bnjfCHV3YyN2fFmg7sY4zU5h6Qu/npwS/I5qBPNjSxdyQ3leE0
QEmIfO0k+Svmmx1Qre+lOcIQlhugUZwyl5jNsXOSKjxOWH3nHMvfDZgypKGU/1U8w/ymSWVdIW7K
rUJ6oiZYpGnAJpLEY5U8G2difLMr9x+j5QCHkPiZtDMrDVhAkXZqRTE6GOXVx3AZEncweLMIpgei
m7G97gmKGD0F2bMdXkW6LujIPdFd7Rd/cUF2uAJQIvZuYx0AjsG2GCzXZmSCQ4Ed5RCbwMC4hfIx
w9OhNSbE9AFQSwTWfb8thzSIxrSxzPDS+Vy4yCRo8B0R8y9OXBFp5V9w+RE8mW3cntbMV5yGeT7p
Z66yhU7AzhgJ+8j1hHq1ytW1pDKxtsr9/QiNOcpl2isn2yodN4C5qR+kOzhtGT7OfkHJN4KwZJ6q
l7hoa23q2iYlU+NCvckLnXaQESBJZi8leTSKYi/YU+bhlrqIzfKbUBUeRK2Qo/eNUqyuZ1AGvTJZ
3OehwRPbsnP9pB7h8BJzMJ7lDJzgXcWHQtF/g1K+gzSdhLLDG4dh94jWrl0NY0lysTspEEqzSjeE
p3idDzIkoWw0W4K+U+cG/9A3NPug337NfgamMtCfL9V65R0TPuMOuHoyJYBBqWLQ6oSS+AqEPmx8
aUpkuzkFAyyifwDltx8AFhtRK95kaoKT3twZ4wWo5zbcRBpw4wXLpXGMeQbTTsqoPhnrtPvJWfHE
zNlZUD53cXkBJIK2/fH0WvjrjcfpdS0oZuf6z05jkrnAAG5TY3mmXU+wFfawId8NvJ4Mn5/ro3sI
dk4/8DN+O8w1ics8uj31jqCpiHf5jrILSG2HUHwal+UM0a+psl87AUsQAHliMMrJxZ/rlTcAN8fl
1Xj1S6UXA6TgFvIV1TUidYk7kAT2iHmW0wdjZFrGEQ11KcZ4v/lxhKzS857AaVqFaJXjMd8VZsSk
sB0yMR4OUWEIgx9avT6cz4fmzK17wh50aV5oE5jnyrapozslLT6VUDRn3Uu8JguLnY2l/E26N2dF
4HSxxn01ruy8BRYUJiMJVmK0idXDlXYizGzzB68+ealO+UiGQJCS+CPy9x2afnx9dLF2g/UFJi5b
YAXXrYwZx2nSnoJfLO8ahsNpDTIboUz2a07SxS/W7/mapYuxTotVXXSPQsGRo58Pil/R40DjvX7v
Qe0KoNhW25/xMDmc17V7f6WEGmA0vBi6x/TNOgZxEN6bRvm7XdhiCpgDIhOSaaDl202oAbxjtdbn
GWygDT+KinqqrpEtd+dwrvb11OtRmgtnVftCgPwVjhG32vvy+LGQJWWHHVBQi+CCsWI+YSDPkvEB
AB5hQ38FPzRYuKOteM2BU+Ueu0kB7Pd6SYg2dF+tbLM3iKMSDe4B6pOV34Ll/jRFmGnxpAVIZhfH
nCuTxeNEWLBrh24wBEtFBw70GyDxON5AuNmZlUAxJ5D8wKezH2SfZ7iXdnC6De02P14vrNXCcfHe
U5OQ2CBAaKTcGBuq9fMjnncwIrf/2OlASySpxojWO2HQydKdP8P64TBkr2qcn31Hy8/nz174Ey3E
ixjOL0ZdboHWvm2zCeApscjBKut4qeYa1Go7Ad9UaRWPCtlF83EMT4/7hFDklatuWY2q1mJ3MdCk
1yJY28JN4ywF0awvVrJ5sVDfBwbZHcVG9Y6YA4JWV0jaBzFOeqZF/PpTGv5nWYtOl8hXPdMUHTQP
mHxrM7n/hMdSt9P9PEfJ+Y5YmwqyXcTowfdkEcJjV1domp67Jn651Q1AdSnn8+iF+9XBiW0MVYTy
Mul4X0HBZBwL0oM6L6kNl1e54NbEmaM1+E+K6TpVCa9PPANICExwgrVGhH9a93lgRN2ITK+lzGkd
xSisolsjhPcyAxgLUcncSpMsES/2oOoCCapwk6+8Yuv8WVy3iGWvxPz3TyYMGtNFZxxrmOlv0J5T
6GtBVhhqnfrPgnkorrWZmZ0l4YFkpXwawofi4pIgvxXShP9liihIoyJ8Pqacf/btmWd62axbjkVK
dh3EQ4L/d0TjBAnniJlB4zr8O+Lx3igo/tQAoCWURdTDMVY39YhhjB510UDRobjnZRcm1D1+03rb
gKzkLRkj8vQvRCL7ZQqHN2LZ8dIdJRdpkwTxvmRxOE7tmTvCiwU25BeU6nkq9BSQAC5I+j2hNzDY
2apVPJdtHeOQILU1zKWcqOBvpYkLpOU7QvUDqrw+2ofHU48o8BkgyBRElmOMKVc20WTmCmaTeaxr
AE9kH4BtmYv5C/1wZ7eUmPjxRJ9cdJczr6kAeVt92vM1bIJPdVXGCcuo6JFBg77hoAAA5kkCEAD1
9rXVDTfiPx+Ger8O+JJyAi05elyhhPEUFWNgYJMPn8eMu0lch5LBlP7NaNTB+9amNpEyw45yta/n
wbeO88ZGPPey6k3fqtn6uYILAPJTTPy81LRyHuvIbsNnXTFrpHRrxaLa3SpxpiQpz73ts/0fIWBJ
h6qFdwffPUBap4xc5vNQ6eYGNhj19wSlVClvdJR+YAU3SrYG5slkGHXIqt1EJMWQa1im93ASo/7M
maEozrPHNBdTJOx/TzhWahtaBh7gh1kE74xnl/decIfGYOcxTTdENsP2H3sZ6Gd15SKEUKV4Wtiu
6ENLIUIV+3mCD2J71mn+3doyXSd0L3JL+bUe+SVuy7Dr22UrPNoSRudO0FBDh2CFElWrPyG0ieqa
/S9A0Pvr/+3mgqxo3+JDuc71++Rv5/mUSaygOlVuoLSsB8UKEouUKr5/bscK3fkV3uX+9A6bTp2v
d9vlT3OTHKmwEBayIZv/cODwOV4InCzY+v8mm2twl8D2KSb3A1hwi9dHVvQ1fqxec87uKm72VAz2
4UE8FKQgMv2IKwObuze6fJCile89AYGyM+XUDvLJPMIuM12bzPUr4T9sM70W+AqjG8LEqzPxvyYc
qcHZun1aqWtur4SdRtDIwtmZsJApQ7eytGMZ/DkfZyQgAgK+HAG/rC/UremuTm4rEGY+cQg0boBD
KQEHlcgyDDU1J021WdGvzRfdc2xRaAx/ibkqwMFpEbdtoteamzDieU+krIB+gX5uwISQki3dpN/q
wFYVGM8BoVpBzO4B3Pjcjp7bJ5gESC4Ra+v2DdPBNLis5HFpOOYqRCv+5zD1wL1j/N8KYbRf60ym
fGaNiDNwkuTjHfxTSwZ7mXnYsovJGmxpVUmjHKnIMcc7OWx8oQv76WcYStY9hFuZ+fO3INlLmVhm
KF3fNN8zMrUkEFMIw6KbxsqhvH5yrlFiWCtQrsQVHqwCahHbKWjZOkJ5uJoDN/8ILJalmCZ/7qjU
c8tIaBBXXxR4HBuz7dm2fSw6h/ieBtTjKHig/wDEz+PXV0J/p6Nk8oI6h/JDiqbmB5RNshWyyvHO
3Bc2CZkrpvKcT0FpDBhzoAelZcduqO5SBPZxzM6sFTqHVLjPSVzcp8k+GeQIA7Mcot2+zQA1PG4o
R/OV4dyFd8+DlOhajtxwopM4Fd6hKs6g/Ndm6z1AwG4K08TtebXOiHAMbSHZ750Ix+/ThGMQ7nCi
U04dhX/1Z6FYbFgeO3c6ny7QPgQlVIuXxiuFxK5dMgLc8hy7dr39zW5BBvU1GLEWzY3fPJw3P5JZ
e+MATFH6jHNC43THTqs9w/sHmq+Ph7F81sWebLrmg4x9Jqq+6Awbn+dif/XcOApQHzxfibkbiB/E
+RufmicpkD4rgosaWPsEkEki8ORTzQqxa38GvcmMPWszI+2CtsVWSwq0WdQC/ay0vxqd/7qlVHkR
3lctP46vPmZKIEtKOZSCzPc/Pw9Ocb5w6olFJiXamxsPLh2zEsEzyZ4cwPEIHYCO1Aw7akWkZEIu
o9LzpvrJsQyYQl9EI6t7iB6jgVKz1+B+6z2aXUE4OIuyX7Yv+H0vRBviGA8nZ/7ot8eX40qHZ6BX
wyo22C6ZnghTD2H1JHAQKUesEBxRIKrxr9/o1sHAxXONT2Z9Zpg0Q/OsLM/mWKhSQ8UPyT/Lw0KP
mMj9ulnEu82Auso9Q7QHSvnsI1J/ICFGPq1IkcY3m3V6UXUM1+Mi03/Zn4NbgsOZffUXZNhYQixQ
eoSPceFIJbc+V7Oj5ZZs1zzHlaryyfsoBgbTKcxRkHwL7X+jH8aNpWXwpuNH3/vPfuvW1WmSzgqz
1G2F8TTYdB/+IGNQ/TP5CySVr6pioBPlmCcJfEQRLHW3piuy15Tqda/vyC1kSvmWunY9WawRAfWH
WKI40iENOsXjknfuxJxpVkIfTy3Sn5lNNaujyDKE2imGKiFVA8ZZPcbeyk8RyByrAnYbeeoHzm2I
XFixTn8KFVCG87BkPNiMXjVk1Y5Okob5VZxiFVxh8Y319DBvISa/1SG9OOX+b/gmLzhUkpO5il2z
CnGpvrnmL+CFJSQ4WwyX1THlo09KbHK7kQg8bds0QOrpr/7KoEnI0uBHKJRBqVd4kSLTjSoMIRk+
IZlyBhlxfX1Hjteb1a+JaCQ4csO684gFdi9V1yv58nUj1Jp3nJIPMXiCOpcMHsywqz5bMltg9DQ+
W4x89MJa0djzzb18htBy6Iw/xK5jNb82pdgUyGyvL1gaV2kHoXHLECZN5lIEllWpJd6fVndlR0+S
RUmc3AXCgr1KX6t9LeAeM0q29YdiL6qFFIF2ikUMZPIBm0tGLX84It7hJ68xjIcRmfgEAP+kah+t
yXE3KBRJ6qkIr0G2B0hOhWxEiviow3a+fL6j73UYYGlCzJ3c043utu7XGnMP0jm0gvya5ntv4CGi
Dm92M7bI09V6HMh1FKmuvmxndKXK6cxVrpZpsez3jkV6j884gpGHzrNIrB2dZgBjQFGCr0UTL/DV
l5kpXHobspP7STPFEm5hrqRGBEdk3/JLzyyf0W+JtkkVDR8712a2NCB6iaH991NRfyu9ZO0nmo0n
S6i99eQzdUZyhK+Qmikg2+Id6weYs5zvxMkYigGxHoLzTW5vf+n8dTnyDTvK0Eq1ffmbirqFkD8y
yt3ls0/bIAoOE6DJ1FfLhLJaXqtJFNrG79ykFPQ4h7p4t5AZrSyApO+4xgZa+1V8O5dpTaeAnLA4
n4wFfQ5OhoXnbo4y/qaefLqmHw/KQYoUPEg4NMs1FpCmZGeYNV+hUgaluPrOWOZU+hm1u1f3wWZb
lKsbD3unVY59K4BB4DhoDW+AuM4BfC3gJW/VpJDE2QAbKXeHqxd7bQy5uKu1clcbGmXjvkobWfwt
WtDw0W0sxnK4JDOwQ8GQq28A8sTa2Uz0rmXiMcOhNNPb9e2Olgmg5J7hVYpxfrrpCcFQV5JtTT+D
Fp9+9Ak0xd12XBtyitg0q9ZT65PcN5krCJ2F7TelTdaJ4TQ6z7kI0CMzzBS3dRNZGZpdVmSVKsyX
VNn/rhOv45GJ4Y8xRfe5r0eyoYT57hpWCHbirPRtWXm2q5qV/+nPJSQVQdmPZpZxS/BUBzy2pCK/
icDnLUpxQ62GbwPGL7u2xGoD1FZOe5acI6avVOy+K6+NcgxMWG/yAfhRE9PSXo8DK7RTDP562s3P
54oKgOYD4T3z6+ZlbtYBTZmv8OkwDx0C9M33tlyMo54OfcpR8h4Sahs+LWLL66zh93a3XYwFVUhU
FOGWfESpIQOnBfenoAKBYkBzg/Qt/71aEtywGvrcCyTlGWQO5X4Wmc6bWTOGeX8CglZkNNHCBY+R
5PbbZGdfNfgmE4R0PnJ14FDDfxmKhtiink5s4FwM2s/LKCLH3qiKTtOkvyDjg5BDOoXMeohybT6W
KG6f/Jyt5CixOgIdP0xlARRv7uS+Wbkd7j28qsgdNFbQNc8iYAS/z6DiwhGNx7WyckFbGOSawvTd
uaUU60gyvydhupkMEEMj+AOXOiAEVfDYVN8haBqQoH0RKWbJqHhu+wHdacrqHiI2difYlFTxgBeK
+YX9XAw83GNDGiGezUdVZwFds2YUNGdCChYBF7zkNghNHsGhg7FjbbYFYh0MQ6pbd7/egLCuCIO3
56Bwp2Y6palFK7VqdtlC1ERTqlEn8EeCzDBTrZCxvmQFjaktyYTpTYOOx3Lil70/RtKpCeZGpuXj
YsrSzeY2IeWg04oaiWyIWrHnE589Nrud1Y5wQwi4onOG5ZEGKKWJepwbx2dDRas8+XcsakJ9A7jQ
AdpXK8EyM6h6CP5WqxYWXTSZMwdpGo0Tv5madX2ujZG8JVpUSDtuIdoncXG1vubntioeQWr9pZ2s
9BFMT3CjlRs1ifaIZYykLe++d/tUPkhmhHtUdjxb05NVicH2AecVfWeHWCJUTx3M0rPicX3lZuHh
a9OHM/5L5aTqh7+LOTwGvL9D+f6WtWdI0B0kU4VTBYu1CjHYKzBlepKIhyWCJffGGDoRUM3oKn4y
m+m3r1jRLSQVwZXobtK75zUl/0oLFbmxTqAO2na8dvmqzexkGqYQL97hBQd4IktlNF7nlkJCZeAs
fHfJkc5f0sPyq06pILvsQ2etnfnFhKkPwIZGJFnbBpcSIBpeD9Wse4SqxRADI+cps9Zt7oLUWLYL
jWAp2R6i0lnrL2QJaoo0U7l5/vToUCG7x6AYIuya+UtcPvjvWlFLsEhxDvfTpU++PgZzy+eSmBb+
wiPObAARXunOk5gBXg0edCSFjEYwf2FQhcXbca9lKWWswrkSKEO2tHC4dmRwFIck0/g/6oixeoiy
3PDUHbZ4ZRmWr7SEOJuX3VqQ1WB+HGAogGhmFe7tpgAkApTsUV/fdXJR70wr09yHVq9rlr9cyCky
LWy5n7Dmd1ZKuOTOik/LybhN2J4XkASOKTMzmXoNW9zaUe5TPSGZiwRASD4PSHcY2revdrVhrH8A
jXFiABGvuaEhI4h66B2TP7WxMmoabKNGNV5yIMhrj24rt45Lh7xH1MGZ+Ekq4a7UNzNdOHss69ag
U4n1I9XifJvJxFDflK957vf5enBuqZOcz8AqUhLmW2g6CLhkrTLKUo4j64LKPDj7wmY3U0lxWCXT
2rlszkJ8pxdjDblDkUC2pX5iEPPCDB9CsL1lg0rkuWhgGkCn48K6D+iTH3alRCu71eQgcn0jwQ0R
7LEleftdIFVvH4hZnpIkgpcZJA3/Tz/qUdljiKsmdcZ93c2nzopGffhzWq254IWa8HYF2/GdMTJJ
+t0RhO/l0LjuWOAFkrIU3BDTocuWTvA/ukmyNO++fg+hj680i12UrGb816Yft4T3FXEHQf0SKY1u
BBDBFpKvNNwHH+bQn5dUvkxOR/R+syrnk9M9gDi1MJpeEUpc6DLC89ZnGI/uVfMW1q4hnHq/7/cc
+b1eRC4PHCiHtBWIzTG+Y+82t9VgFT9+SENJ1hHCzWUVUeC2ALhhMd1I6P6VeTYMYmrqrEXFCchG
TTNXOvI6lcUluyZAJ0/29MOOEzggHLKIujDH7aaXQF5gjXGo0KW1jbIBU4/+e4Sgnnsj1X2HJ1CT
VlzCvyyNwTWsSuYrJQWk313rMJTYJux+7YVQgzkhE/MwpZu8x2Igtmi3CrgrL3+PaQFlU+H994eK
tLCaTSYfduEYo5hpfHZHqGwfNN+urgwOL992byb7GBVL7+DrBF28r135IJJVu3DFwpBUDSr6oG90
VLKPAWq3TqEOUzmNLcxmkkMp93YClfEDEesTT6nmcNwG5XXeEA86wvueXsQWRUgwimRPTBMUiHFI
Yw3pfMWox52vtaiMOO+ty/USB3TXoCJTnA0WMGfsifdp4sHi07h0cpsX3f05xKF83z2KHzMpD1QB
2k6ivAp9fUyi/JrK+ahIqnGLo5ilWWOzHIARwpbSZDPhlZYecUHpvPOfMHrVgCqYQyIkfVHgSZYA
CnO5AJongrOy0NOoj8JG/w8e3keUrXMbgQHnpp8TXHJCXbHxrFm1OEj/QPv9hn05eiNoENTquvFQ
aOZ6crogyZlkcMMQYerBEsIB8CBPgGs76fG1hI1zHo6cbrZyohd3TBnpss6lXuRYCuCpInTECBjr
XZjV0PlG1XJq69o0DUtR3u6tRELal9sie+tCwTwxobvn6rQpIG7ByLt9wQnXPJ9M6AQjbT72Sv0h
Kvg0AZ+NITj2EbgH+5i7yD06FTJtLefXAp2LOIro8gwnJWuSkG1CiP+WMKFAw1dF+FzLqTBdSVRW
fdfLxv5ySNnChXmrvzgnn/OEMbQph8y9gf9nxkyEMh1qAJVbm994FkmEf5hI2+eQF2eF4u+4IeAc
APZ/0jhJSBXGEr+Vwh1hhGFUy6Z0aSfDETOn362R63zANGAIt76tVy0TzvukBU3mWygHqGDDfERD
ALaO4ABgaDFQJL89O9zYJuaStmA369y1x0mARrxA4i5gWKwPZFrr2/L2eGX/1BWyO0hCpggz/ebe
vdSSY1oF0aa4tb6aDaEN7YUA3C0jr2pe1dvNd/d38nkr2+3FkPRq4Vvs5bQbkwdmiy+tTVNoVBMT
nvM1Xg1hB3LrZx1h/I50KlgFAEk1HfeuLKyojq2yOVxoCjZNx5q+R0GPvswfwtEnZYIjpw5v5xzq
huh2y6Ik+6jhwOOJXOqY82q+izpeMp7vdmv4RB62NvtOK5dTMgu8WCbSEhy8bAkkXeaDlhdHlhwN
zgAOJIn7Dj1mQgL+AGnevvNiv8u2BR/qSeGwMW4XfcMcV9inD+w23YTqts8+a/NI2Cd/sL9TE58B
zau81FdAdAG+4h3ctS2IeNQdJp+lEvqysRlSpgBdPP3SeWS/UNceyeym2l8h9+p8b20mn9B3OC72
uf2fcXehDRgac8bNTiKOyNfE2Niez0bpoRJVbQLd38968IvJj5WzUwFx481F5Kb4UkKyv7c18kR2
Z2JMgomnWUqJ45qquWL7mGWq2mj4PRlUQ9W6R9ejd4CPpRwQUGukynwF4RtiwyDhaXb6BwWqfqVR
RgD9WszrD2kU4XUU/pre2/nu7wkSEZc7knJ81tUtk4QZFoe3rRa2iryNXfF+oIdWrk5zuqRj62cD
hl85xWnB0E33nxsFowzIo8yuh6z37pCtD+x5ox0tFJf0eWX53dTQcWmBluir6SZ0NZzib/91/6n5
uJRA7AQkJIINHZI0F05CwlNVZlbEa6OAcDoFuvvM8HHX9XrZxOB+abMRJpR1+8eaXT4Yo0zGWbCv
CVLKH9sG0Tni/nG3UntnwJfzUFoWTr78L8/kugB1jo5x9N5bUximCzP5N3m8i6qNtRzx8rREvh/j
cseLzJDx8NE01FRFQ6nTBPDsYulJUOlhEOasYiFjA7GmU2HQlYg/lC6V110izYewxRZYGgyRgUKJ
Hp3IJ68qJUCLj1UwiSZvShO1GYlleyPf38CvFJ8YicQX7xmcrb9rDM3l5MUOYPKtL0Txd2EkiQky
NHRtLhh65tdRRM1xmDoOxoPKq0CeQoMQ3+y0h/9CVjW2glbOxi8ktKsDxHHmDWUPLXwhEKYdH1mT
3uDHGHfQChpkjcMYMTvqsjzgcED8/fS6TXyn0D+I4pXoDPOfqxsbUObFcO2SMdQET0s8EkKIsWgG
pHBnZqK8fGzEozEU6ut3sJAW1S/kqQebRQQgL3DQXwZjSt31HYvXNnYCkWrpQJe+FDW/iRm0BSTX
0pENBP6DAfCPN0+QQq97JvuYjPpYLYKDU9P3ZX/2wc0s7Zq616VP5PO6xiUUw3H/16lIcPOn/lVA
BwbdcOFv9ZR05VIG2yZtnRbv8HxC4xerpblgz59uAuQ1MwnOSc7rG9/ob3OWdestTZ/jBl/cuSuq
rGXqvIijL9YTqkPWvJ1s7MHbBMWK1f4s673aIqY93JKGkqlgZVoQB4SFNCS2aZPV5JNJspMUzTZ+
HR4cGX0HmV4syR6TN+JjTrqpvcZiPB3vSTMc2wrO+sqzLIznNwu1M0FVpfn0a+sstsPrlCcgMk4N
6oIzJpbplveQ35ai4TgvlPjQOAzWbz/nWr3ulojYaieB/oLRhpKXPaUoarWsdGftKa8jw/W36pn4
RIzw/rwxsOcq1ofqlogCsHSBcAk2BJalTRtNEJCFJRcDJpJlN2GuU8Rc7JSMjEnL2tORDJCUWDk0
PV2JlNIcDFez1Aotbnw1D1EzMCQLWfFMiiFjV6mMsM2+nnFBtI7lC1jV059/YGhcNfhBtHowUuGE
N+oJrpNWh3t+ItCCpSA0Kxt6uvFvlo+qwmrcXVWMnv/YG/tnIKlZJYax7lVlYWZUkstXv+E+TehP
g5+uRWvZMk1jqEjhBM7psN1lvIvHAKv4eS2iXVS3+mossviCw+wowCejqCaMgYuq8QLn5DmLsQoP
bYcchsYPEgAmNlI8IPixOcexp4hI6DEWv/IzC7LV4u3WWjg6ZYpjXpyu6DuTNM1UqbiETl6Eixkd
1Jp/yDr6DUm+XTkKnsAmYIVNA1OgumwTh2XAtEJexwEJcazPgaXC0MvbtT/2Q5TyH2ogNKms83Ps
v+daSx8gLG25ogzcIRu4/8UaUUGNa1aIlZLj7+c0cLyVyzEyS5dmPuWkfxx0OGIvnZUpZ9+26ehY
g8xDCHM9UJ1vnHfAHSM7kgRuosoGVYCa55z4E9qcs+0PlRkTTaXqeUFTlLM5in2xGefsVmshgLXS
9ZUKECAEyM0vZu/ILrOYuq5OGdvODxqdbpnZbycVpYn85G6hiqKCC3h8ktCKVDJoxFd8hTeN8uHz
R4EitCkjOYTVa11ql3UsnpsqNcdhMh4fS59Zp+ywHdb3kGM+9jHvHXVYaw1XXWhbYKig295vbgnw
UGd0liv2Lmsam6kRCXafX4G4YevyVsXw0dJd2JZ5+s6bwPZnZzqMWYGPnL4Z6j8KVs4vEGS7Viw0
z4xe6whskwwyckZFezHhmhtw2jAmGMEh0cE+TDxxWKjHR363baHr40ciHLk/9qQwcPIe7/jsrVmp
X/siyEK+/pjAhMM/Zfl9VmUAfYpG4RkBLWUrji2tSyLKc9dfnyiUCDPd3HX4jc0nhr4B1Wg/HQV6
fn8ccstSG5d9BIiTEW50YN3oaCOV3uQ6rY4OABXlyO+tPWsPbeKw085OYDoCX7VGxR+vn4NVOkqn
fNfadWn1aMzfWdwaiWtXVoZqGOQ0UTpEqSjIMcc632DsPp12Vzns9YHkO90b+hXMgfIiQ1WXX7Ni
uGxmwGi5I9m79bps1AVUIscaE19lCtyWTG9aB55VoWT+zkExK+aFbMH43UxNkj0vgTCavuBhvaZ+
oGKBY2bruSfIfQ7865emSKtAoe245xWPMtAnAyMBJmCTMeUQC1UkPqQ6u9GdYexWAiEBb2GqToaD
SRP58dIabt0vCAOjbuou6aSdm2SqlUDxWNKGZ005dkiPELYGfVoEQ0xj5zwA56PHzL4eadN4TZ8r
LsP3iT1T8yblcRel5kOFIteipnDdaXn+qIWHBja52HiCV8xN0dNnmGeWwAQPgMDFZpM3f9G6piem
dMn+YfiP875hkLKTxCWF1DkgQoVMVzCloAVNtGPMdgVefMVJXuoP9yZDQorUogggwLQouClBR3lp
p7gG3Vby+/WKI7YbeJVToSCSC8TqctivtwEpfrH1Y99bdhmGDkYa/9jqlJ+rwo0wWEvkNjO0MJpe
sqpM7ghhn32yaQOYBxoh+JQPnDIp+ZRr4VKYaBJoh9yzS51HYmvnnS1+NPGbB3FuXLLSyvA+5WcG
6zhdm3Q82OPJInTqUREdFX0lUGneQsBY3fG9sGQ+41JTrRpvjNBimce4EEAhyPVrwdjvivvJptg+
HXSGbMtKh109se07t3igt7USS6nK43N4h/SIjPrwIvS/PKfPPJsq0aLgcoUXA0v6Y30EnvwbQhIR
ofzcUWgk7FeGsvWA2UDChu7BUySWZGUAFiD2Emh/RVmjCzidduhGUFv5xjmo1CNSgzfr18U5pSiB
mh81l22yDtpEQoYknjf1M9TvCEh/8ize5fKN4Vn6C3UMWk36v6toALB0SyQshFray/ydWDt98LCL
FtdJEMROJklliHeTP7lYKPTtKVHuiKWs4JmiG8smCqVEuAgToMqfhDJBW+zT5mfd4JOreUEZzhZa
gx1fRfG+OHPcfOEOKjHbry22p7DlB/Lh2YIRUPTwLS5w5ysp6W5zG6gAZqSrm2Hdd+wSbGrQ87Zc
NASspJg3LoE8jASzvLvRTO1yB4LvNIYiCWVa8qkAagxdgkpYy6bj/7JEKo/nGt59+1ft8TfjqZMb
B8VFLxuS2mBWiqERBNejryil2elvTNf6LFjVkWXze2V7Lip6gfw8uUJH+8laXGv0Pttao7eXJUvE
YmhTgCqkrue6viEtzmt1kbMat+8/wL9X5oom/8DpcjqnNPDRlAPlQSfn3oqHKdVK5LWZ0IUnjBo5
K2i6H0lCaFSMnXl/FzQo4onPKwvJiGGyv7QOYCNZfVTHZvo9wppq0O/gUhlYmwObM4dKEOMTB1GW
H2t4/W5LhtNcYc/wqHcYWz1ccZJ8z4Y4GZnA/JH4niewbegna3Ma9zQfLnWPduBn5lfV8utCK3JG
zajMP28E9Vb7/8RYrTg+Q0uk/Mb49BOrAkFHUAYLlRJSlvs1Ppphfours+xCePLboaVQc/PPbAHn
cl96vG8h8H/GspXT7OhtCn9K2SdU9s3lSvgGuvIAZGh59hJkVDLLMZJxuIVUxeSorfL97S7aZqDX
hgP+P+3ADqU/KExu6lZCYvnLEm+lxXEgmlire45Ewdq4wyOXIHvn8E1qRQtn+jWyz8Dm8OGaLrCM
FUhLUReKZf+4JiQXe+gXx7mzHUw+YmrF4sSOsUho88o+oAokWQ+cxDwfiy0/P26syTMkE/Fw7/WC
YbT8/MHowxzpgz3BEC0aCtUmLE3z876bYahJ9BCGhrkxnk1lp2LLyE5BGlJ3Pi5Fx9/FI+MHdLwk
X3JCY/bairCIZGJv15ZfhzxmUumOEIZEYPicK6xaorZHv2f+D0W5+iCPXr9GZ5BrAxlQSdHa2r2n
nWV+rLY8J6tn56GstukF42y24W+YM+Rbd2In9MX9Mgck4u6no4QkE90u9e4yncF890N4qz7JYb5C
K41BYO8YOZxlmxFGRGyQV04LmbgEcrpyY1N5QRIGwpa7H2tV7/iNM2Z8YqDhZ5JM57mA649TEBGR
8Yo0+Q/HQeEDx/LcPfSyfzITwlyILyb9iMTWe86cwYUVFCyhC4sSwCU++CwhPvktlZHgllTEIOrg
9BJ4YCqMSgfvNqTsy/fYAVitwWqcyZB5S6yWUWTAaUaIhHeI2KYi+nLdW5OPrS5nOt8aobvZV19f
umCK8HahZiqm1TNwOxiyUjpVfJwDSWX3sq18X7CmBCBcmz3JSfXlX3eLAkwfrvpwD0FyRIVjt+p+
ujHqqCeQ1Jkz2lZFTQpbBol+HlucGgrpVZT7m80uRgZ4EBRfnkhO41mE5Jg2ypYX+SCU0o7LV8ZX
v0Pn20Zi9rJZ+Wm+5mYT/pfs9SLFghdhEMrrAt8+311lnKvP2Hi8XjtPoFn2YFEN3xL49BkDfrr3
KvBg8EBdUpVsIHrveBCURTZNyEfGuu2I49nQAxhGZO4lWxeFLQeOX9IfXuSeJC7KzSAob3mdJcrN
Xo1gY0PapygKW9TazQumvry9TI5zUUJbgPUK/FLJBdSWlKp8WeD8ullfoXH+XR8aop5HqkNqLh+W
NgfeiMWMOW60DZAXNZdPMqZUB6/2g/O7e1K2jIIANN1cQ6WWCzZWiU7oTSJDtDBlWE2bIW7u1b8j
Yx/k3phumWGV6EsYu0pqfIaCy3ivC/GS58CSKdjAmQYS7D/8U2NvxgEPO+RULMKAYc6UQESFycxF
/CuHXooZoMm7y0qEG/oKlzVQiXr2PEJSmxs4GVyy+L8R+jn1dMF13Aw2b3MiDBvkusWkBlFpYhwk
fwlIaYGU2MeOC4erZxE7NO9fU4rpBVUGS1W9jfmcObM2sDQQA27d7LUA/sbSj/bKToKn1xhFUeuN
n/Oh0XYQ4o1rfNKLLiemj5SDnAYupGGjI85ZrnAGa3/XaLg/OFMHrkG1Cg98nSSE0P7ZWS5U83yG
pqSdYlY9xilt5UpKjJKMOm9x+sCdzaAVCJrcoagJi41+gCtMct0bASaSz98+sjR75NvUvuDt6yCQ
/sgTIlKUKylvjJycTh3+yxG+irU77y9rZkcilefsTr6OmY6RIg74CG0r6dtdJC0blRXqLMm3RB5B
9EUEPLHCmrn+I8C+zgqIlRtuwgWqlrUpm14yy5VCLJ6SrsM0m6TECU0kcm1hkKSCYkq//K3CDLHc
e95VO0bzXF+1FjJtt6zX6HVfqGuimaGQcuVimrtHYRUyzml+PLNTWKLbKDVg5iKxOPxw/B4rwSMB
U96/dN9Kz46R6RFGPih3Aa2H5RW1+eNKIn6Glh34W3Ne3rjFmdbXHj3bPxD+8dQAcjKwweFiilIp
IbgNFUqtB7embiwkgjIltw28QYqFwn9s7+iJWoZ5fJf3f/MigRRZMdZmDR3laCbSzV4bItTy7K1M
AwhY7AKb6Fa3gdy74S3dCPSPKvomk9IvWDMTz0q931wr2gLh6EGrgNzFzhizAsVVqjqH7wAUQXcm
zM4GzUOBB2Z823mavTwbMRmIMaXq5pL7mWAQpmSPhP0Vav33g+O8Mapi24nFIuLYLu2Zr8Mgq794
cDanB+XxHbYq/V5vIN6bq6fP6e+Ae67EnYrmLVjqWsTZ90GRm5FsinTAYmCSLMwOFXfRx8gtkdrh
hlu2Lq1A8J9Ehq8G39PeElqMHwDkXbmIp9ktYyXhvl7ocaxnAl5EsoootXigs5kGKCvWVnRWi0s3
HJmU51uwc8/89YbT7uiYnrSl/G09EST5+wIybBPZ3KFL0JVPp6QLAaMI9GdRMemLWnmMzHuKyszR
ttfLLWF+WNI05r9kMasZ1kWQS3a/SDDY+76GQFeAj4+QgfOBZp2QXM4TpCY0PxzwicdYecEMQ6cZ
FubCeCDkmUEOVRLD00XIwsoA5BlL1vIsggb/qeL8VOo9f/4MyCI6pdn1laLGYdGTTfrrmXjneTGt
WydT1rB7bG6XIvO2xBK5K1ow9aza7z28Vuy7r4pMeu+jVpcmJGomwIt/1ghYIhJpanEYKI7VwlOX
phN9iM8jA6Or8FJJUPYrWfApD6O1WZw26pqtHj4HX5fBJyy6MlUihBbqroddw5monP3v/aGJ33ne
XUFHvNx04UPV/9oYrQMGDijQUCDbDgS0HjNNZZty5zlBCxDXg6avGzTFyIs72uA9QzxphbqNxKWf
7fKPbMLJA67NqroXO21HusV+ZTs+RP8blVEIt93quqblmHoUo3MzMRdPRgisxDERamMwvY3cZE86
Y2xLAjV2dS/cpCWoZcnK+bcgatFidFXPyI5jTb7pap8HAzCgeOemGbHSMLFjuVVsqUQ+UlVt/RgC
bQ0ssBKUyH6SXJ6YU9IPo1Rxk9YS4Pj4/sn8Y7cS71vkOQY2H7i5/fR1ByZuvVQUZVZGIkFxSSU1
hF0BW7ngALwQy30shjrJap9O9b5b18PthMEsDCs3QbtUyHFqqhDDQJRKMgOj1h/meJYKVf8pPvsd
m1nDbOW6SZXt07kpzzOHWY6puoOWg+tW1KTbdRhAhWzD/5zM90aAIq7ntZIRusNBy7emm7eNlKrw
GNtUcYujTCyiWsXGu7V7pvowU/KCO5uFTQ3ObOglzM6uySEkGYgoMKcpDcfElcz8Kejp/vR7V8jv
nbVVi4eBhSLEEym4YgHDbiCXCjJEgMzNRrvJhu/SBjPsgG5bdeRDy2WvY4ClcFLzbWwsn/UJOjm4
f8HqRhoCbofDH6sDWjtd4Q2GI77G3pMAOs3kRfSCoXed2knLaXabgyROSbtfmjasECjEpLOC5sxN
HyKEQ26HJELIVku4I65smwJzj4RtkcLMwEvgAzlSPBYbw/oS59LKqlvG/aqjPr4BrlBTJL87eJGt
GHXXDvOy/WWCB0ha++3FmG8eyQWDLU+BHnZJVhoe7HageC22mYstAkrFwjrOI9A/8I34rxVyAOF7
f/mnlVDKR8qxxLaXU+gClCSs3gn0JJ9XIYouHTlte7KsxG9amPvIXEIbGa+sSv5Ta44enqn0VtAy
8QNzdvYgW+TPhPrMmUI5zXhvkX0kZszaaD8GmvXoG8q+38jZs/s8E9uwS0kwqRGbv62zs6VBbox5
I0uD7f7oasBG0QEQNtxjXkg4XCsZIeuVB8uippRXf220zA7K822qp5N1ZudaPZJfQPMRlkg/diPo
XFcOl8q0kS35vlveMmQgmPk6+s8/VUAMJi37Ou9erGAzKCGPqSLcIsuMHslAIs+jhAqFpsvcxPRx
F8omlC5yda7SX0KFGGVTZ91BlauHNn+OxXyDkRUdmIqXaGtGtR53cTMRPICm3l6lNsmjzyKZyVTh
pr9/CabmJrRyinq2LREXLs5qVMq4fT5ATfXjdQVQETkONaHsqYpdH1WtXKL22+88wCFHzwJuAoEQ
GA+0AA5fhx1H1dPG1kB8TS2Q7TfDOZz8nZZzyixsOxE4xuidbARHuf74cpnt9zQYt/+MaNs6cKPn
zRYnnWT03NQYP2iox333sTxQmwXSRn2CXaNhgkVTYVkvJ4LDq3+woN7RQX8ll6Gx7sF9i/21yK8w
Vkzdxv428gv39TKy2e2sR56GzUJ4C/5N55BDDu7IvWXqHSdWAsaBFCSCYJoX3f1M5bSTrJ5VejYu
DJpIZm2J25vOADMkInno9ulb7v1cSWt7zeM2wMndu2eIXxw1udfQN5lgGw89AH3xzYr0QbJwOeEf
PDVAmHD4DlUeV5Bo2LK7Khto/wYtfzTibxZIXLqMgwDgL39LafhzBoonNlF5S/H1GJmlnMTCW4IO
SsedfzP6wEXxP1dKYjJM3H3XGASbQCZpwUC2/XTPUdceO7ec06gW/uHDu0qNB5hq52VvZzquY67x
m/fogbaNIavPOYb63fXsPz6Hpk8m6qbyQWY21PZadOeWHDjO8FUFldVonpGM0TuuI++J6HNBF9l1
507Rhn2sDizeC6EhEV4tQr08/iyiQ2wpkzJ+OvNE6puMiscH1W+BeS8LNWPhHGmUK7jQEPEdv/FQ
vZeCpxlZsxOm0yhs9xJoLxw4GbV+kFIvpwK/zEVawhgOhJA046Gg1O6WP+AaTQ2Fmcazuiaf2Zj0
EOJCco+8bAzf9uN8UZquClx0fZvxsRrLt6zRAsa5OJ8NtfekpBgYWutfgJ40bneaKMrPXRMyROR3
Zwg74cIjNFX30s7XrwopiV4hGG/alZ2TPcucY7aTH2u6Gn2shAhILtA8OzPOesJAd9wLxpz95y1Y
IwMzxRwKCeUp7/WbYq8Ku7fWAFY5Dobl7nWD8HTgl0ZwvPgmqSniPLXln16QMlCDw2gZ6TNMVUDX
emvG5TOmnlEfD9SvcUnvr2ZhKzFbWzZtjhfw73iFtEdjXeq/mph/GxKx0dCJB+dCqiO4QVLCcDxO
tgVQqt584Tbi5DoMMrUc7xiX5K8jm3JHfEvV7n5FNOXhLQue7FLFohilZDSyqlwXHBohJiMCvEGd
FxvJqjEEARbjLuci2BdcDSvolhV3nAgiBaW819bI5W9cmom05ekLWsS5ALCUdXtIwDMSJmeWGc3E
3ow/H8pJl0Xxs51cA93FZTHlc8Bq8Zt/vUIiiRIRd3X2OxUCM82Qdcfqsmx2szfyhGUjBUpEHgdN
VLM/wPjwStg3tm753csftRPzsJk/YqegvYF9JCEP9nt47mAkK92iLAxedCJccqrhnqgyQUZhGgqM
uzAnlpV+JsTUHOnuH9rZ6NTrAFDdociDwLB9w+yWVJ1kS4uqWhzsvKir+ondMZRQYsbw6qn0iZ6b
DJh54zSMvWOG6ngf1P8ouNcCPxCxsy8vUjcN5aJR/0B4Os00LLXxRMQ+wdZ1WuI/R+bfD7YeAyu3
gjfC+46tPeJwTMeieuJQlmo3YPDLnsRBecWR3O0rA5RanMke6yfkZMGZ/HiovkMMvAOlRPHc5GkK
CBtxWJkH6lW1m1E5MPdmcPn+WqOkZhpZ4Dnum7zv5ekrX2eNQX8A8yj9RUgaOEVaRsg3Vyu8lQV7
luF0/sVgKAQgLfjisjpxBXRZu+Fn6FYfOlzd9q4qFjSvgW9jAHN1i07lDHui+WyoKeCGM3i6Qjft
5ctmHuB9imyZBz/vrPJSTt3liUsm4iPkMZ0VhpJ/EYglXjC9ZPo1Pi7tOqMm0yanGQvzNcbv28ga
1b0dUqI3SWYRP4rTbJ8ZSoQ4ofb+9s6gJgXJXClmPPc+Sa/8qaBKVTAdzjTM/cdbIn/156FGXDLV
rBHW0BP91oJv2nw1VVX+yCrVUtfNtaIP37yInQkj7Zv/gTA3Rztcdl+9FZFF1Vl7UIS6RzYcMQH6
dJb7tW8QXsIERmfGZA2dpdFNZZRu6ZmBnV+caSK+b/jGC/4mAZhmONHLiBTbCtBgo53nWwpACswH
nFEDEUc5egsntO31dhA2N1uXnIemRsTPX+m0+0SEILvcS1xG+NZsT+kr14OglO/Q/vCHZnfv+vIG
UtryxU1K6qN4Uwmcbp7g0Fk2jRgVgIzByxa3f69xcoyQ4HhXz3d9b6vsmv9THl9Bl78ixAF4ehIo
DZpQITYiQBNd1jmcwhyCLV3IQGAhY5XD2ByERa1x0X20lr6qd/eBwf4StbrWfITgUWgzICYTslUm
lntZ6r9O0X8Ny25yqbJ+6CpsY7LJ2JMCZeF6stpUCW30V4+3yU+HrXwIa+5wfzl7T5nTtIwFOTWh
8MJP0jj7QBBwtPYKLMB9iqgwMfA5EhS4KQ7Sb3803y5Zt0YOcgPGvZop//HgJPQfz5TnBTGEItps
QD27DHGR3x58YcgWADV3EMGoHe0o7bL/4u4rWzC1J8eRoAwm5cBOhDGiFdjPEVwpaHQzNhXacBSR
5lYT0ArpN/LlfB73tQ6Te8JeCD9p0HIx60EkUHS22AntNQrvJ5vIcDopixhjcz19NsmBRPj293NR
lSYNR+MlqcwgBjRvM3wbmCamJcL/1/hQ9eMYNDxCi2l5Oo1apvoQwrQZbEepLt8K+0H2pMSn0Nfv
BzKOZRoYepdJFV0Q3RAOZF0ByQqJGda1vSPw2/edzNhiciCgaCzWkJepDRb4GZFUHMdDiTM6Dnxt
itW19rONAalety27q+S8XizYaFrCSyFzGx9nSi74so9jeDkST2y4JEzciIcDMmSWCEQC8WIYJLjM
bsMGl3UWE6yak/3rdRywBKCZ703FD/ZkzuAEAkALLmePNot37ymp5Aek060rS7ZE1wkmJ435DXMX
XweJWBRhcdxJBCLROX/uQJsVGZpAnd3qu0o0sr3W/MzZBO9ZbB+G/yIk63yLXaQ8GzmR+CZ4wKuu
8ufHnNOsWTW/Jv1/rMsGE0Rwf8YJwk96VihvTp6Vplob6sM3etr5HdG0QXAz5bhFlC+1dzHQiy6a
VezKs6bWuuxdOV4Z9OnyzeMGbHHBjCJAvPWCiqUqNaqCemHvY8HeSuEpSom8LdjBvnsrmreNpmJ+
a/wQqYmKS2AOytBba68cJaWuz66pxVfnnHuJ94n3rju3Pb2FY2LBb6HQCP+NHSWH6sclHsGkkq9f
R2Ce+YJAclXYrKtHqpVKoeCNL1w6u7gnVfHGOKtsD0cpTBYUqdQ+fj2vpo9iiHFW7O0ISwadU6lU
/pEIaUCCL23pMXiffcpZ6PPNkZ4A5ShYd7wu07771R1WlQ85sRpDJr2jYrA8t72GofzwHiGtNsQW
OsoVijeV/7H9ouBiskYYtNgWHlhUMwTTmyS2CpTM03mJPM3IXjOdPBY6hyQ8obfgOrgX4mZJNEvv
ggeGH4yc/rK1iHaUjnN/gLe4VlIsrfoluCDWib7KWKVMuLZy246IWHxZoKHjNvX1oGgfzsdpzHUz
+X/wgK/Mm6bZBzOuVTi5+lNL5eYe1inUO68pSi5Yu5PogLDNBkC/TwXtDw2xI5L0DWiD90TTqn27
8yAu7ONc3uCfSwwcMGrIRTNSXNmErgxdL0Y8qVDl6xsMbGISaYNzl3/kKdwX/8n/+8CewoCXVm9J
LsNrlY5v8vxAykHM38Djz+W/Z1i9QURMzWlwN6cZBVX8mjd9sdyUkk1/Rzgl5KgCFpfW/0xVbppu
VoqmLGyO6t+Z5flDCnK3tz9eP2R6P93qkKBS8pyXk7TzrRe0h6Cnc+A7VNt+qQCxONls1jnkkF4+
QYQhKYw9M7oi7PWSrBumnPScwyrFO4M/Z75LkrrziaUBGxd/xS8sMFnlgVmFhzZgpUaDyT0paDis
GoCJJyOxW7CikB66OX55jskdhNFglrppeuutqEpuMQmT4BO4O+DT0WbqOEdB5UKDjmDbcR6gOHNe
jCxX3IthiAV0r5cayXaeA5ej5heN8ZH8HF4uwzQvA4SlVwEK36gCqfme2tfuRQpImMNT4N9iD2dB
IrD+VfVIaWUw4QwmFhjeKYkOfs8grGYBEWppW0o89apCOZvqTq4z8+Qh9xteefQjoYRPSEVZBuK4
GkXEjrEfpCSyZ9Hv0sjXeSKHa4qjwl2CxdwZzjd8X14/7QMIoDJNK8m5KNSugDLllJCSLhYHuld1
3dt/MzDNFY1l6mIn8nXXy8/LQXdU7BqD8mqH3wgnzaW5XTRczfX8vxX2d0X91/+BcDje9Bhtygjb
5xXflwq0NdUWrz3v955/G8MhemjudflQKqU7zRE3IvTdCOp+M3YtyQ1l4AOcQRUGpSMse29uyeBd
o+kfPDxzdL5PWihC6zFxwsBTbbhANKbFN80YlXgSMbBVQJYp3MHGHO+XUo/2k7G9AI0qZgkVGvUM
woP607MEArFao057wCq5gLNc2HNFjzpg4o8KFDI/51d2oGJWT8X34H7Jmy+/RGXxs/rkDt8wzRFM
Vm2i6GUTxWkrWodT8cB42bXu1iWw+QxYZlszTMDoNNuAfBvnojgtvxPDbf6n0CA/8RrZI8ydAH1v
ovkEdERFCGV/TOzBF0s7q3URwYH6qAhvt0ioScyzOHKaCjLHzKR4nxw5nUcsQFakhaZitSDFzGEl
elp2gcpiWBzaFhrpxRfsuAl8V924dYLkCdAeC+GMoiXVxjJ7+cJ7GCPSrnAqkkqxoEeUcsBafInO
pk+L0jNTKZgYwmEyHABOuosVZswwlXS9jKMJmEtI9obhz0gB7tuY/sYLcycmD45ZUgNbX4GQR/hw
d2WQm3NanqbTt7U8bdO0jnVh2Kjo2KkdIZtVJ7JmDjdutYpnTe9/qpfn+LK6MYEYfI6AnldFxYvA
/Js0Go425T1HtFDnmOipoiGqRCvH64rb/+UzPhAB4VOBnfm39x7TBTeufuTmY+bS+UfwF1lhBC7O
f8lpkLWV1cBoZM8gc5DhTEUhdmYQD82U/J38d+HrljCWina8/b32J0B4J4tI572yIlzujZ2ELT+1
ItZGjqocJICW8pHEKX68NCHbWkCmexrbhb7xmewmnRX9fuozogsAKT7oJOF/AUIm833Y2Ap+M5N7
QhxUSiWNC0Em+sIuhcSulR38KR/x7RXHZnv4vmm+tS8yWHlnCy/KArOk1F7QinWCCniK71ycquMZ
Rh5AJtRJi03XB5QjCW7rsbqVhZFg8mNFNmWKLv3+jBaboDiQniF7X3InQRwcrP4XatnxJHMstAqc
kf+pADLaH+HTels83yO/HfJ4a4iMRwP7zpQygDlV4oNdmtx3kdoL3bb287R1AOaHPVNFSw7K8IVj
UN6me3TK2GzQmGvCGONF1yPp7HYNkdjfLorvvQUXa7dU3L6NKh7/rtaJe5k8ZU9lqcu5xyBWm0Lf
cWjm+7AvTDG1dZ3y83e8LTrjjRjMaalpEKWDOnq16kP8bY7aRZiBKIURd7gM0YIUlJrK+dUIrJkd
8PrvW7v4FV0aLpxc0lDjd0l1PBA1uOoon65mRncPha0+3fZuskTMb2ydF6KQ8BQy5JLuzqa5SonL
UErwEiR07nh6tcW3OadYj6ALqwXqYltCDUtv76cWzbXz8WLWxd3hBNcl3nbgYElJfp2EmmN4FJ9a
vCb6kLv+6N6mUF3FyZrTKxRqmxjHiOw/5M5JA7kxEOK8p2ng1qCCwuwxB0157nl1uxxGShxCflyL
TsO4uKWtz7QVDL4O9pCWkU2vPAR5X6izVO01x7iSlICIfsVuEyUQ7XQ4dBaDAZY3I8jRhMcG9Zke
InmxuoTzG8xcxhDi2LB/OtKAD4M6kykIpSX5Eb3k/FEFslrPleTwPiBC6urHJu5Kz2/5pWypFiU1
MymbPW6ftQ3IjLlgWdNGNuAAoo2DIBUHBFFV52u4dfnpGyQvGcNQN2ypxl5ZWpZgEkB+qlgjEKrs
jVmYmbQCRFGF+Igdhm9vlRatAk/jAsuDNeQ+F3otGyB8IYrmibK3ltP+66Qqx1jfqhNS3uZR4/kO
S3tx6OQnD1PxpjspgXcrl6Cw5SCZ/VKvTAbXfMgVRr5W9qCNFM2tU0idsX68wpgn6zxfz1yustB6
elX8/LtTmXafd63G3cDGfZqZGETZIE7MpcptqgbvVSyaCfmPDgo+QWjzJktzR+iMiyj2ocoqdKq7
rBWujCgOAU+eV+yWSkLejTmpQgFdD3/SnySc94nFxTG3tommdC0CCRRA3kePdWOZD740tpQxpx6L
8atYFKTeYMyyq7IhdU3P3GFFrrnDEDLGzZijJAwy4iKEiuz85RwbgALV3mNJJy5/RLYg1yAQn2W0
aSy7Fqei4vux22f+EfSx4X+gUttdWyzPjD9OCtSEZ+3C2Nqd1PP3ryBe3V+/nVEnCTN4wB7xMOqq
xTb+86wTrcu/F3Pa5bl8hblxpmE1XeWe3KxSQLv19Is+HdqP2wbM+UYladqf8tOrFpGHTiPVKYWq
jLy5FABOHUUlBigyKn6eTBAGlej4PmytHPFQuUhfm43PvRwUR5m6dmtDqL11XpyrXtdiL1sxDgsK
zjHMfZh+BGQg75oWUBbpNrhBj6+KM0Qt/vdVpbhPTR+NxqcNo/sR3/fBcLRvrenC2X9kZ3pj7lLF
dLOsb6ZbedmCA4cYx4yeaNzrgC7pBIh3tIWjwwsEMlvYN60iXMO6Y+qWwRSsMJMI6G0OjR996eWy
Jx0WKoBXveXSH/200Ba9Afs/tK9EB1PlXo9JxLhrrikS/PEHw2KkZ56Rmh41fm/qKpc7HpstkIvU
e1V9VUc1U5vgMGJQAX34i7Vx1ayeoNRI04PZimzJvf16oyR4q5HVW9Z8GVrQ4o3kr8lPMyaXDuQ0
urqktGOF4SFe+WrT3b0PvKBbohPoX3dGWIV6/mvrG+ranqHovFQ/fTR3KRmfpsNL9vE4ik/8aq5Z
0/2jWKqdoKvIGfE3hHXS17m4Dp0X6Cr54KoC3hlKybSe6iVb9G7J4+2gmMV7yS+s/AE2IyHQ6YGz
C68lQJ1gBX5U2hOTDM8L48BGBrdHjIEHWMcXAiThTkodpw8gGtYTsf3/mosnuRvQM09yzhCc2cDm
p8iDLD0jky/LeelePKT/50pIIzYv41fvJ1pDzqe36HrcpE6zotie6K5UKChEDtsPwiY1S0mL5yCZ
oP9Xw+fMr8JDccAWBrkrwaDOSeooDGFSl+LYzt6GRED+o8P9cNh05NtYLI4mfnDEzdHXWzeTFpi+
Rhj+dF8MBZ8eyCyNQfbwaR147yAqn4w8D3lsN/gU6zH9Ir0gFdfC+cNqp1t/e5AoShxaFUU1FwmT
9EguyKzZw1OHQqvm0zq1qCKhC/XstzFxn9qEVJQBN3APNFD5DwTvx7Agdk4pCng3FPYXqOnN6syp
If/UKuRQYXXQ7m6N7J7trGM2c/j6jE8f5017xmvJ0KUqBu6vPtEeU8y+Wnv3uWg2P/MkgshrRb0L
pKAgC3QS/u9gG+kV7b/1k7RyJik+WlLCA5Qh/qTGGt+I7eLQbaf/bV7ktFxpHm7QvZR2xshGlcNs
R/4juthqMLgB8tT70I1dTBc9f5YCOE16H1hb3CLhWwAfJKhIOz0pYWgg6fmRi8izYp8ijoVrr5vu
blGGyRhT3TLUFI9IYhKiaNl+FLCS0Yl6szxW/xu0fCUuppiFkmzlc7VLCgxgqbbM5QFY4I4g9ClH
rN78hTIrodRTjuDGj9IwO2u4ZT2lkcvks6V0idlm0dhgAqSUmN2jgUfnqNHarYAIFmu5xyMeRdcI
ZAuO8j5Wfs7HnTlGwpxjgZ13tWXxOVyVLmC9p1whe+Yoy0TMf9j9Naekq6jT0M8Lw+S7SNNJCqZz
j2/r/ybPB0DnP5WJ7WKdGBxt1IDUr3W6NdinGKgmJUC5SdrD/4Vcv6l1CQ8k8/h9D27jJ0HYfJnD
tJnEkRL1aTscnH8dcY3qapPiSBdu3ZHNTxATD/LaKOwRTpTZkr2ZYAbW2eLhhUe0xokwiseLrmMk
ZYHZ5KtEjVZ2QrrzL1rNRSZ1QrBKhtcewx5/GJ13f3heDMiRcxc9LZoNO/v80Op8mCrzKfO5qkaw
1n1lqByzOEAJm2xQkegjFNJ72Y+YaAK7owp8w5NH2NyeAa3i8tWQqWjlHpW6kM5ncSR8xiJ1JRmB
CrBIFaYbcZmkepMfNtKshEuWa9DcRvsPl4Y1KmOjX1D5oVbe1U/qG4MrGCjjM4nUS7tcDv5khl2B
erL1gTJpf3yKg4UeOWh9yxSkTOjyZDsueMrLhQTlSHuxOlpv8JtJ5AX+5FG2S5j7mo2ptLbmxkYh
qJlZ3Ybd/7G3IaK8PB/mxHWGTI4Sk58gLuYvzn9l7hw+E51nEnJYu43J4hiGZtWJefa3wlgE/gVF
JCKPugNQSGamiJDBTLy1+SQgh/f5uHAi/QMoTZE30BTvaYe/9vBmVCI67WhC1pQaVrXIdu4ZQj0A
zeaTs188ks3a7OicSQculX+v1a+aA7NxXDqIFO6jrlrv6SRbqgNYEl6wCrEukuuf8wegCyqUHltm
+yujb17GujEVzUt9yecy9Yw+C6umATHagYujoFfLOhNkXcSXBF8A/X0RQervNLIvYYUzHg+ux3Bl
cY1CS1xTqdw0XmBhftoQKeCdq8HCL9U32RYtL//FHXvUYkyX4+ACLoHG8cW2kM9eOW3o5guThERh
SdxLjClJjVIt1xQ3XzGGe8Td7or6oJEzSGOCT5MD0AEoZokgks+2dKSezQkbqhmSDDlaUkfqfq4F
O3nOCThsOX8DRtgjGNy4/O4jTWc2/8bp4PjQzt99Drb6a2MnwKGk5ewADfWNHPCPkXwlUsZRKR8R
jEyWtqQgrmtYPZyASyTmqIaoTjxlzs4/cyz3kFVauf3mc+tHBfmv+9MYKcpWLBKtBR9VvmYsAtXR
djuFccTH814qW037vKRds623jpQnR/2slAPO0LMkXcF/MDL1VrdIefAHCsKSjbV0kEgDjfB9EuKQ
hCOYNKsbFhHF57KUGvp5+C8yZrZQiHG+qc4Hoevb5PJW7rpeyjQfDIJzWSu8kZRF3NcomZ5ZyXBU
EKFu/P05jX7VJNFszSOB3se7VPtP2fH28zamDHspd+gGwbBRHq3kY00BV7bKW6aBuIl9e/X892BH
g/aEGMu6bqnorCZO2c0yjfhFfneL1xTpsiGNVlT2OQiHjDI9BOZXh2FGJXXVSlljv9xFRayXN8q+
ukAK16+YJHt3cLPtKd42MemQyaG5cWVgZjzpMXoT6VcIOb4nmmrNVUZFU1xsQ3V4RgrAqboHc0GC
D5fKvazQ20CSI12x3eo1VBYuc/4Q3DTwTj7XNAuZE2hFQd1JE96m/0CQv7JFJ714rltpCy1mo2Ow
CoTBKseZ9azeK0i/H4CsojyAe3+F8oAUmTlztJYTkV7daxR3gcH6h278PKyauHhkIlwjVbLxHC7p
jhOQnzxZiuUsc1zjLNnyGo8GMaYNlehzI/c1NZySb08/r5+B9UXplO8n6girttFnxo4mq1Ugt5fv
fdPuzzkyP8RvJbffUle9oDRBhq15heEp2z/Y8CKpYp1yauyDucRmhbaocRT6MT1Fm71nuj07rf0r
pjNm4E5Ck3vtnG/7OnDm8otNaV5B08pPMbA167xBPMUz0lwG88Ty/ZmCc/dowCsWAhi3sqIS0NUn
CF4n2/biHlC0LSLIA15yQnpzgrhEKrwAEYWZmlRiNOncQVu6a163/WRJmc4NCMx134RBjpZeihX8
yhAK6ouZDaoE5M8DjO6tNUC6x3XHcCXDgnAUZd1ntTW+i0PvHoNPLPBwgjTIZ1FPVCqZG8Ayh5D0
+QwPFNkZr8j4mvmpS+5ojQu8HQU8SewMIhdrZHSXgVyzzIkO761uZNNVtrCQQ7Uec1mFKz1BJdbO
Cs/lRFULy9WTZyfAXhKrmVVnlxWUKoaCx3aZOZNCnSJLHxJVUH6OpQ6mJbnN3O2IgKiQTM9RII4f
N44F140FJXrx5DF4WHmBiokLL3eZiJXz6esxnq7kQeVpATcADzMcZ3B1uDXSO0eJ7IdeNFG2Jw1f
vqPcbAbNexzn+B6zDhT3bh9Ctqj0CD6UgBJUnjdC7r25XNsKedazga41OHa2u0ZbT9vJbGSKsrLS
VhDQgqe4AO1bZFpv3TWjwUP0biJts7l6qPBMYRFSghutmvTIDV3mK+e66sv6/zhCof4AHSfv5UdR
ig650eCFOa2sIXSBE/20/4y/vlm16T6VIVZqofIO2Mu8HX5P2s7eWrj+OOttc36U2sEvZZRQov7X
xt1nwDP1Ilc5PvXf9pJCITioHnU/ouM4wBJEiBekl89/H1ZSGC8rnt0PYj6Bk0W5dTMm+bag0Fe3
UjkwojGpChQdd1Cq8A7xBe8AIIFAjdLZulvDZ73XQmLhg+fzIHLr10lownmB/t691ksIHkdee/H3
b+PBRkZNCRLkIg4CuRum84/dB7krDoh9/6HfAGbL7tIqYQpxPSBjjAbFDAjS9C1CYaCDbTl4CT7w
1q55H+AKpaTQpx+nCu6ZVdox2hkBWRGIvkn1epL+QauOFOPWEm4R5gStfTytSqltV+NR0g9n0dbj
KU++dghJWyZUEjSfDizLNALf6KZAOIgKRlbKY+Ju2gDHcUliGVv31WyLbG4ejPLNGRiDhsXLWE/j
x+9q6T2TYhpvxtWi4bzZFF3MKHaWPGSCa/aXG106/lEA7r3dpkiABLDsXcBKyBwg4CTf4rZ5HaQx
0tPnf4rKO8sqBdKPPCXcGO/kEIQv118FE2zZ/cRvkjN6KYO2ZMl1B/2b3Ug09UnfICZchJnOCL0e
JAONOTPWl1TxUEbulW29lOhSY7c08xX/HkB7JgZ8EzhwFpIkZV7peBcchCYE6fSeiLGTgjv/nVUx
X9PJqvrbEsJJVrvUrTCdqcYM2VYxEaVGTPPXaNA1xSPdwYlJxpwZvdC6uqu7XEW6dh8KJqHPR7or
pUHArtQS49Fg77WijRSZGtmC9TwDqyn+CM1tMy02WoBIGo9QeHZ4T7FHTkB+v45KzgqkNnyk1NQi
yfOtyrnVjS9NUYqZ5VKZPDB/ENrareF9BfPGN3zcAaa3U7AouxevWY7AoTogE4D/iSGcb+5DVR2n
6suaqFrQDDAg8tEoDHV3i27FwB+k+EVwQyXd5AeOY1bC9vy8F15l/LqHyBYWedvC+XmjFvDwvuc+
oKgq2yMagk6dqPNechU2BM8fUoDzkSFUzI3PP4dAUAjZLi1axIIz9Luh0OGenWK22CHsUGxfzwdx
AAwWgm64alWzk/s1Lt2HZTIL5XWvRBp5lMfIiVSXCr43NDQtDH+SAssHeQ7zGrVxBJu/uljbxNAE
5/gIcvAzM+iB71AQ6xba86y7oFj/dLnwcNtFJOai8pCuvPLLpD15+xddDCagvM/OH7APWqk/0nvG
LaVDtHXp1DnOcPl1GedrrbO166M/sVSvxF3CIRWTvwaP0FsvQaJlucwjiyR4eozCsSUTo5BYSy3s
GGHyKrYFW68gTWTVsTRoHYIuBY0YX9zT6AVPlhm+FpwdbUTYcxbLJE0/LOXRce7nRgcTe6DjSQ5y
pWYmg5SxcIm0WAHkeNreVct6UkHbbVnBnYspmp6POiPDTqp50LO1DMUVFWaqh6qPlrZrD5wUHJPk
8xwI0myoiNcN0FiNtAnmgiQclfMwQyUr0UNobBijy1NfglOqlI2J0+a1KvRLq1ZtIlP9bobs44PK
UZsDDpKE9OBg6vFP8Xt0Iwe04AsY3X7ZybGYe+1sKkUmqNYpEpl1CDaOUNvyYpDmNZCfz+W3raxV
vv4FCT5EN1069G2uwk/7O69DYCkQ0si3Y2C0HF3Qmfv27GqzbBGh32LLFz5y9DZjkdkg5vg5ETPL
pwH3OHBbC/TAgh8oX1CJsg8CNkOgI9UiaRdQxZ7KHedDoHw9jzVi+jtEbJjW/x3bNDBeKScZ0jft
FXv9dLcZDrf+gB0hS79ClBSe4+ZDsnpc1CQI4qrPMhGYzGt+4QOVTrnhpDwRgUhTqu98h+Eb5Na4
xRLcCMo6wyb2nAyO6DQHp6NGFX0ExyHugDp4IcMn6Xlld7PWBdnO195ljhgOdy1ilEINZs+M4qIq
sfWHREiDGAkSRw2nbC8np645KycTKTHQvH6aan1uLtYvV0zONiUnzf5WrC72cJmT2Mrx7ojj/8ut
l1SFdeTVS9jEQHWSUpD/8f+2tT03Vb+va3lfCk5+krn+lb3ZY4F+UUFv5K87LLqkmVfBQuA7McG3
WWN5o5jTpYf6zG2GzeI6kUREfW5+FxVfx+FB8IQBcHUFeQJ0pVBdUNSFXvB2VmFMdrGEYZcmoqx4
sdX5SI76Pr0MKgug7uPPCpL+jA1+A6iwvHimvnO25DLhs6JHVKK1/n2leRP/iXjIpta6e80rykxI
FYyVg8GuSc1J+7EmoMlfNJzy0IVB6TxmkOx55VlFacOBXWp8c7jwd4QjWz21bLKtzTPqY0Fsmg+g
5gkq0/pPvRY9Kn/eL7VhMiAEFFBnA2CLYri+c96oAo9mYaHoIZ16LPiUW4uUUieNUa85erIx3gtW
RIdPiJ58sf/bkqP9VCTaHucnY/ymT8PNd6Aet4/lAF5ubMdFhc3U2ILkN3yhO5WXfifyC12PqGp0
FY5H3o78HMaUC0gWzwi47xqY7etG5aB5lA1LA53tIyFW6ejzXE82tNxer3aCW1OYk/HJ9SNnqCc7
yggWRCbCALLRfTGbK7Oi5Gfs0A8cA2WJXoehYtrc6tROhDr2ugTUOlkzEentrG+9otq0oDdRFK8M
TETxgHZHY3e71cemBSBd8oT1x653QpFWVPpMliu77G+FqAMSVc4rHtF9Wc8KEhoMOLpt6FcYcKhi
EZaJBfNx6GfHOgtBRJR6VgF30GUDX2qcC4qYjklVfoxCDwsie7Xr8rbkh7NjykA1wB4T6s8zU5Oz
JCSTdlmpevbWEKARDCTf6/BUBXfCXMcmJ8HScH6a8J4lRyV+M+B4o26JuAl4MUBjKy9cBoUWbxZw
c3RQlTmDtdAYO4DIqt4JjcefaBSZNQlEClw51WmHxL3MqSbPiVutFWV7U0eY7eRjEKyyKLSfv6Hd
zb3/wEaiK4oVvcEpJNgfsYCs06mWbDfJ0nJDv3vLjwV1Y0XxYryJCRTPhenQ48g3iOaxaFFJBCQI
jH5EyTBd8acEf5zKaJx29+7bPzd51hW43kuq5gL0l+Ex2xdqeqDFDNtcPdezK+0A7a3ufF0+jEEB
oGWB2zGmRcjNr1ZZf5ezbndVPWoDeNxnQ7zjdxFEFvbUAZt+kMq5ARyIm1P6wGX2QZl065u2B3pk
w5YXYht9lgzDK3P+ePJg6nm8ffHU2Y2GK4rufbfyibCf9yY9MWlDZ3nxg/yktVzHl2MPHFmyUbcU
ufFkDWToPPRYCI0BAB5+JQxPl6SEfxUdTuYBBZ/0lxtxoNZ7D/3Mx9ECFTm6rpWTVnaAGEUoaiyA
9j+ScE2+U47lDxPAIzHU3eP7IkmufXNf7Ra1HGb+mZuvs6tDvYgWPg5hyJfSmtQ8mie/L61PF/Pe
Ljj6nERpaMJU/zPWbfNMtKZlZ+2O0oSjxSpZJh0ClTjfc/uKL880NC+Q9AuINtBNCIecaxPqzOI6
eede6AoTXbsJFDrgkcCq/KB8EolwIG6IHMGBO7XS9p4/DblckEM5KzbwW7Ewf2a0HGw9qfaqyika
wwOQtSU4pGdhFvyi4k6YRd9U3r3RcOoVVSd6qWXj4FODuzO3vtb7oW6R4F3diuSP05WIdbuJQggh
7f5MbNUlZkk26jFG1qmZ+KHldwquoiZ0A2tAGj/cQT8VRYCgAgaUPGAPqcPlcCmhC8TX4rft7jDV
csNPvCw10HJvshRdCrr3F/Axk4uSdcmr42Q/c+jW56ezc1Oa25n3MJm6J+n6lqtNQwBihbWv41uo
YLs/ZVRL2/iGXSdHXqK4tNONLooiazOK1GTGr6Y3P5nJDpjGOV5p5KFDdEctVrp3mQMgquQ2jdyK
wr7z+r/rFD4jdj2BTvUpTLeHO9v5afb57jC5lqMCRjWrLtqJrfOfsSz4Sms3/Q21kHkTalEq54KL
XC/KkjIvmHG/Uq4s7uXNv5Ze0V7hjR7ZAAzm/5PDG0AL9F1zN/by47qaCP75QUJQCIA/feK5LR/u
3JHpm/aQ9Ci2P0x1txPJLHehvLa6Yg2QsYyDKI5uBl8y1PLqOwR8QHP1oORZnxN59IXgU3NWEkom
mnOK6LakYu+jIhkcHMToc792PuxhJra3ck7FWJoVcIHlO2kJygumuUVWtzQic14yamwKnyBFxmRU
svv9LIrcVn14EBzv9Fo5ggukqGeCvbZIx9lTtpiq/nYUA3czAOnYe6TWRmlNbn23VdgYMIbMZVT7
qAl/rSUPTQ+FC65a9SVNRZLWtkBmr4/9R3MaetZmoUpIvokbUylRaDoWAaBFQBT828bSzEvtKKvY
NdtC04/P4CMJnHPTrT/evhqRec12RMn+GQJbeN/QqQKAJxrCkP6jTF27Lc6d1lTsQCaxbDgxk91i
oHnR1KOkYiiw/+UPY5irw+PGuyjsMphAV5muixCPBxzJP+7zsLKzPSYgl9Z55qUu8OLamhDA/4Tn
5p9XT9uY0JNv65QifeIJp2RAAJndaVSg8C2qGaII/iLLh2ArxDM9seX9YN0QiTXfx3GZYE5zeUPE
Ug9ecPoAmiMilE5sbXkxwIKfEJy+sIStDakpqU4wkIOLkC8FFdmXEa2ZjwktZkrFot2Xh1CXvaFn
dVC7ckdXtjOvnsLFf4+bBwL9x/e6tCznkrzbrMkp8N7gGvBnH/bGnmlAjyybnrcMSNa4f7arRSw2
aBifpE44ooj00p8b29ncs+8mjqU0VREwNFQ3C7g7CzqVJIh4TZrCo1KL0gremRq6426CgBUyFaFO
PMuZtxypqVX4NHQL8YFYzYoQysSPTDY01wMf4U8XiGmeKJGFq3SHpBeDo+OJn1PDo+eA3HlvtyW8
AdR96WdA2a0oV98Mlo7TVqtUBFkB1m7a9aCMMzP4ewxVWmiecWcgu2i499zIrAkqm8uJuYcCgr5m
umdq/+htlGcqzrUDAdF5JQoX+TiMW4rWy1Y6HrkOePshZjJRFXwnjpg1hWOEz21fJu9EPw+OwhaD
UcAJf0T/Q8BxhWS1MGe49GvDNjKjI3X/fp/kDx7PQrmSlD9dn/jIIbwPNP99u6Wm0VsZjHo+2GDd
rU1yd/7qQ2DZwBVI09VluxoQvZpjkCHO6cRkpREQ+ZdA5XTk44UVnXo73SOa8SaSBL0s6Pj9rkpW
C+NlTqLrjZtdbMHQSE9WxSBsnckccllSrmfzo7di24hNlTiLe3qBDFj2MgfliE3R8xb4wwkoDfg8
oCoiv3rofhWG57fYKQ5jUYP+gJ5Y3uk1cfzbraJAXoTsyRBH0THJ/QC5zdAfTS5r9F9fBdhD+4QX
f1sJfFjh4ZfDyTo5RI1CIfeu7j6y2hmrI11Xh/8mhN0LvxFtSWh4BE55ZUdfxbUsDyiQl74xcINh
ndRVXD1kv/iBMicQxM06mgLku3hiPTYegx0KA0sn5Mj/SyXKsJtb0kf5UpiFg25Q5esYPVcqX0OZ
Zw/OELzl9HG4pGdg6YvXOWYOg+/7osnLv+eLNN19tgourSAW4ImfQlTyHlQ7BOGmHrs+uxYfE2bm
tYoznoHG5Wmtg7HtDSefJMuCgvyqIYA2oI61k/kyqgriWWDsxE6iWSg+vsBXMT5thaSo1m7b1IG/
SRrU1MyYwzBFZ1KBHcs6r/KPSek/luV+hHaczVlhg6Opx87yyf2nBCEC8L93CNrvQhvksrwBmf7n
TyGboai6xHf6As7Q2XGUTdLetWgTyJWCJT/aA9pWltEyJQpa3k73O0sMJrkyH/PSFZjjmzHW+zhY
PAmxIxCZWDwkzH7gFxrxc8xKxiKJazC8UqzWFWAssWGmBzpuyDlrsf4s0Z8n2DjM48DN3tObJkMy
+DfOmkmXHL11NadYykmM2wEcJL88y4dR67t7WFlZlzhv5kH+CoCxcn+G3OSzo08rgKsS0WYAU1k9
NPwbOh/YT5qJ3PF+uRHj3hDjzppi1l+hMwRSaSSudhUO3BiTh+qCPkpt8ixxYDyzNcH6xuKXqSPI
AAuW6Zw4LNE3k/JDMI+gaMFQkPLnxmGZ3ZhJ+8aDks/Awik7h5kFt8FQbwTWUL4MxU0R7VFhq7JJ
C+KVrC+UT7iILCxXrfiMNE9gFut+gEYO2Frr0fLq2cba3loMRSHmFR5+BHsD6Q5jfabX5YiUjHPL
rhgXMPS9r0gDTPDvWE25U1xcDd7pYVzLVJMW8aLJbeQB6qlHGgQwQM0thRtCWfrIA5KWAGs/STvC
WzdFjIunSaEmo+uKLc7H73dz1zWVVyiy7OV0zoKDux3vJ0ikc1q7ZNt9OIywzu3ckkhK0YzN732Z
COvM8fXxR9KMs2Fz1DTnoWMAMHBJTNp+lwM2nq+GIzbGATWVChu+vYUXbEaBl1t8mSCjpA3zmSl/
u7sjztSkgKZf5e+GaGrMetqIGh20+1imMpNVfhop6CBCyLcMVQPvecEe6VOTEJgjFztJPuRe/by3
6JGqW3lRgEM5Fz/gI2U7oXsxt/jhOjYI8+rKxku4nr0eXTbjILHxU5zrSEfi0Y+Oz4kFwX8Tfs+O
vEVgsr3+FM4CynOajwCftnb590b4e6LtmRnWmdh4ZWh5kCS+KzY4sG4YNFbRumIaAiWonfv4EA2Q
WGoNFhBxjCxoN3gLtg6O+N7T7SkHopLkZonZQUglz5OnpzFDadg0v3iAn7wIsqmU2nSfroXME+7g
t8CZ1WLheXHjErXTw68dQVxoYloWgRmOtWnuS008XWuImQ6CkmSwVhPsWQWscQZ04JmU+ZE1xG97
2ccBfulekgyr10iZbTQ24ndii4BWy/Yz8/0QMIPY4fSJ+Kj/6WCXmH8RSyiQyLDRzT5tNvnqtahg
vz6lnRnL0xh01SFtePUy4X5QmZDioxriSPbkIUO0J4AUSPMc2urBhUM3j5ZIpL9BDX/b3Wnj5um8
y5cSLozSKgomfpoMw9BjuhyEhNzGYvFvN9ndHSZ/6qNEXQDT4AxG1yXtJRHsD+JBz+q/wdBlNYEk
GAIVPN3VcUIqxJdOQEkOopLgARfiCkg+T3QFhQ9ulxEDWUqQBdTzgPsfM1XdkSED/OohJdRk2p87
WVWdY1LuM5w8fKMznccY+YSuLClWQFw0ejvExS1XdP03QzSRO+hzQd05zKkTYtuAcIGfypXQOsdU
qyo+RcuCO31LhPjVw8NYZ0osQCIYVHaQCexp+miedro9Kr0OaMgNJxuoaUBrCbej342I3YSIL4Xx
kRLrUTAxtB3f6vKU3GP1RhlJk5swxqqTFNjPumdhxV8aSsJ/7U9Sruo5JvIaozikWXgAPWMhEFIR
As6mMHcj1Ouv8IDuK3G48uvScIdKLx5nZEm4WS75irTttTkDsznU4+YNRvmKIhG4XkDEiLFtFWV9
co7yYuOqbv1OxmCyFRLGdMYd27y2zpQ+WioTF3qwj4PeqCA8aCPTdnpFcC9lRAIlx41HH1l7EVln
/9ojnM7a18QPBJ4U5Scrrrk1cqanV0GJwcb6cj/GiWd0eEpyTo9v7IpubpaF16g5WtpBH3+1TWix
4YBTq1VfLhtQmysUKD43NEhJAgKZHuyYsV2LkPinsVbt7wmcD675n9tjFeptnQPpMKUdvcNDnbXV
lNCgvCyUdk+NcMcopRa+YVOrkxDxV/QLk/b3p3h+u2J6txvgJpSOFkYh+oz+cvyYwZtZ7iM1yCvG
TerwNrwqAtGSLMU7juX+MM7T8xdO9O95RxyJriIg3z+djWsfsRVMENmSNaN7Htd8ptxl3eeag9Jz
5nXoIMClVmVyzdWNQs1GcYH4kFFXC+F3SxZCh/BMz+EDVycZxBwgJiV3z7fZabzIuQehn6Q7CnKt
n+aELc7e1IIlL7KVFbZLAT0D6ti/FplJLsDXtDyJxDlhRAE/ARSGCi+yL9c2YnElDFuHsTPdTxuu
ma5aC+DzprEJnyEhQSTWcsFHZ1aAFbl26ja8DaR92BId/CIUXz137XaONUHKriiBmX5eXtLWLwej
fTK35QpuulWNKWRdIkKqwN7wiD1VkI4m5xh51VS0D01OqcH//91CLyAoMCRqMBBHb0V2meBKTmMq
5iPrEXILmofqKpzv8/vF04OT5rRPlUC5uu+8TsCVUWgs+JcGLmBCNMhA5LmTuH7Zleznd/RRvrHz
TYd0aoKyc2tAldYs9Zx7iv/F0pqsALbd8AddDDiVSZOcFcrt2WDhaShDOwrzD2Zew545mDmgzo6/
9qpBDJmONiLP10jnaEELZJKeehdET3Kpgwnh+Dx+Bx2dnntimDYFrYQL0eZIUUGgI4sjZI/lpNeI
g43OsNlHWcHNUh2oVA6LKbG92cYjceiywZ7pyQDEoCvoQJhhRy7RsZ2IcevpHAWgwfG1iT/NNKrx
h57FAU4fJurDGI46EQfM2nlLdwxc94QnZXgy+cFrV0RyYYsozMoNdXaLjIoBw8bb3Xt6QgLhhoLA
xHOVhM9J0j17v3xOYy/EuoFkEtdfyXz+oUe2O3s5jJdDTi9egD5yDCohY0B8vzR+UnA1PowJNviJ
6vFo0NSNFrJUP8HZOCxRjndxzZ1qsB/Mp+J/ODjHqHWF2xdzk6RuX3QhrEhzOXJTPAWGG2sByKfL
bYPv/9i+eGr9hgt6grrGaFojt6hkUwhc6agnKN8EB0L5oWl2oRFEYIGHEzpX2/HdpkrhT7sRikuM
lEIfj0El6sxaylgnr2ae3muwSgOKUsiqQVdCgbytI2AMlWx4Tf9wjTJ5IUFXP/SFlQWexsNZ8VEG
Kb06y56E2v3VrikqLeRiiDrGG0o4Ffj/fcrCS7/+ChSGMlcUk4bg70BOGz/sfOxCuB60uKTnwnJa
2pnjjuqvlG3QcUtUcPzwgYsyK0w+E0ZhdeDXJYIfXm8zwIzAhGiMVPxBW4eGHq2Dcg65BeDo8o1R
honNPu9traBYvfAZmaHE2Pye4c7Fjp/Z9uohCgYwPwk5h5v9BrGCoqryWwWNl3p1nN/sZ1Zfz6Fj
0YDMUQC2gE3JVitKXcAFwSZVgvz/W/YhW8nDrOf47iBdC0TPCEpogIxCtrLqoHbXTVqjzcBPPewm
D1VIhUBhjHkAibiBsiAa1HFZL/NRBQOWK2DMLf3WBbSgFLzSUotysZ4J7F+jAFduxtQW7m45IQ1q
ToB5Mkw2aMT+5lnRavDk8jZkg7Cn1aRDMwiOCu8ExVVlyOxO0x+v6ScYq6HJ+djRhxEyXcRNN0Rz
QBSKaKsdow5C6NfKODaAx4FUQFUnxBm9OS1roxaCjGwSzBHJWqT0z19u1bz8Vrzo1m1mznaMoCqB
L8dPhBvoiWoMOqv/hfJLQnAYtwhEk7VEc44oZ6bc8iLp5U04HB1aR907txMvnguhXd6JU1T/cEfO
bR9TpXJG06bpyMAWrQcbiyRj6JK7tmPF4f3tlZH0jqxnk/BerAYobRBdXcqUWTt75/cONafIJnDz
zcURlbewmkW9tig1t8gx0CO6bZL9IK8a2Lw2x0RtUH8ZaHTz/4m3x83tyUldXBE9ukQsnpLugnLh
Uo5JKppFSM0r1KgmmUZDIuYowQ2beMYad6BOp/5pykzlbX21X73fvwscQ97sKBCbbyR3JysWm2BA
/uy0xipMNZr4bOx305yZZWTH8zrG/ItryNeuUdNscr9H+ZBCz/SkoBdKMR8bWiAKE6eTxYXraL81
gs8ShKcgBiWNxKbWv2zFYI+P10IVzYFkDot6XTSTpCjl9YBvf8CXefEz0PTFAvJ37Aw7Ks4B5OiV
lZMp/jUc8b/sWVbXwTuyW76e9vM3RavQiPSD3FwuM1n8NHTT5KpB5evbNsTr9GQL6fY2JxhGxrCm
gR8YqG4us11Oq8VRUFXvR5oNWrICd8DwY8GgBPKlSqF/viZ5V5lc/vqC8FxSVHh6M1JTluTBe2R+
FGQRfoGNoMU4kT4z1TffstEWoe4BfmI7bEWiRGbeqTmS4XTjdpU8em5XUexY36xzrXKIeOYSz0/l
ryQpOVw1TEusyrcqTjjrMRgisk8nMHkLUdJ1ZkG7hSRzmayErFrWFLSmlv0r0M4MGul2rYzDmDEb
SWqT2c4x2ktsmSMPHCV0SsoOOYJe2XDTol6VmPEDEjZbgNOpfkv2Gb2fLvZ7hq1ps3IOl5rm1LxE
adTvS+VRwb/jg7OeC9GyUs+zKbYuCyBUzpOecnn2pndrDMgt6nwg2PZdkF6BJ+BsktHW4QlOT3v0
L09E6wMflN0RNiNT4qwvWo8bSl7DvZj4G1Pi678Nz9vV6OwdLw6rK9i6fcxNwKLTfi69/7gm2iSn
B/Dk6YpGGQrRWlrBzFiW9QuWrghStirmwQDg9tUcJrpUAJPWuK1QuZsRKD0pFqR6JF3bTQS6Mfyg
F3vlhFwpi5+e5EAYv5DEYe1TI0r604pskI52lWibFSXROtj9sosH67WQqTleb9s1FCFmhEZNmJkn
TMWsH5iqQ9zefvsETQ7F65ScZaO0hEtO7EnRlw7TRl++CN8RzsCJNsoZRW4fsfpIW+3o/m1kdzND
U/BaPrS16uWm+dQn/KolL0WHKHN592yESotmKl/fZkah5LpPmseridougls9/Iwh4UbYL1IOfHfJ
aRztVmvfZi6sv/dA9tSCC2u/OdDh4mN5E8d1PGV1071i4S7VW39SzjxCdIz80NsjmzR39D0AODih
q/PftSrbyRz9+n0vufzKLsDKZPkqiMZ8CfV3nEi/9H+4kCXJW2je438N7+SDg5Db9+UI2CztkEpF
T9nWxIKtZJQqNXBRHRdngkH9go0dNQTdofRF0ZmNk0NXHFfOCZUWSuiyWOnXIDp92GXZmwQAPVaQ
bpGb9UomekwlHkfPl+s0nuXGsmhAG++bR5HX5GbR+meZsOR2kNjKJAbJxtMKvs7vtBs+i+nWkBb7
/k0zEuwxYH6Ve4ruU0xG5YVvaRqoVwJgmNWn8aRsVkXPBhZO4OhplF3QfSjh/YIiat//z0nns9Wn
bIIkXaMQsfxcy51XJZSYTIs2qCDRAFkTEdpEt0Daj4K/9Tz7K0Z87ngv0+RgKD4KEDVpOtt/PehR
nVcMX/EPUEYeLJOn6DZZbsKX5EKifFywLqong02DmlJSdTx+j4xSgL/v1ESQpA3AHJm2LqzRjyHq
yWRi5jD2huI2CxXr0AEzY9f14V5L/QApyj1GB9PdlOTirXxi5Fewv5TDhhDn7RkzWUu8vCyn2BRd
XOIHi408bJiDJQ6+IVIUV5mg5wPkoobnMFHUbVNLYM9DF62D/2V5kWUvth6YoAa0lR79e3Bsrqq4
MeKdRR6hxTX9MR/41o5C/IbOGUVjWFHwjnIpsL1jn9vvnkLl1PS00zV7H3kov2eE1qKNy9pHMFy2
L/BZc5zYKKodISrrvSKVgy2SwzG2p8aeNT5NrWbnbeXOqh1XLy8qO/yzlQkDuM++DunXBUEX7yzN
QHZ6ZIijkSFBCgUsCaE0iQZETPUuHMAIA9cbt+jY7DpHTPdBNttn0JTtLrJ6hBX9IfROFHxUgioO
vrqkJIoI4VL46XyXK5xT5GjV+QjPbY+Mg6w7irdAAJiPzR1Y5LlZiQvDUMlPK9wosDI8oDbKMR+d
Y7b31HQ8wLPYmeXlvmRiUcRMAHfJf6juLqakeP5TUnd90PJhlBJuS5OGkQfp76IDgb2EM5YVylp0
PdTwFwWLkprtjPSG2VfaeL7+BCg+kZcAI0JzI7Rekt0K5jz5gYmswcH0Ubl0WSiEMqqOseSlnF2c
P/7nLI4v855Gw3T81bCn6N/CrZJAG5UyQacAEbuPkdFuh56qOPKImsWhziSScqy9osdXaUgnnUk/
6VN+K545MVR5ThfVOg7EMidcuX6Av5bOjdRHTMkoA9b4Eol906fQ7ls1new3EFrFQeBRLPVrQL05
3kiGYJP5Hsgf5vWESA3/vWb42G+bSw/z7W2mT6L4jLviMdXnV3yozDVdkwE5JCY2txXwhSJbtDwO
y22GeBRWcDU05mbJtCq3f263SveqgU9kDGLfbswTWhJg+EFZLCBQnOUtrjrMcCydbhMH52+dDdew
O8amvFl/Cs4GNign/cfxa3hn7U6nBBJ5wgT1nv+Sqv+cCx+TxSByLTnjnGIWHIclW4U5AC1anHwh
R3Swi3xh6prgCb0G52SUdf5wuDFnTayJNrFGFV8yS9gvIjbko03PuzzNnNkY4TLUWvM4PBT2VM48
c12Xs38KTnl/ZszHLCFd1f6EfvJFD1pqd0DhE06CAz9VDfcGxvXbEHMt4OkgCZbmU3RmWPc0vMz0
/xYAuWavgKpg4mmgk+YLXn/mLDcz9UNAay6cnbqjxDObjmRZHv44DuEQnxh3X3OJa6hpD1KsrVPW
nacdHCXGUybK39DrUiWNUwEIEK4Pob1J6fRozez/QQYXJx1UCaaiuLwD4Vzr/aJBc/HrZl+LOid2
FAPwF8Wqlvd1GLVY/o09ACKQsCqSzpHnHdtryzJSTO/dfyjmP0K82JIhfG4toNi7hI93Ozf08e10
UijIGTOe+TgsYj2/IyoSnxX8sCRULDWGJqP2dejfJtpjEqmFwIWA57Z/6ecclTn2ncnLFVLReDkD
1V9i4OdIyJ8yg/bc76+cp/BreUGZ/zcT/UCszdYsEGKrMq1SdXs+x4ps2R/AovJYt0x3x0/gaHvG
3iz4bTJOWGHO8fHTBxJ2Eu70s7y+s09DM9J72G/zFQ6Nu4l25UwllyszdjuBdUj0uyKsVzCE0Ub3
7yyWN7CwoCimgutVgmsFX7h01MlAHdsG0QtSh+WhTSIwkXXxhZ4AyRS5Lxg+uqIH7ts3EX1SeywX
SPlDXukKsjEgEp7Cnr/dNWdQsKxDtKoT/rniZgCFWec+5+94JDNrwx7vpGh3SdCho4p9qILlv7sJ
74rPXXdktxzPEF3BUlO6zDTobwabpxx1st7VodFeA8jPCEoJjuZFu3ENyDoAKSusIi7garKlvMmA
GxZ4kBZMmS6kQXfEB8/HpilTxTfbrsYCN3K8N7k0C5UddhVyZORd+f3v1Au6Gy7VBDG14P3mzCza
z6veNm6J935A8pAMmnFYfyNsIXnacs6tJYma1y7kdpBSoQ9pKCNr1f77e1aj5td39GNia/2s9kXX
+QqWmUiWMVEOL4e/a1X9ZrJdkAm30lJbkdPhFkmtutLBofIeqXK3mrb/vnRYFMUce+9dIYrMKPbF
RqWjmgMj9mlT1J27cdX8wzra8AGOR45POMO9ACXKXCpwcXaz+uGT3UgdTMu0zCuDYMzso7QXJ6+b
NRvvIBCA/m7jxmoMbD0kjk3pHZcjxpkmVH9ldAoee+O3MmPUXS5I1fa9NfmX2ZMY4829vyiecEhu
SJw1X7jfGfdRRTHHotx+y1gq32/TBQO6f+g1kMOnSJp9DWft4MNUkmWw9M2G4IrZwM3gkkW6ta/m
SIcHV/4nFwq0JmrNbmvfvkXTyB+GD7+blK9xDrIIy3DmY7eZdhNBB4wbDghWzQ1kYSf/la7E0n8o
Eg9qeQ5kwwPkjoS/eEzkZ1/uy4vWiSQ58kZQTiXDlT0qXHankIhDHctGHmZhke7gGi8a0M4hS3My
RmXuyHr0lQhNp2rbSnK4lfcSJ4PS5rS/uR6DW4z6mFz/NWh/ROtwBMYtC+Ob/WNm8yIhmTUiu7+g
PsSk356gIlqEGBn/eTgv66NPejdXMNX49sFudA/mPl6jI41u5M5fk4l9DV+nEKZhOtzPS1gELv6w
mPmXmjtAMsWxhhXp9N0M4i6Wa6qDkT1OBlXVfa5Zki2jQZrOla9Y1HPLUdRA51dKbdzL8z4rAUS5
R3oEzc3ksfFUYiRNtezXvALbtaZDJQ7gTjkNDDsEdpFV3R0F21KJUpiY9bymmZjkb4o0lCsTpqWZ
yVYP2Cw5xqKDMw8uqGLap8tgIzwqhvXV7ch+QlRc52VftrnXLBqLnaQSFcZ95HaWzroCQzO6N+SS
PTvKMmJ/UYQ8X03ETsMXfqbpYNr3/flB78+X98nrfUXHrvjBXHbluM05IoVO8e5kTMa7EuH42Qzt
mDgD6oGNwA14wbQLY9c94tX68cBcuRrXoujr+LqzvTdKwln9nX8o8yRRLIQmaBAELILpileYLPZq
DG5CC9mPjPm+ixYTxIQy9HtleqFIebeE+YMvVi4u6k4g7hI73HlN1D+gQM9FaEnTIwCViFhaI3Cx
5a0U960DuwZA0mIJ+Q6/HcwU6x5AYJfvjgKjeuHvzs5MtIdXwRH9IGRsad5PklfsfIu9lK7wmxQg
PIWHSXB3ICZfi/VLHuFP6hTZZFfefUpyCeB9Bfc1LranOh599jv+imYLhsoqA/e5DTY+xgJVwTgo
cd/j752scgygiCo9yFQfTlztL1sxlwRQeS+C695ZxRAWOJD/iLEXMJLbFbdn7ZZo30XuIdzDZOKA
jv+8w2OdTm1L3U6QmQJvx+dvKEtBS9bUc5MYLNobWHp7kTGvt6s6A1HXyN5siFpnVs7+LanphOz8
zlTqSKdyAxik0Cr/0CvQAC1kyCZ6kyX0bpPpGf1XYOgtKTGNCISGxOnzOQaTG7YVxUL4ekezz/ZC
p9rwUcx15dhXO1gHnDo3SiQA95NLgCIJ7gECDrBj05eGOqi7o/RXukf7oJ4OVdSOAluKMzw0LRdi
a/nguaAdoMrp6b1PfWcjoMrg3xbKsvLy3nQA/A6BSyXxusw1Omaf+nvImqBvmUSBT+bvAeIuBjyb
+U/YKB+kwZ7t9Eew70ZQvRDoKDbLUtOoqoCFcop2QZEOeDLofKehN/RHb0s+O5ku9e57YcqVLOWr
kFOStfNL//ySFh0DK6SVV8pqGPU6jy2hjoO4EFAdYBWY0DgIvWmqHRF5eItDBqF7Tpz36N2ki8q/
wa1zo8De8btUywyY3j0VGjn/G/UY2p3fRKguwLT80eDCra93clrwlei6EA6DIca6NqRvNAJO5wA+
ln2hBCIcqOu+5+cSCUy3nVjIfqK5GKY7UvgiK60qg/BtwDa4OvdFUA7kfkubvAxqf/Y1EE77cQOB
rACf0eivttlRUBwHJt5Jr4/4AvYkZ440XhvnIDcsqOTN2nZMfSW7d8vC1iyYrYTnMae4G6WIueU3
5rwQnJ1ZqQqItWpn8D11NyMPVsI7rVrLq18rVWrLbCTzwbPJgLGSJwSfpSWP4VMvcZ3RN4JH27X7
RDN52SJUzdUOJndIQThZcFfeHyUCCN0bEAY1048FKxYTy2ejghDMYQ8kty5KoAx/sCuWZnzFMknZ
5KUcJ1x7Cdi7i90xPd6kCfrsiQti8X465iopeAYB+5pI/BqeC/fDDXDsnFmHHIVO278fLEtMSLEt
1LnLAn3+hsJ/uzRwwy+u2TZeDQO3E2Jl0CCnEqnKWdPuPnBxxgorOIcPFI2xKLm6UmQYWvgje/l7
LEUYHh85ExtDFGGJn2lJHbtbTINHbArB54/Xg17CLWJWfX81sELP6HkBt4V/P9WjR/Fz/OUpriYe
iwYbZQQKM7fMfts+QbA0fiCdH0sMqJrS5jGcQ84afJGFUy4ra47kYvqb7lZJnHm4Zwsy5AysfoZK
PkAWS7jV02OAAWeE00Rrb0Vr2CMRc5nG7vg5hslvzfkHQA/kqmD7ZftXFPEhLhJjgyRx+htj/uiW
wkIYMIhIHe4L5ahE+hLVZjTG6DhXv1JEG3NkrVh5bF0E/9DURNfqNl9VmMjYA6IdStCrR45VR1tF
1W2lOsYe6Vcrxz/NxmZ+XsC2PnUCYpEd/tvu5jqAAhL5zlZUVdW98Dt3UhGOlqnFV6rCCZJNXcTd
TXEVfFU4d5WS0S0GBJeanIv5k+i++8XNxqPyQIxdbVpKR6ZJKxXQ8CtrEMggnwlm0HukbqC/5Zoy
sYmdglsFvbMMB7cfW0KlEP+4uHlYWptjb6dL4ySWoL4tcD3ktymKfbmhqDl7dzM6VgxoeP+6vcyl
k9ycDvu+CfL7pSoq0TP0KcrpY43I8gk7PZgIREMM14qL3xmEF4ZnSlQ7RphpC6epAGSylFqodpNI
va22pDkYHy+hfW9bdrt8P5ceQKnb76VRg2zh5+I16IhWzqHRUHssYuc1gLtleAnpAQyifnZDQGWe
NOk2CTklaNUCbkpIpJ5+xT31wpsiwiOXC1TuAwhOWONEreoSmObsSvbPpVfUT14OuOxL/U5HDBdB
cUAG3LMOFBrC3TxC/lgb/A6+aVZqnkWdkvnMMIev16Mcru9F3JP9YwxTKagkQZ0gkO+Bsx+r9EJa
iL37VArjWMgaJRmFm0Fl5Jb8f/sOQXeWE97OqlsOn3mxUFng3MUwwAKcQ08fBvw6Xg/RHyX/uF9W
hUTx56j8IXdcDF2/U2O+gQDhuXieeNmcTXTdwAA2eWqMlE8FuPnSZ6riNUH+UYbTtjTig9GXZLSI
llyGSBMBnjnEa/rwjmt0OoTU4b6zLM9vT8EKZlGYFwSyfgsW3SbYWZ2BTRaJqgPhKo6jLfVu5AhB
Xyqni6akzqqt6y/YB7dDYuCuB/mTPVz6H3+87Ho0BsnWZBDUEOcSkXYSoBQeYj9RVC1P8i9FKQVM
yTH3Ivky7FFseNAz1oimdv+daZQnXxz1io449Q7lFP4DV3TTn9DkfF65kVSQZ/8759eUABM+Apg6
TE7TRzK7LAcIhrqVnYu0pNRgt+Y1B6clW8gcQtztrybkfwowX+FweQoj/GwOBXjEapTx7GD+3Wf2
TcurTeLjJkGFE7HlHyHQKQPoAjnYzqgXujq1y/oo6mvK+rREql20PLM2P2OyfMr7oT7lr1wudTzq
TQ88WubQ9s3oRFGnm/SzvCOLzQRVpv84LoBYtKG1LhmtnJ3Eo7IzUaChQ0SeMS/WZNUk8saumur8
sm9mjynHuoAuQF6+2+UQW/ehPNMVnT0iz+umcmmU1Mxrir7U+HQpuXVO1zbhDzZq9jZxRgG9B476
Y63y9/PYaKD1hBUWfcoe9pvhNoBcqKy2RKesvlXaNB6KVaN7g/FaydObcyRkhYmk6aOfkfJ4pWPs
J8NT5TO6D71LifYEAqCUd7oR3NpOK1wSRn59l/aoURUCsH9uoUPWbybNygKSnlPDn+oQAGZV/ib4
pv317Om6W31F9TBr/fHvvwRtCa3GDiY+iYVll1zluVl7vFUEiKL8DVqV1NW8KZ9CSmWefSRPz57n
Ywqim42xz8F8lIAp8d6Z5yjcGCE9mir2UVWk/w3P6cBt1hG6Dem4ooC7pEQkAVhq8qnlks/cCcqF
ULYkX00zLvkM255drgtW5Agl7fNqEz8yEJYXvn5danjwyulrskgK0rUWXwKttXoZG0qkwWCx+koM
LSD2BQ6fDunw6k0wv8FiEA1M40fR/gzCMWNZ2hqB7SY5sixxTJQ+KqMoeBNMz5fHVFRb59TLoksD
sC4psarww7MvJqWH2Qzb4zx1EMbd41gpNYGCjUMxQiCxiUJ/3+kPOkOxWkfJrhL7+MGouIGs7cin
+A8Uw5+XIOZRebpmbcjarQcJe36432zKmBU918XNMfgIkwZxlXwRurNO4J8M2B86CIos7Uy8enoV
oPzIPgwe3yXnTmSXnKZWCMbNhQRHpS1c0uMIHqUInNqW/z7TaesZKk7C8eempjKFz+3ikUgkNus2
vycmBkpLkq05BuyU4i7i3ZX5wsJj+T1czHtM1aJbIVQUuBBzq/1FhNZvIqKrP/aVx9I2+3nRmqef
8oKT2cVnRluTAJV7lxOGr+Xxcc2UmspOaHGEi6VVBSFEcnM5QFcMt1RK0i5KoJnm8lT+sMLszbTX
kDY8CEP4vZZMHkYSlcQMxnk2m0c6n1/Mmxhquig9ToyjkebAoOcxI3tI6d1JZIRbAwWFOD+xOnwM
vtdfcloG9+xdS7ffmpB9o8ajjk+Xc+cuI/Qo44pO5vsNpZIdBlDz8eyYx0VQfQS9bNiP14AizAxZ
DO5FoQnM3XQhjbYnBsvRn7Pieosu/GnYe2bm9jB3qEU2oqlvr169yr5Cvu5lBSsZ8ga6W6lmz1Rm
YIXqxfBqX8hVQtsbw7LLrypcg1kPRZ9/IQOtt3oKJslWzOS8YV3+NL9cAxod8b0q/oYizGX0evi6
O4/4ezT6GKAdAhBEpmD75LLxxlDeTxuetk+Zb0xNihReq6Aq/55vi9uI6Ds9rXeuFt3srPwlulLL
rKSK66U+8q/HibZYOeM5d5RPDZ0pt+TCmuyjVvEyfLwz4i8Vc9GKjSNQ6crvZidhTe/QD1oyu5Ks
iFDgrqQgNcrsLtVXDsy40b7rcdg7LJW9CCRCSitvLUAhxZPc8GhG237kQR29frjE4DzAPiV59fUA
WxjBOa9LqLZ1QM73f1YJP/XRrGdner6zrCFmnZHdf7wzAshNiGrMKPSYAkPaj08P5HJzYKIE9SHP
d9sOAju+PEA7NwFXMDD8TVHm5wgSq4+jtHyQ8lET4PybzxJ5jw6UnayHwkIM1i0ZEJMDlDfGIZNQ
SuPtzyqT5tinNFWENRH36YxvTYFv2Mdg25TO7Gncx/IA+guo2il5pRfgZlKkjmHp9QFEOGlEUI/O
QARF4PgJZ7P471i585NOnI4blbfmLDHZTkETJuq9QkihhBD620yTBGmrnsBDyLS/BTDfES4bkTJ2
vpoN5j/+geGswcyJ00WNEN0sPPOsFEuYhLBZHMOdX9ieNnwgC0s/2YmQxgM94t0qzlhWkfOclK0T
4N2rZTlxTqfPVyYpdEOlg4pH2JxcS0zTzig3xMfWPqvsf9X3HSns1EG4wPswlTPAsgANqPwzMm9a
KddPEeggnxwRBo4sI/cdItb5oE+XXEezd+MWI37rP+MlGpqn2+36sMWQ9og0xN0EFo2/GtDRUkPK
Ur2xAD1VqHL16NoRH+hHctNPNpVmpabe12FaSXZitVlEw7zn43EfeyNIFdoEtnKLzfi6NScZFibX
/HLbRiU9LxAwUQZuw+Ujz3yAzOGUEjxQprr9pV+ZnJwJkI2E9ImYXiBdWNK9Js3nLXwfNN1YDdtb
On8TQYymCHx0yrNQsyA0RH6agAchTYFfZ6D6vFI5T4C5po0GtrNGKDFcClLQ8QPo5l2qk13Ui7aD
hstLzy8FtLA1rJFfulL2Qzj5zx+QOHJTl1m3Dw5V1UU8iqVngZEXvkR25briQE2yNA494XOnDXtB
lQatODSm9twGzYCaJyizsfX46EofNoEs66QJ3gDcmIA+WQi4Rv+C5tYrMgN0yoyaGvQmn1/FBKnb
D7+FJW+4MCv4AenuqXQl1rSSXJuQU8NQ4s2pUzeCxxhBCK98K8tkJ4XiBWL8YlImg5uAeva+jMcq
LKkc+EcGf1gyg8BlO/Sh0HZiogmy+VT3Vkp6rLNDkdAt8iIzjggkWfdvTMAoV7lp1awrHiCW0p8z
ICGqzb/xS0SZpMqhNTAh7JIYByfsnRbivzOGiYXi5ODrJ/W179KIiV/wYYUjX9+M2M7JNnGfWTGg
uN/x0cFbwu2yyYA84ZGEWDD0p3MvHwzeRRtHlM0c8MnCtLXgQ0rPXyXghTZ1tL/+RStCTNYAUbV3
ons4Epi82dfF8JgNTSWctJ4xARZSuQpsGKF5oF2Mluu0/OJQHMj5++u1VmJAJPm7o3uJz9uHyqjG
Usvp+eM1EP93qYSFMAk5HEGTUPSKnf+luIkWVunYMIuVW11fHeif4ov2YF6BcQs18T4e5HKX1rG1
Y715JxAR1lQyrVcSBaWlFHP54Eb9+/a4wTYsoKZsym4EpIKqFsPl2SPRGDBg9ELHOn+das4+thWt
bZBCENCeCwXeUsAXCQme6zplehOQY+qQx3/qn3wLc6E4DTVkr5eUQYugrKVy654vP/eB7Zdxw/DE
gSYNBOWYooN8SMiMZoW35Ad808yBiDgPrJao8WUzLsETBcSTmq1qsPlVNtfjbx9V4isXCxXKBhbS
j201m+P/EFDGsb0hc5LUmjJQrnU5HPBazMKgwAxvGBm67HWPXK5irY8sSXUfiEzL46LWPHuBCGK1
NY8ubKK2+R9Xyla5Prz6iykX6UY5V7+UxNA+PPa0bPsB+3kruJy8xSt1df0P6qWepeUtwM87hQtZ
1C3x+yIAj5pDcnnbuzUbOwgxP5C0wSuLK2DLXkHnGIuqEvAbDV4FP2vrMW8gec2fnwXP+EZ/uoLy
a0KEXKrXsMI34KDF1u7SJGe0L1ZOflyebc2ax8YJrdHkcW3oQWrLC5RFaOa2MYU4NovFzqkxdhuP
MQ8JZVBp6PiFLhuxxV9seJqh5X6bMhaVpmX1yJ9YM36msIVMQ9n6RWTCc2ZZ6A7c3qTgr4ap4Jlw
1AEbv+0yPi1Io+ljjsujo/38ALqih1xNfxfvQ0D5SHQyCjvXmIslFWGdc7z5JS8oxJ+UIMIXP/7b
R9jHqN5aYJNJEcleCKzNX3xCRyKQEyQiPMYIgi9GFCVf0Zbi9EhwCcThDgArYhcqv1qVlkn/i9Bq
2gR3VDXQ7fxQbjd89xj1KAxfOkMPqueFG6hLp7ovSwgnpiOm9X7MZdSn1x13Tg3+EbOE+wkDx8El
WgYUvGED0DAXlkV4CE+CokHfNsjI8lIDvSF5/eHxk6gG2fzEBFQmTElVsuLVEbTFOo4d+LEE7m3f
TGRGwDwvxZIWUSC9mHfBjw8SfDgxhu6Wbvv5IGpKagrldrF999vy6RxPj0eT3tF9umGAu4sAwaag
//7jmdW5efIK0hA38yasjbOv/ONxe6uLwSlqMsuhAf55H1nOafcOrXy7/+QG4vJO2SMNkVvdYV/W
ILPq5FPV3FKtcTStoAol9o1X8pZWWXBrecVKlRwW+mOn9WTlq4JwEx7mqADYRgyVKAINzV0eHu/n
R3obV3ztTPLLMFDBwYXQaAOysggEDsM+No0xUcVmElZ0+9c23U3gDfn/dmGmZVTVQAW3PrjhtyDt
MByfgBjxZqFRlQRuDMECxEXvLyeT2JmgyPl90Cz4yZZ53EJK3FEb4Q9SA1Byk9cp4OwUlTnYvEdG
Zv9cRL57UWuGvEFlruOqz1c+TFE8W4nC7bg0vHflGBNvKQ3K7JkpKkPgrAvs/Ve0+IngsWsfo2sp
OZNdqGcc5jQM2qaaXPkWO5B2AsmGs4g3SqxUMwIBFHDKcmBND1anRM0SV6uzbc5+ZDWoOix1eA14
dpdxvwrMOmn4fZhymIphiec2d0yUn1pyATFCrUZYwo1VyQHpNiIiD5eWZs6h9kmn97XdB7g8WjsP
xGJ7cgzPxy7MotPk4ui4O2DvDWkdNXqsRdfcZ8WnklUPkKuATW3NEyIX0/bSd6fN7rpGfK7/Fkaq
7jRMVFzGQuS75/9nwaVZQbFTsAnN4CYmek9ypCIDpaVi87QRJixnnr7XyxAcJfaFdx9vVWgCPpCi
Hd9Qrax3cFJeLVb0IFqYcWJ1mXk96xXtDdwqI6fbSbP83g6ISXwksyPd3WK8LTUnreL7nbQWIih7
hFjs69nlmlgKiFkbWVcHeA5kfMWvY/TAjPqL0QVwBsYa82Nt9h2lNfOx4S1MEmQiuMYDWa3N6LOo
gvHdLBjVi3DrxgD7VXIIktz8mK0TQYSHPph4ko/UxVniO0k42JOfMC3llUwnbWkWU9EWUcZ0tNfe
U7slCWLrC+IWmCdwT7OHwYh50xoBaD9Q4yPw3vIFBMZi/Cm4ecC4yRgrzqQP2NaDryJnA/9P4S2w
Fbf95ahbAwF+Ln1qj/jSi0YKhQPjWHw/0JYieSlo0O+ZVlNu7TO4tgH4aurgo5LNoPTo5l+SeIvM
e8eu1W+G3xQ5i3hTbuYLgcwj8PaueZzySNZTELvtM3e1l0rju/vPUcIxYjm/Alvew7umfpe348qp
GA3wxmnnIxGjLxatw1b1xB9aH/sn5/O1sjrVwFtRY6cTL/kLggFUfebHQEkifCG7SS6zdzafxnxB
z83N3wlcuywEp+d5hYqk71dQxc4YEvGoHKJb2bsbUiT02Xrv2ZhxQ81iWl59wiERPG16K+Ewt1kV
gQA8/lYo9nctDs2HG9af4jN5vyyIIIfD73WAV+hyWrDvrl2g2Kg0eWN4HJ331nIhVuBvUpcHano7
BmiqEseQQts4/6SraFufvlycc7xXxUvIqTOe/eiAijQBclgokxKxwtKZt06QNTFkJDP9hehaholr
yOAdmTgEV8z2fsnsXDwC1TC6EKAAfgs1j/MRlWD3JlieGaQV0bZxSBAEg9jb6LbBWdwP+YYaj1ZT
5i/oKYYorhirBnzbkStQ3nHNs9uR+p6MyHxITtPlFIhS3urIgmm1Ji38AW+Zguv3yvu3gMXzBAFA
vHZzffHHquGVjz20PlevRvEmwYbglnNLx9YL5iktSzE8/0iyMoNOupvcrEs2j5O+frL5qC/5rn6E
g1/zelLI7HR8y//kycS4EgtztPKpWamupqJC/u7SN0aNzfDzsk6GOxACGnjjvj3BJAjmEGPJlHSF
Dbf4bwSC4Yn3/byjHsEiRFqglMgMCRZFdR1K5UuUSdEgg7GRwFMTyRJD0Un0cRe/vUpVH7E/33Vi
MVwzV95ihTg0XHWcddjPLrtWNP0TeK5e4M2IyGiy7FZr22abwi7FpnjlC7ydQk6nwx0oki/WE5sZ
l9MYkoXgQS+feHOUXK63ZmX/1tozhf0pfe+BJPeqnG9qqnUtm9LhzYH7i7BMPdPr7CI2NLM358Ym
Mhd1oDJjNRcwhBq8O6s+L+A8gEZFdsW2+WnZ6H5Hu1YYi1MAcEb10hhkgMs3+WpXDDxAugebNN95
AaIS26N5YMBaGkBvFEkiYU7PPYllI58aMuHbbYBCIAf7m95q1t7yvdaytOto+LdqzbzTOHR9FeI6
fZPNgdGndLGrLnw7WlqQTfjyWVUtZkzWtDjmy2jO4j5Nvj2c6gIbR4qEChJ/zXzKvRzIU0vVso5n
nVz4VWqescivh8O667YUw4geK4mGynht5yQhu9RB/Iw4BfPe8WVKtea+sCPUzZkpXjb09wfpqBYB
BFrVIAxt0ix4u5oRApXvR2c51A0oqNsF482+PhFvl7mPxw4tUYWsYnT0BYZeZvvsDHrzsb+Jws5v
w5AejNtgx+ageawjk4s2LAroJBNd5Q3FN0bOeqss3g3CdHPq2c14KwAkJF5CJ+ymgGrKE/dlgfFW
E8wbVJrHiBh+T57flMlcnqsKY6tt6liYBLKmtp4seGPC0DlZNdBYhTU+herTW98sXlmY+Qhz/LPW
Cqd/anxr8+ZvsZ0xPcApA5JJrJjYdHOpPL57QoisQuUW8zMptV3la7PXJtLFAQTaSmU1waDbzY2O
OwH1eUYVb132anRhUrnHG8Pl+tVYLSHsNYeVDVMGmQjw//7MqvhEjg4Rg3h0HUegR2NolB2PPvDO
5CMkFTweRlpEUMSOy7NIoWcS7Z6CoSy5HYQTd1xOoSGqUU1I/TMyIjmUj4hqxWGF5Wel957tBL6Z
9eX8PFL2XpdR2nk1IoYcagy8BjkR4P8Dslgi9JXi8oGiuXX5exHGQJDCXi8Tu6fjiZ5KSLWq1kGc
NgLWXW54YgmD4jKfdNBubga8LN3AlEuQBDiZ4woaqm3eOJ9XXC/6OrUzXYcM+DF4e3VbXDCQEv6/
HlQwUhyA59kChBoNsml54zX5yhyJ1cZ3Iu8EWpPGYp3gvEaG8coeQ9z8cKjmIU4quvqF4kqu/7qt
FUCZu9XiV4zLRkYjiCijMCBESJ+82kfeJno84aIeFqnLgnM+SbGkcfPJ3Wis/byd/PHsLAOSQhIb
DVHIDaZNTOwpIT8N/j5ovOYrI/hcCUh4c4qgJBhAwtjGTJlbAHbgOtjH/EWaqOjB5Dm5H+fBj+qK
Vk/iLZRGs6EPeUvkc4ifN3Xj5jbZ+X7BxDcNj1qdF16Ztlfu4IgjHPAZRrO5STpHYN9fIWTZi5HY
MnnffdfUNgikxYI61IM9/5qfDOq1skDhWgk6v4OWFxPsnCVPgLPrNrQuQP624da9gvurftvHW70g
j4xi6vSeVPDgmprnwsSldEl/wcGvPsIh3jo2a11KiErAxt6jxw4m9PFfJIbIyh23GkQpYZap+qfj
wW4j8ijA9zbG4IzFmfnYD++OVpIZ5x6BqjWT5mRjQYT0yAuMqlKEQhzLf38GRmisYrWYIlSX8K5o
MZfEpALKIq0u/y30VJn3wPSUvU0SZZAK3YWbL+ed9Om/i5Xd/dsATHQXjgdhyO3BchnhMy3PN51L
CS9tBEEnn3x1e04vJKoYqr54PaEMJahMriuSrmtXqtn1OY03IzDpwnYLaJHEoDRcNpoZC4JE4s9U
ICbx6tk06lNMSxLCuJzCxxmPvtVXY4a/L4g8n6evBujTvvHq7l8XzHGVJjqy3ggnDkiE4ibJdQvC
94bRVExaV6spYK+n5C5tf3fpj5gDmcK3QMvAEtyvsDfAcQRH8y6JJ6U8Kpqecqi3EhbBY7mypbcw
eQaRI89pRt9OdGqmGr/UlsDQu+FunGBmlUrMdavfJ3D0eJ5jC9CJt/ZN+y9r9D0LScn1iK3dOySQ
pA1gHyixnksapwHELpOWaBf6YqvPclYvN6xPZJJdnRkzvJR9L/3jsp3LwUWhYu5krbNoRZthYT+Y
Vp+6ltnlI2ugbnWDodk7O5Fxd824HHT/L7Kpd6aS94ZR7WkWKfRcDgpR/XxP+b5tfKIfdVpPw5m8
5cClukBG63A7c/K3jCDnCErITDEmLpTuEqdtbcHmqTlL81tReJ9v7BOEI/FvAJIy44yGNQ4aV/O6
x8im4r8lUmsZa5UAYFOuVpaYAbC1dh8BByvw8nuJP+ycmiOifIP2CH4przi2u4JawLFU0nm0MWYn
KGFYC0COLvP0pDGgg6b0JdI8Jwja6NlYN6v04/v4gK125T7Ie0Wq9eDOg2eXQ197/xs1JWBWH7Ze
Zb9AyuykmMqo5Alg1WWWmwHpuwPl/1Sj/LaP6292N/mZKXlaqe6hRjoRNCLbUQDf8ri9/m/0Y5OZ
ehuxB2frbJcGAqRO+Y8sHv+Lr3bbxEEbcN1nK7jMvc477HwxlJjsLyhwA1NNptNerw+1+6dA/HIc
SQ2nTp9OHjc9XwtDPWiyFIShcLrbeJwwZYe48sHjYGpNo6hG+bkn684F3fO5tresBY5wVRI2sJqQ
Sb/4JIXHGM/4X0iPt7/Jgs9jW31a/X0+EPRJ/V7B6bSpGybyw8wovgY8Mpc+n4bxFjoMafA1P6dc
VqeMQfx59NsCMepm8D8SY8R+w6gdTYjiVWeacK7XqE9t1q3mgGy07BdHfTlXjh+8YB0d3IRLev+N
QxxesgJEtAGUvRY84oYuN+yTnjiMOU39IIYibMIXdzBLy144XLznn7qNLhMTJg7g5kZBdMeNwpIy
hXY2x2v7gC0dLOSVbIu7ewFP9KEubmtlIQJV8DL7FUqnPmN1itZjWkeCiyuVUXsvuapgyCbYaq7I
KzIaCTXnTbgEPF3bDQQgtjloYmvjugH7/rRonrd/SU5Mq4WPHyZpFshraPI0/dzaihmkj/a1PfEj
djyspMIjQAQuJnNed6ny1fiZmPo0lO4sGbsTqUsW0Xg5Ezxyv7NqWt+tvhw4Z4lcNpCYDcbKhhHN
i+uK6RMrKFbVyn41KoKSjF6V5ksj4V30IK6YzLG33ag+S9jepYueTrNX7KZinDZioO/y/t5k03jA
J8qw+5fnsyXXBQfcKNkEEv07vMpNJ9ndMxHvrrePQxlnp6yegBGeYE+t7aOaxaOhc1T6/8Upz4u1
baPFA/eoEuIfDc5FPizUq8vlyGb9wk7s+T+yyYTVowmFzvF2F+YaQ+mqIM0cN2zwE+tnuIVapGdL
yy+avGIzIwWvqp6AtTAooTrbVwz3hKvqp5LdlQxT+saKeufPFvLVvqzoboLJTrBZHc+F9DOnlzYi
Xl2dctalyZy+dAoMlI/asY4UxbvyqjCjVPXXJ9wd3ui7exd1FhGPRsakfoiEZfFwxBWSEGN3huPM
RaUFXf+p+NYgf3imr2UK6CzOig758H9/0yZjIvPhb2XrtR5kzokDrXnZsWyL+RZZlSh3ArhysyaH
4EFjaXvQa8lDyWwLSqLVBP/AkFoAK6XslnHnfVbTh0nRoqDlYYa8G3Kt/lgH3ZpKRi1sB/KzYZUg
CDkRh1KSCC398T1ocgZFn6rP0VijyT+tCspIp6konzOPAiacPmN4OHc3CqYJhfyiOwZfIBGzu7uH
SwPoWq3hGDuYAAHcU4TwkmZjbvkp9ZZW7rTlTIiYrc/dUK9qHlAbjMrwOTtHm8jCO2ltHrNZlHnq
Hdfo33vBUjztwj+xne+gSQQ2ipyvqxFFUPC8iIJAW2cMLnaNCaAKFKLRKvMReYRzZ1Z9YURdGHq6
mhjetAzJMLN51NurLfu6PqYUuipzbCxGdpRrsRLghdg3NJkOD66hGObSfvBY+x+B7+fIFf2JtTsM
210hqp+Wfc82am6sSvbcyOx1F1eCjLYZvIOiggVbAxrUst6LY5nKZky8IC8PL7JZobT+HlxTtWJS
0YV3xetJ/mi/2ECo/H7MK/clwqCMVguPE0MgXBfHWSiwPVP+feSnV2WYX1zhAJpa8Fsy7iQM04I8
sV/M3I7MJP+wqt+SFnZDRLjSiaEQL34L6jMozxA8Y52nKqdPGzuaHR/4r0Odlwe+eRLSvQLQfDG+
AYoGMVAugQYudfM30s5BPOotTn3XXJcye4TY5B/O0jdT4L8OMqIMrlz++9jppSLuuij+O/tOIFg3
oaamtAOhLbNfWDy+M+y8fYYObqqJtGCnPRI+gyOv9KIGMe4eslxRD/Bl+835fhF3aBqhmse/0PB1
LATjZ1dXMYgpnxuWUDo2hgN5HK7HoWUGAQ7eadrH7XMvjcOrQhAGCpqQQwbn4uGkt08PrZgaNfQ6
l4tiC4zwmSoDccEpvH0scnGa9iiywN9kiABuGjh6fYIVXCJSrb1MQF0F6OqQtEBqPQopEMrVDvrV
snY8GUngK4emkuibP4vS0SOR7V7tIvXMbUrBBk07JVpG+ncaTU42cBihP1hhEU+W73tgUaKvhZPD
f3M6b0JMtUlAMfnjptyc7EUdg+oFZkAjEyxzT2XekNBlaikhiOB2hYPkafczWqF6WZL+nyGNOp4r
j1h2sXIxj4Qn6rANl4vzi3Wrl3LKh4qHymE1ZqvaWHBSFs2CtfpTe2pfisJb1FdCihsp8KxaS9uK
bspFshCX2UiaDAA16bd3FV7u3mvaV37hTu5Y/hLuOKeYPj/sjiE/4t6e8WpPzgc6IAoP/lnRH3TC
l0cr3/zFMErI2r+jipprN/ZVTy+FH/9oFoVvZL71ZlNpR4yEcA46odgJv+9n59MnyIk7Bj09/apj
ZjrgUAKcwzM+/S1BtOJTavQiZVN+y/j80M7o0p0cxtwKba2jxzqnemZYoG1st6mjVDQyZG5euH+7
lexrXBdSMAN1LylcjvEp+cSxXO5Bsc2DwaHyi+TtwRLlWL6wvi3bB6Wab/yklbjJavLo+7eZeiAg
xl7fET84AiLWXs7RMg/JRKfBHP85hKTvYmw+0/eMKYtxRjttPGmKHzoBOkKiKqG9EBRciB7iPtuZ
+bj8vAtENCi7NZvarEquG7FQcVqxmDi9IAOas64MVG/SLfNwmYPmKVjbgFrTcyY407+vf2rg/W37
uf5cZaXIZsC2N6BdjqQrvOfy9zkib61z2rDqjRnh2BK1ffsOYzNWmJIw45XJBqzKavMa5vEP9Loe
bCQqTpEtxSG7KVRyGRSCSZgDmkavZ4FpMb964G08B/lcSCxLn9Rvctlq0F9jkTjD43UF03suOY9N
LRiwWjBvH0cq7HpVO9OgIcGTHyfybTgq+Je79QMJ6MG14Y2gkzHJWjjC2QzIndgmNzxRB4J2oo2T
dqkLtnGbw2wCWXziSns6RDwtKuiFpayT1j4hZ1ggjFg4a7t2u80KWBnE55n3IIpiJSdfWBB23BqE
tmsgzJTVsSYztKHkvA9OpImHXwUrROFhasE3ChM1h5fsNMXKai4XkGC3kCOR2/LYhoUiQvrrO+BW
VPjErUFZYKLndfP0F3x9KfkAQqfN8n0QAcGepctE5bUbFuicpShUWroQK4AeMLj4DhY0dPLruUsq
k+czDK+K9gvDNfSbIwAVZ1QkDVH4vk0fl1TUmOC0jiz5fMd8OOQaf3jfP7Ptd/LcEBJjv3uotUj8
DgVqZLWHAg5xQvzcxaPeBU3dmsbCIVKPV5fRRYrWoaKtJ3XVnHJdz30nODDm1wY2cnoIzI8JXZ/+
ADqYfVEsdhl5q3S8wbDjB7R3auTlDUjFB0Q4jg5AykTZtyyk27311eCnusnGkWA1sc+JJV5lZWdl
6GYMPXs+WGQOldwfuHN7W7tF4ARiVXXVsr8kc28gHRGBnsWuFhgAazh1aMFBRgrfw1F1ujVYnQ82
9lKceAon5IL0Y0kyGHeRVX0HvV3Qo5TTqz3xwoTWy1LvGiVLafN6bCSgVuOOupEdOB6RPG+pikn1
y1NxQWmXYWXUsp+iL5tLczPXaaOePmGK5kGHIX/mkOPSYOBQeKe0hzjE8oW/ObI2BHMWphjMQZFh
plZ4t9Oobd1tbtXWNuHZw4I6blMQ875vqaktDG7smuDcBOkFtBJDDvYaLEAnV2enVuPBP1XB/z20
H7i1K4s26Sreeslfcjf0sX4wOwMIJtoKEosCivlKBL8la2SuhbnKy6Lnu4675f38qY5lxrqiylEc
7pFJozS20YSPtYHnGKdzxa0OVDAvdc50zqakDuTfXLpXKw07dygYnfZDiEsVFPDAd6g6GCsMRxlm
eCv25txHynyik4VCsFHwdnLwh2iuk+icBpCltWFAzUnbvR2erfGe63pO3RgBxSnS38MWKRjnsFUC
J/JxjyHAU/NvTN2GyosqA3kCZc2gocDXER13/PWQZSdcB5ilIBlBHZdH2/rAqIMkh1Nivtf4Ox9M
nkUdP8L2UFW7n/+OLMQGR0BXzvyTXVa6xwweHGhigYKHqLTmXVXDhI2DDtxxmwel1zv2WL2OoApZ
H6jC9gLgJqCs7rU04/xD/r8J14mhKqIK6d/n10EU/ZJMzwLtwsLapfZPMbjxy4VuBB9GDDVY8/FO
z91enmRlKRZYuAyU632LXUWRlMxCA/SxEds/UTOZ7LQck8iUdA0DvMBHlBHU7uqyLoS28RuebZZE
URbf0IiGFz7RYSv/yY5WpxJHgFCcamNJXo0YFXH/hLNCLcHKJkGwdEXn045svOO9TmrmBjahzagW
vmC7h5fl/anO1qokvmWO8EeBrUBRf0eUAab7/Qd+B9F0krEQIU5XK/egvUZIGA0enex2aXnaoaSu
YdL+VOkZ/DWFuJxcQ5brMwfF/TeXRMcsGnCu2KnL45TeNvVlEtzSPHgTD5ACIpw/c+ubyzqDbb74
FahWJLzc6DSP7YYH7mJ4qt1C1ncBLOU5SmytGRhqqU6M48vyhJJGR+Y5WytoOoEFOgwjv+DsX4ai
UhZRyhmIKSHY10TXv2cm0OqDcEjfh14jXlebKLorvzJt2+bYm6rsu0ab3Eoyqo1T2MDBR2O3uyR3
2WdasQ8Emj3QSrpYE8z9VmT1Nfy2T8BAbXRAWN/z4w6CA3IhrIBt9ZWal77Wql7AuEu0gG+/YXo7
CKQbnKezzktqTKPM0Xh0Vs31wU0GsOcT+4BzcVNyxqzGEcUbAWQMTN05LhTppFOLb5u1gsnoq74n
YMkkxxKAnz126PTarFFUKyfWwQGJ3HgmQ9SBuRRx3AuffZpxHQ3Be0MNIoIXWA6g5uKulM4ccxO5
gNWTJ0+3uIqaiB4vYte+vjc1If8vHAncfxM+neeptS5MfdHDnUx29ZgV+eyiW3REwNmDho+qGp7S
h9PEmlMfb4KDxQHvpNquyM2AKV5AoBV684ahubjnBNDrfU3Od/kBvz7X4fRp6QjQdTvV0ATG/xpv
Jx8z06XL2GUW+e81TdDR0zZYDTvVqrY7nlasoz4dByZdFMj2yY6UeYDS694YRtveSWdxSNl95BUe
aK7fu6IFa0xInORYOAWOxpeojXyAqQREWfiQrKMWU7GRtyqnuq/9Ae64bWE9QHYxQ6h7xOjefIee
AtmVNemm+CbyFjpjgmYJF9tNivyth11gOTZpx6oxiXUg91nWKTwgMHV40NcNO2IuhgZbL2+dgIYY
XWTb6J2y+5Qlc7JZ3M28nutluo/aBC0xa1GMRW8o8EhIPsBVVdEWFtMUWG7LvDk8sFmxDoO3/fN4
YG1VfeRPlR35MqXLsXI1f4+rw2gbDEEtM44Lpfrxq2XiDiTTJUPP683JlWaAcQflwHDODrMTpTI2
oGeBrnd2ViGekMvXJB1wf7Mu0XTdvXSa6Z30/JT4p9iukDIzQaWheceBhcRp0NialkKcORe0yRze
NnfTXil+t7UPfXKdfoMZu1I+Sfu6vn7VUyAgmuy5LRgS9KxabzDDexw3XfCkurZCMTTZjXOZ4EGJ
E3OaAVOvqgJfk+NNvTWetvujfT1/WAG8rI4iuSOA2nxTY1poqiYz/QY1wGmlc9s+1hL7937cPDNC
/B4F9CNTn0d8DKutpGqdOTvYjMKVDrv6oP5zq4Y9ANXS0VZs3opNzvf18Ydyy+IiSm/flhNCbgVz
2a1YqDm3A+tECCkB4DLEHY4fBQPg9xjBomj3cDKNInzr30vxGK34ZFk0TNKc86yfVMOewJUuNe+D
tH8nINFlHL4+KGg2BAWrR4uu/XiiZjPzhnCvXNje1t8U34MG7U2sZsRtXGgdsxUTKG2iX0lbV8bD
FgFXfy2wKtoRd5G7RTT5+R83Sb+ppxBWVv2PJGcRp0RcyTBATDCsk4crN7PW7yQsmEAOjV7BcIiN
YOeuTJChLFIKuJOO7Bx2mXlytd2ORf5oJfd8ZwKdc1o93BkWBGHDssj6WEEgyzsSrhbS/v/Qtwds
mH3bZ1AXe5wiu6CZMdsKU43rUFAYymTyVYNbxv1E22ARprv2FkuT2SA/+smCxE68MZEBVqfO7pOL
CK6WyYc2SyOC0Mgz0mflbLG/+YVCCAZHyHJMS1plAKlTz+C2uSAocPBnHQh71aHQMVHNjFbtkHBD
TT0eh2XKAUx93qqFTqZwLiNJ+Rf1PDD16fDNDngsMfV7Dh1wJVvLL3Vt8LmvE546X44kJ0A/dhwN
HJIMeFDiqIs+6r9jYel4uJUjjscuQ+ARZtmYo0dTuMzLlwELiYQtzg8iH+seFTpqy5Daon8GuPB8
IggJ1Nmn1TvZxgKuixIPZG6Cb8bufEgAOpbdqcv1ih3GbGFV7jAoIQvhyk2yZ0eSPO1NVH6ctIsO
SCHs3kqAlG4nrEOD742UuiYiGF2Hi13qrOxdV7RqQH/+2H9oim+zHAchlXSdNThVHwJw2sisbSXl
drNy1h+qe/MLpMU2avGS1cpFt0Ynda+5QcaCwkMClIGs6zvqDUVy7UkjX9HFnPlv7fkl8hbt/8rR
1qr5/HDctRdvsbwH3i5cx2qpt9M45SnZfeyDZnZFfyC2d+cFqOfqHuCC5AvxPpCvhklTryepqGp6
/fQbtSr+bz/I6aF9E2ic0o4wUDhqaD9Oxm2AK6NKiDwtU06uuDKuAV/ZMlOE8gRTAHWrKX6kVn3Z
usK2f8M1IL/WqBomDW1FY9MRNINXSnKrhid95h7JAv/nCg+Wtf82jK0+aU7uXFzgBRSgg4FSOx9p
Da/Rs+szl5aU1vCcB40E5q8epo4yowKpK83E6t+KGtr2tU6D8YyblnxW0N41q09tzmx6JYyTw38Z
tYn1MG1eHuRekP7FHFuf9nu2be6yYkur5ZGUL59AfWkerofGIKUjMVj1+ngoOWAnx9zGZmakno0V
RIOmgKRTcnCqvHI8ZS8Zw8nV+aaQP/rozkkniwE8YiSYxXaf1g/ppOwnm6QyZH5lq9yoB3XFq9TM
MjOVvp6UeMPsFfoALNpuqTKfk9xYW1MO6/Bj9I90BZac/2ClOnySC3laPYzALXFGZggWAPtRx5bx
xTZk01tLbxJJU9vdpzuYTEh82Zazs8cs4s5w6uwQQat4xlAtrIezolIpiDCydH/sLsoOWDg62/6e
y9ZTzAYKZZ5knIgDg8P7T/7WCzQTez3sWerN72owbjZNW/9LXvpw6xbsD3xpkVYsKybtK7C5FTx1
Bg1IGeKV2+Z3y3Knk/a8rLSj2n81UHS7mqNnbDyYT8mRuFrN3P05h6T4PZWuuttwks4sCPACRy4/
aNOAdAa6uFHPZMllHz2L81f1fH/dXcSNLNZHx4jKCJHXHadTlIUw+cVZIyQu24SbUgtp/M7GmQK6
9m8aMnrnpfAe/1JRjFu3VZUsBrobvT+57j1vzclVtx3gkHquG7/lH16ybfSLT4Ax3/3epgYNTAvx
98cvDjKaR4I//QrHg80js4UCjLHTHduvE0XXtt4iuD2/YjtugnaV1IwFL1OHVjArRVlaWRxg7xHW
/FM/Qbob+INElmsbOqn0EOUE9uO5mUT2o9eXZ6g6z/dcsHFMI1tJXVfDpiodwYWHhyIg+XBmHFR7
cQ2XM4NGEZpFJGTYrUJB9unILN7/ODDgSzsSZuDQv+OqVm1mgvb0+zTdE7JiSy3QOstRko/7nBfP
WO5MtXV6Ngaodw5uvcrTXDsC1s8fnL3Jafs3wFAS1U4qr6u8N/J0RVQBEi7HcKbQxo/vC95OLqUb
alxm114DSN02zeJczFnNLRnAcLN/XpcKV1bhAohQ6Y8r23KanFbOefFvO3PXikvYjNAz6uQCRm+b
eUDG7pzpqcPhwa8jBPmfbkS9jTBzsr5Miny6Oi2vjKwVn05Z/rdQvQDCmKsAImKF7BS7om5Qwv15
ILWIhwmTv6Wan4vceImohLGW6CDrMEqkaCsYdXaNrpscHur8kLpg5lL4FGGgrotukvnkEJKJ6/Oq
hCXRIwuKUJB1QDhnAsaIOQPst+jDbdobczQUjsxUXlbJ9RckjkXEPwvDw6au2ZMQhib4NJdvuJ6f
mr8wgrRHpOT934lWaf8jCewHet4zvXyjnLTHj3t5NoPTITkvkMqLFjAb9QyH9bOFnpUa96jEYRry
dKQhD+p1vTmmuKHuujim626IU9ddjDhfwDZPf4/kC6+PzR21G8I1FI/aHns6OzR5X55AQeDEIojh
dA9+VEJKviaUqr5KoSa44EhX7hwnP8YgeR18dwJ2TEH6+ewJq/0q+kTDc8tjWX5bP0CGTDOoam5K
VoMNjf9TbQ5yli/zN9tBAZQMvjyMmgIY9XWfHffgAXi1BVbXnOGllpOFegYl+hNtSTjetC3MPZnE
O3XG0VpnQfsbzkcF19k3kzFQFUaDNyREL5xG77SVsA3GAhcw6Kd1bx+Pq2ylHONCk2i2POa6jAQe
uCDK531Y5RQXMiDdpzzIK0/WiaTqFp0AAHUu1+0x+IjON03B3HA0f2pVGxP+PxF5SqEqwc05r29h
bMMhJCzCTddrMjq1PXemtYq0h+oGXMKJVkEee+nShFbcjHaiPEpFiYwUt9ym6UUuAgtWTtmeGEHk
aZoSKdvH77rccH4Majm5mmLS46qxUYsh0fOSF8H/d/Lew4Xo8mU/TYGmRKnN4X+A2bvhxrjmPhSz
B0RNX/JORMwjMgXfpDiHtmSKI88p0ha5tsY6klkqQWBwa4YC6p5mLW+Nr4flPfpz/R1qd/wO9qqU
roqgmhrzVVHs12oJMKGe2v9HU2KtvqHk5RrNWgr8/uksqsASkiETPphJ3Jyf+Nzix1ND5lxOQNfw
QfsqMovGGc+WAY0G8xEt8LIvAf9pgOkFPvSIQfBGqML+U13ER1Rc4KvP+A0/Dz27sm6egPaKw3QX
qHfMY+hpkYbAhgzFluq9+SCWKTe39/w4GpkQ7V6XujVm0G3odXoJvYHoOaAYIpapO64xlzNz89DI
4XNQHqSyXZgbVKg+NGSfkRD9R0hh51acQo22Vli24nrD+2Nj3Lb8xNyaswOQtdJK0rVzqIFk+LSw
DWsnY4x9k/Maz33w8aaEwRWqVnrwG0Gq1XjasIdpDu9VeHLoG6CnorO5GeELOT2vGpbUY/8AWrd7
7czvZC9z47POiMzsUT+GYush1Su8shERXTG1K96eIvQIMIWQEp+i3zzIBTrIaWCOE7PAitI2HOde
qfnj2OSuF50uA3qKVYJ1WG6prW0zYET7TE5Ze5aKmK+Zf053tfqe8oOsV6GqAU0RvaWwCGxs5kru
h3jZygOariDZmElcjUjM6+wP1xPo/ANnGIDtYbCTb/IOoIMjqBphxuWuRnbZgA2qPjr/wx1fYiy+
8SIF/6dpez174YoN5PbLdr7kEuhD+1D5W3DbfDn39N4+ZdC9s4LWIznxyKuXJMUpibsj6YFEePrQ
+0DWIOjCtRJUQFrPsIjlI5YId5nt3CubcSauACUnUb6zIGB0p9gUyLrbPwZJ181+PaGs2AqyJfyo
1VxNYeqOIzmeWw/SyD3xz/2kOezUhvJ0iYeL2+YBjg3N/Y7NOFECiIA+sd1QBD3s9uZv1QzXWSEP
f9bSxyye8W6dTVFUumHdSsJXNoAxl3VTT2sr2n1iDgvwPiVUS7LW5dLbUQkBP9LOcgPxccJCo2iT
Qq/tpryE4f+Jm6s4bmXqLNmWiWcUJD1cRjlzghHrppPAQLj0sTzdFXeyRNeQ4DQ//2UrMysRdqAM
DhjjnjXiPbXG43+kFkccugqGD9iuCi7TZg+JhSrzBbA9iulx1gZcNMAWpTey/CmDQnfCduVg8XsY
ki8YxNcaM9MwIRJ+h7YM9nWje59fAvCDA9NRAOjTacS6h+CC34s+n/qtrWBfRe5eJxViLIxQR3JE
l/e0EhK52ZRwHtwLNi1Tg3OBg1l9hPFkaJKQwLw0wXte9R9nYOd9VvchYfp9O6+tFGKUCEgFfS7Q
kftXiHfROUTMaSim26gGO0SBI434MU8aNJX0E7dKI/lOiCC4GBSMznlIy6M6gR4IKRy+Vx/Uq8tt
uGbtBnELxAo5nya6yqeG/dGnLp1vrNc96gEnThx+hGluvl8YytQpCEfM5lvrkTadPXe6vjNm5JXa
zVXY3d4Wg5/wURh+/EBdOlqzWs9cl30ptSoBQSwZxRGbcqcg0ZopjuaCbKnFTxKzBvKWty4Ppuk2
2697QZWPU/uHrNMJ1NoakZluuJpUZLoBP9zbd9QJo9y+TIWi+pfI3nIiDLuYSwyEkXLzCvndkhb8
y7DVHRtawbsYaFPhPNZtAiJqoANfyWE5UAjn3qVKuOsHKX3aDHCNhc2QBuDF123dRh1MeDWtbJDt
3/OxdeR3c9gVl5UQwPFntBfxFv6GlOvt/kNS2BN3GQFKaP3M9NyRQb4EC333GZB9i1a3i5dyvHlR
fUAb1gvr+mwlVjy79a2r4rpv94H9FTDwlqR36clJbB8adzERVbF41MjPIQIUplqaaSzpsauHysSv
iKbmQcxPOEaKM2aypy/yGEH/5lHqMMwNyFSD/iemeMsZgDsdEwC0qjROQnTRxxJb2+AsMP4FZSmS
cYF78Gg6m8Ivd37+p7lY7M9AgwcGTScN7WcBZYJovrQfq54HK7g1sc2yamm9S6/QDLV4DhVPJQWB
xAgVTfTGmNCop8H1LwJ1uyn0DL0gTNGHCS6FoZn31u28wX4qa9kgIVLYJLdT2Ikx0vIuPjxWcJwj
Ype8NHAJQmcbW4H+NeuTA8Xl5thzr5nOLqKCK3N0uFmtcI3uqy5Tg5JxytnVTJg5eO9k9h8Z5Xo+
q/lVLtG3C/KyP2px/SDo4qVKXitxW98Ur1uHowhu4/ulkIchCmpAZOxWPpnAJJAOA/YZevgkE7ka
FWtSP6nFeZ32I91elanX4KKA0oeFv2R/9Xqyji0ioKxYIrEP+wwPacZ9ZLmHEDx+7h4Jc2v9dIRs
9KZogT36yopeIYooWbjtlfD88qqq2q2V9/jCC1APCqe1IL19lTKO2Cv1ZIiPAsS9UgMgrEeSMYEF
DAEJmVBH/eMlNdMUTD1a5keWHzto7eMVjeOWNqRCoEUbmSvGuGGW6X/VDNUqsscWPRx167QiPVDG
P4UB78wR/JY5gjQgl8nBixOtIR/wLljtsLY28ZZYP8xGf8Tl2HRWcn7m0UhPdQG0zQUoL8tdunrl
sTkDj0B7r4yksNgvklKqJdbe9gmE387NpExHTRFJFUx+N2Xn7MoeoqAC6tD4bnYkQZZTQT/aKydU
VWdThbW2Ryx+sVeTJiSZVeWvWUlpKHHHzy2tz1fMrZA1S8Tq0IXJ5HDEwQiFaXCKU38ZCUg5Tv88
fdIsop6KucE0Wb93KrlktpkRbyMYxjhnVEi4lPBr5edlO4VTQdnDYfp2spb3SWbFIZ/gqH6SUGZr
CAFzYBMjsBi1UcKLeyr4GyaqQ556cNtTwrU4U+x2mmnMeGNYOw7KKUnjWgeC1OkfqjTzMAiGXN+/
mLSEKyx29tV5Hm6YaDXXIs0T9XqlzjQWjm71N3yfju4OsjTTs2/0olFREb7aa/vJWdhKseSf2Zx4
8gcW6sB/yac8aG0fKfdekpsvgrqJnMRmvwfgH4gEK1Tu/sVEqV0kx7INAhiAV+xjwqoxSytW3uuF
jxzeM9tGjdbLkn7k/2zeofJSXLXHgeMSGgl2uF44bsA/NevOWzaAqZQrX39P4cWWt7W3k3IcMfUs
iw8CpWft9/uDPotWk/pS/R1aohvyviVGqVr+Ia/1n3MrnOlGL748FCpo1XPYavkmJEzq29/x1FGD
pINpSCyPA0GOKGOtWJM5Adru7m/drQelx/nvwpt0tYg7oUbByIrzKJFp+q6Snao5SaPylNJbsZF6
4HN5QWFZVf1ya0WYBVhWizFD/QyVTAIDUYrgnO+YVk82MruvvWI5folBMPk+EdiWhgvl7HAAbXYM
i/gKUzTjV/UQ0WIuVeTZ7szER9atnPHJP5so/Mdiw0tBt3A4y0+sSRgbFLoOVjwzUhGrjTnBC4eZ
0EcUEBCJHsH3t8wRp/VHGDVoUbE6W0Ij3XRsTpHtfLGe2vaK9aRH2aEp7i+tj2mBVLJ5BEoY8Bam
akWu4y3ox2ADLcr8dzcvBpIC7bOwSIDYbbU7uPNXAA9wwClgUbCkoeyGl34k7Xi6uvid1Ds+DW81
xmt0UMF0nQdYn62Jup6zR+x6cn72YSnvVYrcD7p80GsJnYan7TMRm/c2AghEKE73cBL4bpXNLv1J
edfejCRO+uO4c89ijrog2CHVJ6zbxFZiCchX7DGxlcl7I7TdHtf1CssXc5vGz2UiR1aicRIFixdm
XHBTBnIGH7S2rRKFxuPfObKq5bOsKo2zd65tPriABTPP8JZfxtdJ0Ua+bpSvqf3ZfNBYSkzvDwj2
ioti/Brw5ak2PgM0nIOtJfIuCSCclTremLTM9AiPtts3zYF1zRYtXCg/xwnV0SQqAaYuAuEGkEbP
pMxqhXJ446i7u2tCDMAoDlN54I5sUyR8Y7YMbhH3TzgfmriycJvzIt3a45PSfUSSArXFhhDHHGRe
69lhsTFW9VT6zZlkeniz567JlAqb9AdTcRbSIBY8k7sZNqXrVh3ZCVWM8Lj8omkSbPmp07frjDKE
sBA314PiACy8HvN1G//OMQLJe73TClO2+cafxXufjct1IRwzbl4Rbc9Z90SfI7Y7AhS9Mi867q9x
KbCTVF+YnsqKo0VI9jYZNB7Y10g4TvFV3eYPOWP7t/yZtqpl1eiLU0m3ziiewVu0O/MpBPYmO2Xj
neK/0ZJSiCDdGHw7ysgnLoBDDOHLquec5U/ZjIeaFX1AQbevv8FNCv3ab0PJTz83NmJFftXI1cNT
vTOda3Tj6Udc0Lnk2zNw25vpFomo47/+RH+CIXjGd5ySvsHiLTNDfrJoqkLb5se9ZqtwFsw9HqcR
D6LBUVMHTo0H1iQMX65G/0W8wPdFwrm1MW7aMuIdtlM7cIg0qByt7r8LldyzKRY9TwwSQdzKj3Ga
pPRalfrNI4QKtR3VG0j7pHKQ1ycbJdYCoXzH0+ba2XiD9qDnVfmghJOp6RcsiZdPIY7cBRyYD1fQ
g6NnTcXORGk/xg8iFefnTLFRA22zprX4I6RCpZlwK/HZdHJjdt4lif/sH2ErZIfl5mlXYmcS4Ok+
LnTqvwrchElXTw1bidwHR4667JRV6R0z/V6YrAB3lKRC+6WqkBGuYHJ0mL5bo0+pcN1YbzXM3TmZ
2V9we7hV/7FXwDb0jzwWMUYSYQIQ69nj/tN9v/I6tv9ulN62De6pqq8ouGTP9dqbD4/E7mhaWSkf
nNqn6lKY6WU6xraoRUP4vrKF2hYiTQZOoccsw160Rs5UrKlml6K7iFEw78NUG8LO2+EZd+uvrekK
/J0eWU+nf18oTiLT57KV+qVnoqbuRe1feLQqvZG03a+ONNxDBZ3EZAxNf1bSrEleD2Y3QeBlizEm
izqnSTzvZhKEF7P0i0RMs+Lbs44XNFD3aJZf2wMO6fivpxE0lNavKZ+K/SFcwEy44a+9+7pf2cY7
+CdUBBvWzaYsZUEjOqrBIC5Gaceoc4+PEWT6z2mm+dKxIKwSl0fbrrc1jKTumdSLsrz48P4F0jgf
a9/r+p9DMeZlrQheyu5VayyNzp5ol7ziflLzEzTYwtl9YCY2R0zIIyBQh7gDzNYwZdI8SFuSNSCC
tq2CDpDtEp8z7rwQ1Tdyp8iJ1gBWDxZR/OPbcEWcQHvTBtHz4C43FvcMfE49QGuIYPXanZeTwmRD
Zwk3qWR4BXRIcyIqCYQ4V2Bf6FEQB5kE1p7B9K8Czl0KdvJ5sSSfmak9mABeQnjyBC8r5u6JSC6z
c+QpBrYcc8hQkcWU2hwe0t7+W8kGr85QH3bwiqxrnl9WQ5SojqMH6s4iJoNBl3jY+lF7TI+jyAIO
OLkpKiLrUQzkjZVeQWWijcZffLlz7xG78Eq966WiiD+cuakXHLAcniTe7Q9sF3Tj56hDJ+UPBHQ2
dxmdd4U1Hk+yTg/kxAKF88ylkx44FG8Hv29bC+Gv3eqpNyeyvBPVOVdvcdbilPMrAArQL3c6YPJ4
t1dp71b9VHlJCPWP8vW79v5YLYLj7kOuzKFIjLZvzvUj6CLEmO6PaYasfm3G/xvanaP4EvXNBMiW
GS2MLjL+M8rc8t8eB4Ie0q309yHP3li1/i7hLLImZwWId2BcAIK2dWcvPDX4mzz5DhcaCi75QExN
WGSxuF2j8TujT47jn1xegiEIsGJ8ojfKmoW6MBP8A+UD2CF7P5K5jdCVc8C6XbjvhHjLiOGcDqXs
hnoFOBz8UMaTyNOuY/McXYwUZCC5xFnKTsF/O9BlpP4h7CLBQrj6ieelDspUxVHEhyKoRrOD28YF
gSE2BgV6mMQadf1i4wO4wFNu1Bjr8umNi0hbVuQ8lJ92W5RySghHEmUhgXMfX1Isn7lL6Xvbey6X
tg+bQfTtC3NO2h9hJDPF3mkegOllX46b66z/7F3SNRm8DyNzhmPzWe6ezjDGemDjzn8wHCI9EyvF
Zef1em+ww9G9VYqYFdMUn06uvN7vFKQQYdgCsH8GKVaB5MkMcbJnqIDQ/Kms4HzfIucclDIVqtwD
FoCgp2CPzhxBZUzt/IjKiIik+B2TgOKL5ZwS3RaM/KlTeWhnnRM5E+Z71Jj5sCxjmQxDG1XTewT9
wI3nnOxEfeg9eGrHQ3e/tTgbGqxA/GONtNf4zrQOnP0P3OdIAFeGnZisHN2teBYlCmS4RzU7WcX5
2t6o3c3m+wMwA//2M9Mkc/NMoqrfOBM/wT+pIADy6TFHXJzWsSn8dJiAcSprAt9HLMQweUyhoihx
YFpwooGYjVN+TQhCXYKwlF0tvAxHdnxEmdu+eBxHqlMcJhKsa3aXk/V0Acu+YQwcHehqBml+KTt9
SYEX8JNeaxFQWd8jVXHZcaIv4As86fngsmTqU98hXauCmz68gZwd4RKBA01Biv/ino7CetcoeJ09
2D8KL/Nn/SN+tW1GAnPLkI5Ldr8dhGMc0I7uyNUibkpZ7shhnt0apeJlmCaxMBavbgmgRo0sv/+c
moCoBbMdmP7gb+IaZCU7w4SjUP3+Sv1vPBh7N2ckWedEEerWWPAslx7E3DMa2FwysTXfYnK5r50L
gXAyZl3zP7VdYFf0peHsSeA85hcldHRGFmNH3qV/6JKWgm+sqemJhw/C5WNaEBrVtauKGmQbmaEj
z9V92ArDL8SKLe47fyCcVVlWXVcx+QyVUEOshlj0RTe8Qa7PvP4LivDwiGK+F+mMBuJi7m9l/hfq
BxvutiCcnR7eMhGZxpA/vCQrK0n5qYahgCDxzfGyFKPrfbRzX2RzKMNjQ8LU7+DNPEvIbb586Ekr
EgQ3sTdTsTPzyhd5Lb5gfRcVWZ59R0uDpTfA3Y/NzmcMSHtO9RTnRtR5iduusV8RwsWEps+/GKj2
I2h52LveM4I0+KfQqsljCw0P1dJUUJSQcCP7sqe6lo4d/I8+w1oLII3EsX3dRV1+bCHhah24BAhV
z6v+T5luM/0x21ivkj0L0/1mRKl2QOIbBlLb2xaZKbSE5xE40jKjSTTnXjfxLAlZ8xV3viu5gNtg
pmkajNWVkiJNvRi9xEsDqduGHGeNj5Yvui5FrDj5TrKS9+MNh7cl8EWjxKGVUlvSD/7r5DuzNznO
0xlE8xI5jOktNjKzzGrB5sBE58U43VOiLjZcU3XEuiVfvW88ZnvwamlA/jUe7TmPHt7loYNvBAWz
TwtNpwT99fyFFWUhTqQPKsKKNmdlpDe62LoQVU9wqoUrOIrBkjnR+N46eZeMNNL9ITVPHjoIFpkb
Yh29fjTrf0JLJ0Sv9i8r2vvq5kO0/un5XrSVZ5HzmJ6yByUrAqD3KOkgKSLqiSsFFk23h7ErhHNq
cZrzp3YbPsaPShUTToUItsKMLmrBSZ/u1kcnT8KGaEvyuXcoF43flSa26+ntvIc8U1WNGfamN+dQ
ksfG4V6nATlNLsMjSmX2OTZq9btb26/OuzHqZyNwTn/hrpMviqIT56RajbMMLZL+BHAb3Tiq+sDZ
w9JCacX1hP8rcslUYUj/roehKjir1P/HjGv/4n5VbOvWc1k+Irk/DtZ+Xef9Zw7X6QSlMpPLXPz3
y/JbZY4zoSuL0CL0+S5bk3gcLsbr9MKqeQP+VfH06JAbldazd8Z5jFq6uK1wpp5MHE1dIdviohSp
4MbT6EpjAVkNGISfwjwtVRH70vTlX16cb50FVMN4Q5ASHos6BZZKz/qQMV9tYPIoWdSfS1M00aq5
IGHUFcr/B7pGtNg6h6qw7gs2Yyh8c2GJKtnEwrCMjKGfk3ld44HyGiArrTpkBkHFghXN9i3cmFO1
yT3ZPGK/ldoEIf7nDUinRjopInbcgipJKzGix2pwtx5pRxRqXUe5Auu5slV/nBDEZDgjpkhL/Ps3
w2qj6SLdoeLACUCsJ52Ng70SLArp9VtfD2ULwAo92zNf97T1a9tjJYA6T12hhIqwR7hbx8mhBQcJ
e9HYHrucw/WD4Jh26SJGwhLUUzqUvmRhSztwgqXdlCb3OhRfjrt3p+Vy1mEoATguq/R0mTVL3qSx
1DDC2DFKNS1xpGO6BFBglLfdTlgr86804kxkgDX1qxt0wW+9vquLSj5XKPF/C4GC8+J49e9L3C22
3cMpJ1jrpzPddPZ+fdRTEhplaZykPZm5zCdc+MmDwD4d9D81azUi2P/gVZBYtDfoXaB72LTVpznr
90x308ZspklSMKPxRFFDfSwV8FDFIccVwMXeNBju+boHCJdLGDGnxZ1Is1Y5WTE0uDl/28WUo9sW
/MjvqyAYL/ddhAk8aHjZZZdhiKlZ6sWirKDRQ+we47kuEwxKbqTe7/Ux4JyL/yzAa5hGQ4v1yjfz
5KpkcinNB+JoLz1rjoukTApwQDhd5tVsgREJ0JiW24WJ3IP0kayO40kyWZ21hUP1FO786LDjddsZ
zc6ULXYEpd2rIGden6eknF91YFjX+Ibz0A9HC3P/W1rrMAVRhl83TmtWqKOLtSibR00vWscufJck
tUK9WNiKs6kjx/ijS3Gj9/pFPdOEEV1xRyFFsg6FagsfW2ZolppFXx7+ALvzDlFmDICDxuFP4mEA
y+UEa9CY3ejfhCgPjtg+S/tlw4Dbrt/7wlVUAz6QFVbeTifrcDNwKvJnl6mewoQRz8HQNu24f0Av
7Esx2SktY4gQKGU4uKfa16ET4VpRajXz4jzCa7T/4pxXM9hPg+zpN4GuIcmqenyOhRkANpbRdWPf
NWqgir8IdlD2uXRUl3AINTaWQ6CGedOjXNONaYKQHPIYLxXOsW32liukaBOSjvEIJbhIpNwrJdzX
ZUNbD+CJal0FgWBGzQmua0oHzNzvVvmdVo40p3LwpH+++6Gge5ViJHSp+hIfrfcz8qvzm2x+Bf2q
n2AT6blh6WfpzBg1zMZc6wYh1pAqGz4I+katF5diIQpuGQu9re+8WZNeufgzGvjvtFkKMhToS9/7
ENmQADScRYuOX0iuvF0ppU8k6DJAuRdKrK1vwdkQ1OLkQayNQ8wFSvj8gDdv3z5LneAFN4pCdiMn
QiSDeJIC6dxczti/neLvnG2g6N7KXSmpBx/8E5tIWjUx3H+dQMahREPsNo0aksqeoV6KPf1Ji5sl
4AUE4NimPUUdFgQCyxyw5sX1FISxu0tX5ZImBLkoUTNxin+uUbyZP9S+r//29UDrgfE2skQL104X
NX5XTfEZIGBcbU1LPkDYKjZwC12wOyyDah1kDf4Xe+qOD9cfwefsCb1OpmR0pZSbsgvZkhtOG8j5
kAVZJEwbLH7nPnB+BTw+T6sg/JXWYx7z1XHOHNP6uHWpQlLvMcmNdQybBoMYtkPWStk4dnWXtdV8
vXrXIY0noceYw3pJmrHPzEDdSZDFcbqR9TG1LzVzy5qho9gUxd4rOiaHgJJ2P+Izxvz56XPtS+q1
J1WYfai9Hm2o7hdCt8NY+0IVCyJPqEC0NRXJJ85dH0DjoPak58DrhH9Fqwa1VuQ3CBPEjYvYlu0t
UKAwImmXOakn7lvmf069Wf8qryGW9Aw3QO7pcJLW9k6TEj6V6iJ0Scrreyj371Q4Z8s7WTgJ/L0F
tVOFlRnBbU8gZOMPTJxLPO78zd/QE6aaCm1UNNNXHPM50vydJ5RuO1kk+/JHzeG7sF/yHmbfXWFC
1YYhy1aSQPCxutuD8krpZIuAO4SrnQoQgafP5NrbwM+edNh7JODNoibv0ldo2kBUlKfpqmR7JBou
Pv7BJPfb1BT8QhNlP7uDnrpxWh1VAlBN/eovcHTlzNbDI8V3zghA73S2nH4HNpNIiuZX7F9GZgvG
xGnhYsQkREdMN5dQDIJqkNRey43NsRlDUmmy2gIOq5yW/nrdOurl1movQjHNrapxAv2mQ/4soPIi
E6TFY3Gzi1RsfR2DqWmRV+z6GxvrGhg1hGEh4oKVnVhch1RcocUetlkvVKupZjyar8/l3grqU6js
9RWpuDAlywT3v+yI8o3fkeE33svQfZZDvJgpSFD/WsY6D7TnExwtFrEef3KrG1mdwTto2AxhYlQe
IpDrtCJouXUuD34O+HaMeBCTmFL8PM0YjPzPavi2d5k5oWQCJktVmsUbK70+jfG0hk9BNEfBke1K
7ctmL2geMaYIB4qwNF7+kY6KEfSCNRNen8cfaK0mM5ym/aplm2mGd1sAsBNZUilAGXzEpeMrIKQx
/qMSnNUwKr0ipGzLA5IDq6t2in9w1t51mqbVJDcQeW2rWEcOYCRK+FOrwLiaudZgvl5+bUiFUp7z
ex1tC8hFVXHD4DamL35/3SHHkrFuLvEXY02Cr6z+3CsbKSW32VKKs4hLHS8kUHXJj9SXo0kiXBjr
oxnC2okFVKIGFip4NLBxesTDuDjDSwbeJjoXj0TeLCPu59MP1gRso1/DNzU+Ptl1j5r0UZtZ0lTh
PSk0vkMaFI4x2kSdAUjddvrVa5mc1D4gVmUmD+HKeCZkSn9U1M+jM+B+kXVXltjZ9zpI2tdxgDuA
nPtXRb7hMOCVW/g2tUksyL3g4qvIiQpf3du1eajmDbrvyzY18rW9YXLGGC9kxaJPKvMl5q0LGIvE
pg9j3QgX0lkrqhyPadDI+pDxR0VmpyEEZ9JFB/h1KeZwIpxDIb4HZyZOOF0b/N5rkqXgO6jii+5s
DrI39+6lEIAmRDToi7pjqQD3d8bHYt2MlvqU0rIPfHdHp4q9kIMSlTY6kuFoldfq9Z1UBKjzP43s
bn86AkTtlfB8bawZlvj16xefzqZiMO5ObcGWuNWmVqTCKlPo46y6QaAWMbRPhsVDY0Z7J2XppxnO
C9F/GAu2lUFNvtp2cZcherMNeWLW2uE6Rl8GU4d4dmeZCeDrp0SgMwW+Kq8B0baRMwvvKXigArmv
2QcfX6KnPY/bcgqABZRQujvn2gkedpl583N1qpy114bRwavQK+Iy6lNQoY4iZfzmhfb2QjTstydt
oh8oR8hFl0yCe1IpkTvSgMb2QOJWOQk2crSphzpqakLM6QdlzKxYNH11SBICRXiPtJdgKE91V5GX
3GiW83k0yNfYXpVEmEdL2LrqyaGxgWKx3JqfjXKd64Nnn3V1rpcoTmfuK4UfKCov9P31+GWb5Fju
3cV+m0T0nFTnyZXAChef31c370NxXuUfxcteJpexnSIvPFkgQgyzviFyJzBtMl/ifyqgLUqHt67M
u6fBBeI3OXgkcFCCvi1kr2muwYh/AUXL9C/pnmDoKQiK7lrIhFAEkzNiaC5sMvhUr1CqlyxGjBxN
LTaPXtIAs958Mwjd9zEB+F34AnDY4coxPmZ7RnM7wf+fvGEjodOMq2cI1nuMLQPuSXcX2Q+FbYRp
5Zv10Is74YLcwN+BJdBD1Q7AyVPXSSVL5PeeuiN7IwNkQgXM7c1YArotGNZy17d7afDLhtvbqJUY
9Ki0+mOdTantMQ2QT6DauhDrEwwwybIPQ4zapUs3hE0Cu1ABMU1kpFlRzAuezDUtSttv8Oif3qBX
9yX20sN7Eq3ix4NIcNgdKa1qhy/JwC+UDr12RcSD6S02zkm23piBdmAbkcTelDdGNsh4n/aMC9OZ
zZnI3ouaRPgCGK5tOBirHOatxh2Hk6PgWawTcKaeFYq7JO9c3K/ERaDvx4ih3rlKilaAV9banri6
S7kQCTaWIDJCQVn9uV0wZFuit6QulXoIXWRvZecx7V8zRrp9FQ2OP+J4wWO3yIwW27l9h3cZrE6X
S2e6ANy6ZArNxrHRJ097ZlAyD3xdekI0uQPa+Y4QPiljyyeQK6hiUSsdo2LYmaB3rdUj9nHBatgl
3OMOnCmEiMctsmgTsGZzL8v1/xK/qO2mGuS8nWLJ5KmAm50zOT3lX7VCueEH+UiM0+dCvPp5FIMC
SJwlDzx6H2OX1WjSjF6QI1x45k/pwhe8xUVeF0MlQlerjbtLqK0rc/Df5mXZywOeaCULimE3zco6
b1qXIUpGBrZF4Lg2MspT466DsyRmg51M55xmFHf130hQd6b8hZlaG2u3XMPpLEB6DldYmYNn7WYE
FO1D/0Xe1Ir/AMeSsdOECPRTf2uig+6TP7jrzCr0JCTS7gACSnBy8TKiYgmlBOUOog2pMByrDeME
Pycfj+YWPN/zRCVW56kEeUExxj6mUjKLuso+k2ZnHniSgH26FY5pz2CP/2nc892k+bIv5rut8jBV
U6RgXIL9x/ABZ+x1EDMZlgSqKcOOAFcDuoNC7HCWNKZ4dYd5lgDlZfhisdta0JMX+5qha0f0I16/
6LEhrom/Fme87kME6duMxGGByjGdZ4zqRWTe89Wea7+TkR+TiYj98vX36YYOvcUh1VRamF/s7ivq
zng4dwHm2KOslANoWXKsFNOXEJgK9UJOnVMZIr6FZUE6Yn3+91zKA6LKhO1SqEdZ0WkI7Swvin9s
xSP5aN6oWmbvfLcbMFYah0yd7KHcwhovEfKhlq/MVe5dYhYqe+wNwWbue4j96ifIAzB+PMZwBW4E
bgeVqA36MbYHP40YKGDagABpmsF0Tdyqt89YlPtNllNMCtLq5vBtlvk8c72GN+laAlMFxXlxuUCd
Z2QaLHXcai7E6wu6qZleRuTohbkbuWkBER6F374vodtgDuh2D3euYLNTGZLM22zFi51ywvDqdMjh
5NosHECgyxVb1cQqoMXgrOXpKH6psLobX21MMEt3eCN8iSMItfQEywQnEH8yJuQKP1BCvVkVpbNC
HKsQjbSSG7amTe7RusiBhObWNQI3POlEpechuNd1ntRbMCSKHII6o13PBf0++TD0xHWhd5/UEfuZ
QBcSuevFvc/Eh2fh8xMDfiB34RJuYxj2S1g1AZ6+GrCNfjuRgaA/WEqzlUARRnQiUA8ERlRIJzGr
ZoYJzRtkYiWY4EWLb88mrhErcz2FhbtvZugZaRGiIubWzct8uiej0pFslMZi5qSR4/2QuXI7Huz6
J/t/df+MsG7AzVZPqYjBRKC9scRkH3Qu3uRJlfG4u0YSMu3ccFZvz20OAu4/XW08tGdJn1rM3kH+
AnFgCpQc9+Z1IzUoG2tKjjBkYTc/eGJmt1WxYmlPNp6leZ0XkPhCbHzrjvBindJShct4QW5bNqdd
qpXHt+jQwBCacjWK5U6Vz3gv5QBhpkHJrrZaxI50qTZbiMZvYz5Bur//gOeEyONPumGmKqXx/DGr
2sbkZUb+nRqJcmoFEXq9VhlYhjdregxT8I9eBe8DIz165fmpClU1oDpSf1RX/h+gvka5cxODUald
yk6k9l98RvX01pLARU3nWDQStY20+QUwghDMxhGusLYoNV8AaXYfEcmYU8sMVu1MBqcSEh3JBpcM
bgqqqByqKTz2qWqpTDeaeqhgZESGwnZqXpxvaIdFqazmpowKQPl5JvfVr1sAqHN+WS7onHQt8dBM
U8fmTUCKyEC47c7ebiXXDAXPkHdFXr+CxT213bHjut82WsKlatVyqmmcyF4eynsz+mIk7xt58yEY
9h0jCxhekOfTmjDh17Pi0/3fWhcJcecfdhACatJV8AZfrfcOAO8pAhSTdfJ/1BG5iAGnDRtb8+ko
COpYlJC5LCGVxiua7x9EYuF7dGYALxsxDRxW9BmBQDBgFno61+KsMP1FLvEY9F6ztoATxHDTQos1
ZixGqU8jyZNWIWJdfEOQP5EVQ0ynVpx94cwH1+ucohUJwQ9+vZhGj3Vaa3YSs1IL89JV4oNojeA4
wjKVBycgp1gkCrZD6NYCCxAgeDVOJx9YYKLW57e+OnlKXV/wDlpdyfJkimH/Zqa3fmMU+M+YFJnL
VjUaLpaNMgSNqB3yPWrRwtQYSHjjsBnDkZqsuu7RakXTwBRp3/F47XmZup5GO1TQAVYDv0wwuc6l
DvR+Yvl4gKEKuBP9yLOpryQBrTjlLxIy3X8FxoY88czkfS1yCziDAjbJ95ZPu6Y461ZOIgki/k42
lF3ATtV4dewe+dCDAET8mXlTepn1RkHJb08QywDJiWujcEReJdjt7ETMoDbTMX4ohPIXZuKdBWN6
B/uxWb8QVia/dPASecS89l9TafUAr0cigWSeHIaZvGY6SE4UikYeAxaiG8RRn/T67JjU8tNVioul
4GgDfWTX+RXOzvfsvUWrj0M8peAi8nwfqJC+wXheXOz6Uh5TYaUSy7Z3dQEwFzUTTpHebTxSbhsH
7IYHCKrwXTx6BA2Wdt3tRi3TrFTfwuro9vXU0bmjlDwSDXtAfVbfT+VjwmFbAloEpu1fQqkfkQj8
fTGKCUX0NJePBP1skxUaMJwJZ4yLuCKo1hdrDL/fkgEavyAK65nhKw3lGcljFrwZe6mqXd2F4mnc
DI/kNEsjCQfXNiW49lY43wWwFAwowiSxNuTZ6wocmEaAjfrf65edimcNYEOJ1C26wVQxKlagMyLv
wwciaVPOFC8mCVWBWabdEOqeBZbrizuLTwOUQFR+bHi1sgDNzibkICX3hTs4vlRj8ek9LOYJclsQ
pTdFuShAuFUHTD8TqNsVSEWJ1sgBaqpBHOvoetCe2hpov2GbE6lL2QUB11MIbXsejZ95pgfTFaUf
grFua/UCX5mzP7JMjc2CD5PInfyRiSXqDk7lCy6vM3gYikckzvQF8uyvgefdK8pn8LG5RlPguEzG
HjF6wJwNCORm8jwKb1PaO1CysKhlU91aPIJ/nXXmE57TDKYdiHTtMA8jDltY7LmibXItekkI+89Y
siRN1nJO+5//9juF7ybOHb6TDvW/bW3kyJbQ1e06Fa/+dSZyI0/zqqdeBWzJY1wPqE9XeVSRRoWh
n6h89jRnp8SIqbOBrEV6ytgqpD3h6YGXeKUgEifAiC0yxuDCa1WKhaqTfIgp/tbEmgUzXF7fdGov
UkWT5PaRKC/WBOilP3zT2G82NlL2vQ9SP4Gmf/E3F0KZ1zgWBnALcDKQZ63KrtKoh6LNf/vlSwyH
2N+XHyIUqOWebj36coJDhk7WqV5yQkrotCbnlaOFNcGUqEoZTp/kdj6CasZh2FkN6f/2o8YiOWOn
fDs68TSY8fnvg2/Bc93ebq5Ev+3aPtM4PYbEqeWfP61vpflTEAZQOtJ2sopqrduyuRogWHL0r73J
FHzM14CdjFnVQ/sYIrJ1F91F2OU0VG2WiaVunGc8hkiZxqyy6sxMXA8k1pj99GSU9hDRTeoubTiU
4gnXuv5lIwA+qKzRflFp5759U32XpJR3tMizk3LDsGHfrzxKWPQhVq10CaohMU7jZ+ASACCLXlbU
HjacMoglRePohZwV8TjTWfpxWmAR1BBJylFdPtYb4htTebF5JrLRyiumHmKTymvmgDSm0pILpPl5
91xBmqiJrNh4eaf5cH7O7OgmM5OOvMJgtwRGGVb1ud2Q6I2Bq/ZfzILcnHeHNk/n1Rqduacti5iB
5PSrBTeochGVo9NGo2bAVNuejOhWfh+QFfC3jXhifDYnO4pm4kwUipWZz4cy67naYCb6lt+4txct
SL4zntiosV5d4onnZlNOMFvFPLn2P3h7tzSOIF1ndJf2UNsLjPnIq5pLHuRaGlrudC0ha1NjaXg2
pM2yanpSScLgmeEmHOT+AMtF/p9pESBRwBct3s9z4D748aXTO5R8zJog1obu4NknNj1LhYONz5f9
D31ZRkSFJN9EM3c0p/4J4PWjQ0Feg/oxsyaw7a2wwYdq10uk/A77h91pvEO7PurQs2WK98zcTGj/
pqpKKrPwt5DhvFRhHa6ufWX/o9XlW0ynljQkJHjtFnblPsFehw9oA3iQU7grrzMZmTHKh9/ImWAZ
MXaq53AcqzKK5rDnJ6IMe9Ut5FKdI79FoCNY0tocNfwVerF7h1MdIWQfTyZPhCxS8gGFm/mRw6ix
YsSMLCl2GPfs/eHMqmm1I+7S/oi0VTAWvQWUlzldYpma0qiNf7zjW9Um/HYHhxz6M2xumFucr8MM
8sXkNyoSSKkCQ38dLIL9vRjPgGKZLB+bhaAHstnS9jB7YO1zUTPCRzweWFoIyk4SwFNS84th1MX/
ZjHHn+f+7JZ8lFlChmZcTWNCWOB9nZLa43x8BHzX+jETilSKk25YAlD66wtIG5BLn3+c43z4UYTs
7CEA4AU4CySESHh6EvUkfNUwzB7QTu1qtnsne8jEkDPSxqcWAv+lD4dmSbLPm+advFzxt1Wv6lj2
3Xrl4tXFcfumBBUD26+Cj1P8lQXXtCO9ASzJ+APRTy8VKwhVxJh08HmDzK0gf5RhtbJtC31YUTql
b0WjfG6KPJL8zOcEPcz8kwRFCe35WELXDc5SDlMAwZ5tpxROD0XDh+zOPRUHp2mQ7cEBkECe3Up8
ENEwhcfiNx+Vh1p+rAqL8wDGV+vDgMXnxlx4IYPqpOmXqzzrHutqOCgMTo8ETqBfm7jvSz5wwEkq
5tKcOv7/AZxM1Uksniqk03/Q6OjjlbcqmDC80vCH8GFKV6Ag8vKjqZgT95WcUK63qk0e045szDwx
+UXIHWhZ6gCcuCHQFYXTnePDhLjYawIXv0c4utFjTBsRl5Pq9dDV9peDQrTifU1VHCoGNS0/EVmp
PyOhUA05SRzinz02letrfszlt5ZwZZjDvUjzMn6sp+vLo7NOfBtHG2voHh19SKdI/zrALxipNGV9
2+9YxhnJJ7M9L/iRj/LdQWvNjrub+WuasWrYxajW2UkfBV/9EbkkuNi0dIGP4qvjZGlIo1iUtJy8
XN05tcXfkMO3+eLxtSV/eI7XogZdqgDDdx9ZM2MswcSwp3voaK/UNE1VCnr0hueb1E7Ao7VbTHwO
6Rme9/F96GibQIjunIzODNFJxoEZTGcssvm2pVyrubbSLoIiUCWa2gdNxk+F2SIXlwsdIuQn6H5z
4Xy+QzdhKpW3F7QV2Eq9KNn9JxfSei0vyCZ6jS3271JmwT9m9P9b2a6JHCO1I6OYKkHRW2hzrsVp
ySJZkvX3AZOSaqydIaGTgO9sO7USCZPKtm+8kJjBTj0vNhZJf/No+e4L91zMXtSRNzOHnSkv0cbr
ckfMHbMTBPiemkh2NqUWRaooBehgnTKaf8fe8swTew6h5jPcEMt7NRx3yUhw6FcNwKrtuulJJQ8l
C+RJrBMWD2sgCbEeHJ0BrZwAmT47qDA4uihvkmtC+YkqRFdaaAAr2fyX6TnkMeJpSQqND642VHEh
sWeUVInSnQfgqO8ZpjDEqfBLm2gWDeiUo7kzi32MK983NFtShBSfLRY5oBMHCnpSAyNYOZKhs/Ud
/q8hb+JXER7dHUAKlLlouOYFLycrqToqyf+woQ7heRmzIhJxnh3Ztk4xUNO07ewi8un5XwhdSD3h
/mNKapawMq0nTrrc+FlPjvCekiWBJjckMYA9fYeLgF1DcJv0qBSeZoW1SQuaq7uP6kOgnhvDiSJ3
xiWDKvSWBj+/7e3B+Ai4ei5kQMWMkEQvkrTjfRwbCCGsnWKQdRPsfoFG65eywCIPGCWyCdXVy5MS
gU16I6rh3r5Dv8KDG2Era8DBFRTfRJfl70me+z281iOouOfOezIfqktIr7RkCTqR739gUlof/GpP
c1V2xlbWxT79sfU0X9a4Zy68TR96J6v/228bwc7wtXybimPsMiASg3IAant9QVU1MX/4zK+9gUpo
XbtmghUUzV7eWW82V4sb5EmZRdzB2B50k8W7wzMG9Fd2THPA4ab6G33ctJI+AaHFXMz+QkXiYf2D
NwxZzNYzX+K1bom/tRsLcdWfqhhdYYxIE6hhYXyhqnvQA+kpMJ/PZku9jTrGbbQypxmERlY82ngl
uIwcTyWSDQsssLBQCrAaN7kgEimXW21QuPj4SY/dHMxyYDyvyL+QGx4LY3g0XwCwh+5Tt8227ZjD
kDeE04h63S1dkKgUe64FLGY/9FrTY09NCyadeCb7Ks3JiiWYqlNvpcStHgmMGx3N3krRCwfXcJnG
0xBqD/BGUuRL7U9kwonQhqDlJJ0oFrKDDC0DL9Q+8FOgpC0KlPYiizFKG8X2/J/vnZRTIsicVv1S
tdtr84hQjpWZ+KYsmnb/jToRpJ+kXL3na2KwnwCmAOW0CKzj+TNl/83JL95SD3OpaYuE55YuNUiO
FXgL9DH/i0lhdJaVR4NJTwSmc10PP0yrtAVFTnPxyNfW5c0NqE0GlBC/I8ZvnlM6BER2EDZUmbBr
sudbfuqqMUvGJqbFwbh+UM4X1fhpo7KtaDar6UM4n3Qn6b+jOZYWvWxO9cDCQlTcVCUJ58dtyaWe
jt1AQMX0ph3y0cEOr5u4CavVodm9B2bu9QZgS5tcQFmG/eqBEZIFw40kHEGcXK0WY5xDL7O/g3Tz
mDQeiOAM+/idhgLBK5fYkAejfOsE94qkelx1OOvhoL8L3agUAYF1h2I3PCfKY30Jl60TQf3R8jpk
wgYuV9vpUy9rs91ijmXeZWQlQ6wMIdk0L4V/vAtg1r2dHUPhH4FlQ82abIjD1FDrrIzwYJuV8w/m
ZiMs9OtI9z49JcwUcYvV1BP5iszneM03/YUmcEbPLuBTNqHFQZFLOUAELqX79+3eVcb/9pH4GLL7
halVMMdyrPY5aGgDmHJLdRWUYJIuTZRAzx5wcx8214is0TCjM+NRM3PJeb4LYDQbh7S4qj9MuEcw
NtSXN1z2O63dZ1rf9bgPULmsDOrHM7XqLx04cPdPOpfVvmuzUKkiPx8anNARfW4+SjNE0XYnB2gR
/gmbCDjoaTc718yQ3KUzFkgm9gNkDLbtxYxw58CkApJ+C9gQAV/Pbiptqhb5e/w5DJRBBGNZlXsO
dJV5PC/S12nEI48iSbWUsxEs1sdn1Tgqqc4v2infTdOrxu8FGp3ufgWWo+mDYzfn6WqRM9ycS2/j
en1Rgi5vHvyqQdQH0fuJKtBLqZ4RtbHvihFt7nZsl73Opi4k+KbrVAfCrdCRdOVSFFLYTpEGi8UL
oflrQ+LV+6LNZhjGTKryXbGlUPVuj0emSds2SGWgBWc+HjrJz0BNuOUq+ySHsWmqSeAj4JEPCJt8
qRNJ8NH5dDr7/HuWiJuR9QNX36c1f9irx7d22XzG6Eu3rnuHy9Tm2NaeKvzBJ6+UMvBiQ1cfswtn
gIs5qk4zL8FgBviXufYL3s/IFobhgWbuk6XpKzp6fCEo4v9T2RalCy2MF7jP6InOkvlOI4E081gG
loPeBLJbcoRZItv7maqibrx3pBzfQ00DguuMDNrwLvDQdGiJdf3CLXKuU8OutDkw2bAaWb1QwTbe
OnbnUqRjrS+KAh2jaSfMVA+71Cc/ZLvy9qvkbmj8CbTtS6NUIc2/uJeb83Pdag1oSYdQ+pACpUX0
0j4LdIiWoDiIv2LO/cXQx5ky1kWxMbcPgoQVQE0lZrGUUfwqtUAmly/R/jis2Fb6HnOhdNaWkxzL
97SzZB+NBg4FoMQSGxcJxYYSCDfBiyhCjRYb39SeJtQnq8GQTglDyWeBToGHqknMT9/4H01GT1TA
2M0JL5NTVCe+b7zgklNltr42HHewganEkZF4NR02RWjh80MT66RbQwjrRV9hpAJkzVMzS8wVSDYx
eN4IacDiUYtOoe3W14zqSHA84zEBH7WzZZYUS/5IqEhE5mQ9/wG9omxpLn3e4mMhCHKyN502xM+P
GJR2DnefTYDU9wWxB6PLDNm82hcg0RuqZA6+w8jLg2k1Fw8mAezFHE3mbLket3yOxKIz8rSJ8V1m
O3ly9vHPRaqZ46Pg+OSzWIjqKJr/v2SyQWHs6wW9J6LU5/jsVHzSxVZSXwalnqtEcxZlwLDu2Qxj
WiPs1IxHx8LCajFh2XmMSifzCVv625XQBSc9LNdF4n3OuEwMmi4MHo/Bcr558nkpcyaaVHDZB00X
GMSBUy/klVpt2vd/IvKdXaHRuMTVT1OhVsz8y5elJ2jpXOouOz3hng/zCWGGiaCyL+ybsSCjhwYR
vwASW6qPciTK+MBY6UF2DMsJlhIfksUba1GCnKt4BOlikQ3zIkrfJ8WJx+JGf51q2l6uCq8DSx1o
QP6CWjrCml5w6NrV+4lPLoCqpsKWdPAQZtn4qqYeRjrRabLjt8HuMkdICz0WZpgNXI05cGUtlbFs
ILb3lBO5eQRKdkPXuOogxwq+dbMgDCaxxLBJahULaqGYWBYsPto7n3vBEuQKwtZqsNZSBgm6pi6G
+ROPlmVgapBrcnK69UoilRPxWcOMhZN5GymhbbCgPl1ia7tncym5wihLDuEfrt6P6q4e5hb+LANc
lrFjbKeFedNVlgOibvu3qA4xywMNkgLnrYM3UeA41idKb80k7UX4jldgc3zAf/YxbZkIpHu2dM2D
RDT9ARbgR2NDxNMLkCSOIylxJT9c4uwnCHjp3p5WZHooaH2fXEQkEBGMBzmdRsGqRQQWaP0OdnPo
BhduRHGfIqRB1qa5bRYcvEqSW4/uWERps54aVFqbtG3WO3C9HepfjZeKLwKiAsgr89uuIJLWW9Ft
BZlPksiKEjv82YOuqlLLx5H6a/1ynRrkd3nvUYIdr5PEtdR2oToLtrn4Cof0nXtvw/OialJMnBYg
Uz+Wu2vzWXYtHfKKQ+EmAvc2b7s4H0y1CRxxeY/ZdLhb4FFABvMylIWFXM4z6qHvsjBpeoyqplS7
OKrbUuf+VWEG1MGXsxUHHi3hlUPgMrEE79wLyHMPBwhHri9q06UHaWB+sylc9FOMVrpIxmJGoCfP
t9ECwpHMJeEoMrMgy3tAUsIIBSPnx+pXdh3T4qtaBq1YJ5wF6HMbBQ6El2GlmEgyQY0SsCRrqFFr
3gtpHyeInp6CG2IqBTQUqlraHN82jZ05kYOOwPjVRWY9cMflTWcEBVblBev4NsR3VmNnoqBessK0
jS0O21V1jOFXIg3vYvqHbaLrXcSNTElzBgBa9Sb9L6Bboy9LWBVzQmp/5nVfE/bH7ycvSd1NZVwR
VUaLBBhEC3dI3TfwTSXhVf+3JL/MhnrrRIgmSdeDvAbE9nk/16yg1E5NrOoktfe7dOcD9Gk+VXaM
KTjD6mNn/dyDNTqNBDHfVSAx2EDY3umqs1ElY8FE5/GiNC9mrBY2S3LyTuc9UBHiFhLJRj2dUUaZ
RSFxd7itGKI1FmDo9niC5qwl4JcTorEOTN2YvsGBPQWxDGrzuSh2YquRFXDVEyQhA6RGoQUxMJCI
Pw4Yr2hyTAI1eM/HOSFOw2H8y3DqX9UMh+YhrdKT12TV4tM65K0x45nB5mrGOxu6D9PwQXJcq9qn
nPACXSkuohm14q0Qoz6PCyOOVZOGRHHOQvELw93HkxsHIocraCh9YeUILlZUm1XWXZLyhHh/c/F9
bHIxrne1uyqqDNkTv3gu2VC8oqQIMb3genN28o2aL8toG0edvXTf7wLMzlIAisk8Z0YNrV9jyu8E
09Ue3oxnrxUXOJOTswmw5CQO85lDkOjHnxNDXbegZQxLWwbelGglkY5YwG7fXYxBbirnU5fGDq7o
23LRAoj53Er9afiqy9vHYCtcvZ1j93r27izECNWRCirCNVwzMt1HHnBmk3kf0TEt0IKrzz0m6pRw
xjZi7vjUNRPrTokBgL/mCcSv0bP1PwwkZ6HbMzgJLfRyeCST4Wc4ByHAr+rH/EKcYdcSSBT3V1eX
QCc9oipxI7NlyXtuDQY7qYOq49I4UBCwtYWdbsMWPxVIpTsaStdki+Ov6BPQ59ZVH/kC3PLlT59+
WYyM2NdBWtw0jK2G65+4Y3fASiol4d2KeiCbvDi5Ld+vSKk29ElRzwvsiSCSS1EIdX3lfX2khWkE
Z8j6lVlcBU5Kffp2qd+QxQl8Evh2Yz/HHXVIJDic7tMKb1qwvKDglfE95kYYGHc3VlRiK/h9ODFg
/KHiiEiOjp7B9R11hUXMTnxUqNEzsY0EUz+3t/3hvY2cimyC8u2J+NUqjjejmSMLrGIcfeVD2Azb
O4PXBWNDaaM6/rg++zfHob4J3uoCOf1WnYS4t8yrMoNK95treMRFC4ap3JBOYtRQAGwkvbwPQAqE
jEdWytQY99ki0+7hxjdLsA8q+NDOWjKcQl+L38UwAd7p5fN8L/uD/N5OfjUBcOMvOvK1KzTb7gu/
p+aoLNcdTusCz9neE/BbkBuIXsvJZkOvD8rn2sc8izpzGtV+ncc2UXczA1nfEjonO4TjOAKnl6cf
dtsbgMGaXo624SCQLIMJYn5lVaJKGCgv15Fyg8G7YYLCUW92vprTalyMSYdx67R1NTHZG/5LLTkC
ILw6L7No9p5bQtYeCbE4BZgUUkkKOiiIAZ4owowhJ0Mpn4O/HcK/UOtq0k8IEfrIWVWI7YX7gohi
HvOBarOxtBoLi1JvmURndAW+esk1Bwa4JRKN1euRYOoJeWidoYwdRiKRR6VS8Ct6GH+4Dqx+6dOM
kEJ+HXwTNqom4HlyYJ/UT57Edma5S+awoloVsluTIer2nGyG2bq4WRn0JpVDuoyET0yHEbsnvKmk
DHIuuGP5C9mSC9k99Oac81sj8M0QXqu+L3KU1S1/HTUrdxXujXo6RJ3RKC7EHWrmlwTvkNlvSfIc
L9uPX3L8QTsDgrxuNCrRmxwC/wEwzlWg2O+C9uDWz2QZuEco4m7SdKwxuzPPMm+4VsvoHyM3Kck9
DR7DsBb6AfsQrXEyHaXEjpBYV13YU5lavfvf4u0Y1wFXSY1HT60Wm2R4rBCZ5m+AN2cdaenyQ6y/
N1IQjozZzPZLFhTTt6Hcpgv5Rj5PmHXveAPnPVEsTH4GDtt8e81Fu738J4JgYQhNX6nZtf1nH10P
2BYYqsLP3CEAAdLgPUXY1EB6wVufAjMlL2wBYJYf3Qtgbxzv8sQa2NaCIGKpBq64f6lx+FBwD0gR
yPQVjJTwUv2qoM4T98bjVfecfzfP95Jf8CaRhPbz6rlSHQG4PsIr1IO94qNV9SAlS9J3RsSZIETL
kqCz4MYzmeyP2eGqWgDDx/JPwCmEDkE5zlmvgRgYCZRiO4uISdpjeYsm+QAqxMIyWGyBESEdVCfR
P4FtevIomIsCSx73baOHmV8qC93eZcyOQbIVPA7lI9diitM70ZARFOZQKvO61PokGYX8vNIp1sq3
tZx1Q/lZiYxRS1OFUDlTXO0w6jQm1PumJaZcvCneOe9buQgOmoab8hSmTSyRHxGVR3RBhyiUuDQ6
E3EfkxJ5iPhWmny2uAeSidtv44jYgDecB/ar9fyDtpgmt4472HNDwBsgFY00UUENY/w8JQq9dBu0
pqlS6heh3p8u9rRklYYfG2LQdxiZDMLEADbZOWztSTXgFzVnGJd9tV7VQ5j8j6PLNnQodhG7BRbq
rZaqzScr5CN0xykIVQzLVnhmAnnMuET2T3hUs2x1ZXUpzXTzIWWPemIzScEg7kZQ8ttDtuQ0l3Gh
+xYLXOwShwTS/8cFcfAPOfzGSBRAVMry4RhwdIHqB5QL3tlv9XKM4IHHMxbwnKJPXuECwUWO/YJG
f3VdKEOZpjPSVVm2dlLhVqk87gc1L6y+B3sJKDL33C6UlJkeYDzY3semPm7fuD8iee/iqUorBGsq
Pr59S81hzexvJkxXCCwLcPU36HcDijUglQDgzB7L4MVxU2D+1L3r8sUA/cOuLXE0URJK4M4Ug6Ya
SjJqJbjhBaD27UakneMT5LBNPfcdMLzx8OvMXVck+LRX7gu63hnYt7rSRFpux5Vo9wRa0dpVJOks
N9v7CPKOldNqHmt7SpCrvr81jDEMq8spvr67oThuiPBZ362zKxQZpdxGS+kaQX49Q2MzMZ/b+70e
2v/8jLvwdgK0HcMRyR539rf7xJD0YRvY1zB6e4y1goQv6bbrLHUvoYHxpJuZ4ZQtYwRLwBtV9n/X
owHyy48gggrvCnb1N9Sf8h4CH86aHGNWL7viRzBmM7tKtF1oXfV9j1pH71LGNgxuW8yvq2H14dQD
4O8k/tU42n69n4x7cvFtmk/FPbvhvZ1kylubc3IRMA7kf/ciSDWz+v8GgX7C9C22Ws4LLjnqlSQe
fAUujVeBw87V8e4VJMlYPaMvGYain0NMOQobiu587tI0ST71ekks2h0INl6OmXv6IfQCpzJLKyXP
Lumn/fWLyifw4dldm6U2G2L27ekjwQ4OSKG/Fusyru3QTpDOjAgP2OjbOQLL0BpxP3P0mmDwuCmr
MtVNnbQaasqmiB976MI2qdvg7xOtJ4tJTdPKswEBBHUWbpfz19fwhGhzdfPiTCoxDbsIJe0IN46f
cNoVCd4Ln0D6qt3TuohrfChMyRYmt1Qv1fUvIpmoJ3eERUbln6eXG9yDKXcZulFiJjOKm6R+5XOJ
M1OhUp3KnKE7J+FTR+kjaAUIXIJrANRKdVGjI5UNGLi5Ro13NR1sWhoJm+4z8Yk9Vmq2BUVfN68h
UrF4lChljLFPQyItY4rru6TUEHlvl345Sh958CDFKZ1CAhtfC3KWlasGdIjbpQKiSLBoDigrJAga
YgYKp41tXAbCQugGkMwpS2Jpm6OeB/wrtAvR3AJNY4usCihnigKIVsPfQG+4jjitz4wbzy+UtlK1
liNk1/l+HTNDqBtsQvBTwKEMdHXBit0IgGgBaZq5suBRY6V7FvTHmp0mUQAka+lsBptHl+jaHcbU
Qz3QMJdsMRVBLY2MxmwvxQJHUnlHR7VtWNg3/iPjsLrsYypRnmNH/ZCXvs5RNWjEdA4dzPQN08vZ
0VlebYn40tCkev9qLR6FNayoCdR8hh8K4FoyNxAF0ZXs5Nu0N9g0P2k0fPrucnsmjFmESKaQ2fd/
kHIIBZPUe7NMWOQSfjRBfcUw2iJZFZIwLQBMoyqHtOzu0R5hb8RsHzSFdgaskwEfb2OSM/CJ0Vo6
QJxiVp0KbytbU1T+vn36lj+xIYJf6U8xkovThb2VdBlwCpp4Zk838O+iTZHD6IXhI7XbV075Az1v
3UphBFA+OcuZWkCi06elDJeOkeHsxo8izOg+rVxuE1zwnvM3rtxSssQuKlt4k1/Iey10ymnJXPQq
xw1LzJIMqXeKflVSCscIqhNR2myr+AWigmvOyl38fkaOOpFhWAVKq9wLzbMKDJKoqay52rElkmET
m7Plb+0IOLszTarUH9a7SptFhyNhREtJhyTqfp3sFPYdl+egB6OkjivNwO8d3V6fgdHQLv5AY837
2v1+Dy8bGXkFrKR5WqC7AflEWTfeg0sXEVrY3ZLOJQ28eKfjx+SOFW+45gzbzK6bWqXhtXcun17P
T3KSC1YK/Tcnxhg/XpJI2KDcnyOw6553E1nHr5sU3mBX5D38aMfYvvJuqrDb9vlevAfAo3JNlRyk
FmZZpRmt6fYtAMgFDiK7w9C6c2kTrbLCHvdGHgwJY3s/3FSe214AmPAZ/kc2lyrsBOEi5ia3d3ji
K/Fjb6aisSPG4jaeyd00wQeI1gP2Y3NFCwLy8HnlLVT/xT7oDZbamaRmsV59FEIj1A95UvOSPnmm
+SCStgFtXODMAbtFp8lChaxTAoHEr1Lc/issbl9WzXjHD1k7RXT43q9NP794DoZUwI6zCmefnMwG
kUKS/Q9HAVuoQza9iWoR7LJU/a0V9OBQuzav1mEx9tZYWRegGboz3oHA6AxPZ2PKI8gSmCvRDYrL
I4OGaAL8B9RZzCnUbBsge4+Z5GWbUN5YmAGtR1lUrrOSb1rysGY7ZSS++tBTOtsZEXi2Nca5ZCcn
GVuHyEcdnLgy1SzPZA7mShcCQqtUWDmK+n+y9UPGMJKDdBdf+ZRVq144BUMvz1YCe4nTeYdyCayE
BwwZawV3l5RfwpUOn7iKBOHh54rOlhtAEY1O1cUdD/RgV0h/Cpdgu0Dza+/ONm0ENdL6iXwB2NTz
bwyhyPkEWVAWMpwb7dqcPt5hn/65IfoOxgFj3pKavTUJNcyOda1yLW83zomLWQIN0EQPEhn2J5nn
FGoUDC6Bn3eBjLT7YzAEVfdQZB+ltKWwXYr+8r+ojlM7+RvSOgqjHPhLc2O1GbHO94yiaCsj9ezq
rEu5W1iXqTu1BW3/DhQC7Lkm9OMRRsUaXXBP4ElbYmKJcayF+n4riV0A8Kk1WWheF3X23auztAwT
J9uPMThg1JI0v39tHKadcRpmj59AY23xr3ScjI6TgfEcK9XnnQ28XbPcx4oV8JBQVp0a592apPJO
97el3tcxCffkKY2VwgBNDXKqhjbRLb2aKHSJsju3ViDLFA4RlCgd1eXXpeSSREoW/qvLDsNAYiAY
Ovj7uvv9biw5lHkgVRa/jww6QY84XyZFDqVR7rMbo/tzsfU9N+as/sOxWNAapREMYtbvZV3XRL1i
HhtiFGbgoySgt1LMXUpUkKFEN5TePDdkPICeaeWTWaIE12VBNZBbufJ+jrw0qrJBDdyX1MD4hLqb
FRjiDVtLtO7qNqdy3xxWd/rerLpvGKi38Ko/Xcv8AalXz1yyTs4lcNHn/TBrWD/NP27+7hRTeUhr
aueIIY9tXWFDAoyNvkv+ZE0ehU2n64ZQnCILPjF7ZShyxfqwnCdRWXK097FqJMSRSvrxbaxTIc1r
B0ufYDmPuy4jut+RDddSslVeVJJeBfbthyfq2ZoGLbuhXmEGeQfOM61CIBWa0Vv7hyEB/NoF0exM
JExke5xvV79e21GbppoUfA2bjqLK5nCD19b3IQy4XhhGNLuvRTa59M3XORRc89U9bp1xRt6UkLVZ
6WZkb/Acv7toVFAYBZtEiT3MoX+29XZNJmhJbN40JbrgdUb0gbcT05PEchcLCaKlfBffbTyhT55K
QtFy9fHdtgAOL9Y+sKKGgHR2jSueIWf3Z3znEWY7SYL1A8YZeFc9uir7I2YolZcZDrF14k4oeBUW
T5XGsQD2CTKEHSwgTPcuOEibAXV3F36JQHdUMKgxdGVf99UI0Sfr3loerdCog8yTR6EiX8i2fiLq
CN018HJdfMKensUbRHJow8yrFNYAbXxE3Nt0Q4AqDHybURKnO97BXAehEN65xEgXJunRdVgQ1RbV
S2O8WfajkRKKh502fVfqZJj+98X9MJw0j6F9q7gKU2OONL3VkjJINBTBNg/MKfqBOsxcce0CXcrl
ncS5ncrrBCfJmh5SAi1Oa/Ma28yaAalxctZqVOL81v1G3iSuCWndaYTzId8+cADiFpK4DvcpVFjS
AkGPJ+9IwBEHcurCk+y/AHJ/oAdxWxn7QMeq/pBxIDh9TScjarJ6Bx83iwS87tJH2K82J03TQYfm
cenT6iAdIS+Vvqwl2aELiSciZwccIsxlUWWTIvcX/+SBS/KMNaUyfq1eIImyhJQ202BSdm9MDCdR
pCxTv+5Xq3dLrfM97W7rzxfWLjGawSlhYH+VfBAsjFlF+LiFClRTgAEyZRYE6zT/+fQap7b/ThDz
zil/UP7fpPqyrvkWWGMasSL0/c+B2uaeMsH+2+s/N9syOxct+ZDmnB2CZvJi2sAGHNnb90quLYUt
UoYiLGMFwp4OxYWmX5c+/JhWdD7ZjFAEb3/9XNIWLqooZ+ZGO/TCJodcSfo+Cz52aUqFg/x1RS1W
OAlj0hs7vYDmFq8iSRUpKL72dSZN6WYr3FsrcPRFtE00pVJIMJ35s+7YQY6I1/i1mlImiIKaFn5r
frL3T+ZzK53weciUUg20LnvLcYhT7IAhxxNz/SW7QUU2Cb+iDDIV2Yo4yvi78QU+pCtzM7tju7AA
ksvLRCRIFhNyiToCSPCAaYkTfk5w8G2v4hGw2d25KNVEWcEvGNJfQ1p0jG6VgnUDazP4i8MuBbvN
T8Jt+KOseLQURvIzlJReMUgsORjAtFg5fhUgQnBZCJBQABTgiT18gt+R/44DB5Jgmb6melgyTgUy
dtrSCYQrLcebSl6Jw/aPZCKgFATNNNCdxuyfUNTJtnnKOoa/qYoqgGcfsy7r3goqBwlY4EOcGv3y
x5Kw1m4z5lYZINIWhy6sEsuOXZYl53x2dpT3l20U7IAHi479ha5unqbeykkCPC3R1J/3XHcsDoPA
g/1w7sxFDKQfBALkh6xa2/ROVpmw0LQSi8bZMqchuVWdsHBscWqCSs2R5F4leIS3qAeikRE2cmZW
WUg+ntBPfuKvczTQ9z97/jk8lp3g2cR8GMZg1njecqpY/oGhBcW7W7tqo5OJE0Oht60e2CFwymOZ
B5eu1P21cqYZpoA5eQ+wUsrpZwHUHNlcjnkKZWHd/dLulOl5b76pNc9ihrxRql92NwV1AAwCKelp
99Rhs0i6JhQ/n2rI7i5uVf50N/CWU5WTGFEleu/yvpkLszrWz3CqttOz5TzgnFdCw6pzwFp2Rtyi
yrClou746rqJ7gWeciu6Za6PHdB37aQp7wTE2LDjjb7jQ4kVgH0JaUnurQ1V5NlSWVLLQOpRyGMN
DK1mSDEyBGcl8rVYzwFD3e44zqfwIpmGjTqsr52ptl/nKQ0EhkbNPBwatUxrt0WnL9VbzojsRXfE
XdAitl/YXb3alVDNDnWyv3BT/eSaEpld9Vb1J1DPNe1QO8mx9pNfgJt19gju6UH3kirfwcH4j+P+
tmv/gY0uvxh2NfWsNMMWL8UCUk3z6+liowD0lXDwHte6n7lEnbDPIWaZMSyEDwsConSd33aeFjSZ
hsUKpbdYmqZku9Ob1gzt2kb1oqRyLo443EJLkgdpMWYs/h8GHc6W6+I1/mOUAV8wfRFjp+28SB/k
EjTjdI9/1uvHVeyckh1k1dCBd/a4B7p0nMD8GqaYtIij0mzwIxFnsUQVvF/crRvw/9hYR/MRPmKs
ryq5yhRnSdQS6RLqrrZ6T971lLTYnoyRW5eazgzOrt+kZK4rmhHc/+uGYVNdpFld0Gg9r71a7MSZ
WP97Zvg5Iuy2HTutx1+otOsAWhTXkUfhjhHywh0lqHpa5GGQ5MwdTvQR2HiYvzWyThWRe1jNMyyK
GAvaTIynObTG11OI1egBiMRXtIuVA+Rb1H+H+3uzWiknJuNm3XBu08/aprSEypFhD8IG9isPcAG2
SbStWYkfxbTtJOu+K4xhwRfQovx2kK9j0P5YvA6wkE72b1Ou7xKY1vwhnx2/ExYQsNqRna2NQpH8
LuPyVUsC5DMJzKVcgH3OZ41UX4EvKE8dQNtpHoJM0Q0qrPQLbqValk1afB+Z4LpB5ftIjjZk3l9p
RXhIr1l+ORAkhNc5NTGwB+m05OMwnfzk+cmh4bsUHCvBw2N1efL0ZuI7ZGF5jjC/CWXjH4nSqPa4
Oth5vTj5tfRndrRh8Ysi/192n0W9VdSE1c4RNkeFDuJ2clWMCS/+Cx2Z0VB0s5ltNjgx8FcMYm7s
9WMccaKs7RX/gxqY7o/VB52haUFTxey9ZN/IFJyNa/o3lJy3ofHJjk9E/BBZeIesEPSSWjYEZvW4
jS95GkVpFaqlbcFaGBm10WWQNAWcepTQWK41NCGk+cM/HrwJhe2ZiXDWLBLsF7iVSJ5pgesxh5xW
frSexwCRzkH5CSORPHcRsiYxc50ERA5hcYh5i3ecpeI7hCj4bZAPEkVTD/56X3G2/I849HWBS51r
ex4aHqwI3uar78ghh4MIP8gA5ispShl+i8ailwQLURioUUKw34JHZQsXClQPcKnEcjyFA7SCSrG+
D69t2qGElZ+rUYNgK2y68j9UDEyLQV9PwAlSLa7V5pH6Zjy0alPFg/F98gcjiWh7w/dFVq5vBq5s
cUI7253tS6kACGDJ734DpAPJ+3yU3m1ryrkSWe0SL5E4ZMbHgmHdjqZjUspMYSxzTs+4GEfZ4C3H
lwd4aOiJ1aml7R/j8+IASLebQg6w4IxDmbn/ZD3Sf3kyKblwamsr1YQguAALipD9LRuHRrOqNKvd
CuIyv5VdYznJr2Z1nIrXbyRPGk1U8iXN2pJKnahoRUx4OCyYzE+6IC0cmNIFQgy8ls+Dxvoyr6BA
IIh+J+DK/xmXua4OqpUjCNoi8pzdOestu4/7AhLkOMmBuzO6x3AB/fc51FmySN8bfK06czqeLIwg
fXDvaxk8GQW13ysC7PIBGh7EZVY7CpmqZi8S/8NYOFl46OnyzckD9X2ESdnmobZsew6xdJHBVGbq
Mt2zEdjdSCA1cftucNjPom/wd8BukMtCvU0T2nlw8KYAf0H2cAr0I2pvxfkuVrH8yyUMT7o4fJ1w
sgb/gtEbQKSs6nFlu5lWssjByqkK1IaD3NWoE5EC65gI13jGa4/U9b1mh84YDG3rlED6TJAv9V/b
moZ8A4YyBQbQjOD+K3hyC4QieAnW8nKqQFd9CJ1vrPoq51bIZIZEkSM8Mj9oPwr91wEatiddSN31
EpilAInBbaUTwSDmgWM+tX511NO9MEQZ/L5J013uJT9YRxP6bHeWD0X2eDNSXNoU/ekXfDoV9Deu
rSxgzV267WfQan1wTCg4F9BYtTCTof3/wp3VehyRuPSuI375GekBYGaco0J7elZ7CiO3/6YTYg+W
5rZ+spP4tQiq1nhkVmB2uxXSxYV2p3brjiPQbLVhjwralce30UfW1TIUj0zbZ0PEgViPMjQQ4luS
0eZ1GJSvUhFQjjwX46dGloaU7bblyi10+QNPGjTiOA/7BnnEKKqOHmHyffXnNzMR9nt95PYGYH71
ZD6O/Ik6WXekT6EI552FnQ8Y1HzFGeyysnTqcyPAo97f5/y9zaFiCgJMnHCkWUKpkcpj+CZsZQBW
tTl+1AYPN0gdh1d1RS3YLb+IvRbv2Qr3DeD1BYyTtNf31SyWS+nEucKKGiyzJdNcuIL8ILuwTmpw
lw2pLJrJoVxEGczDZ+9EKaPAQsG/B9sfygX3+Fzx5sqbjbvM1v5oCj2ebU/83QIerCTU6MFIeqac
9o2fJbwutwMZ8tQX3a+SwZKFEK+Ue6WV8rBqcomc/uiIpMaELfdqudl10zYnCcEeLx0tT9Bt52qY
xqUbSTK1MvnBxpChtK+bNQtwFr3wzjCXb3R06NotpGK8xJYhwyjKh/HuExSm8g7vrOOtO/BZjMiR
etZCJ2eHhFGijpAlRYd2f++JWuBPvRNwTSTReqVbPAYxn7JdcPHpWRg3YaLurSuKhXWR0lmWRNp7
/W+Z+9g0iZjyFhcyy14McO/qy6Gmux3o4rNDlO65skquIhxPCqYG/6YdbJ99Otxod+oUxhzVt+t7
Hyd0DO/NG8NjtCk5K4w9xOqvOrk7Pl8QQJmUG26/kOCex7r0FZhe+yAvLgERrj8V30ydON37SUSV
sMTDhEVExsJc5jqkKFudVi1xYEUvQW1xCOZ8z2nbzByBaKsC9nYBV4u0G3j6Y4uaTHVPDaRhJ3ZV
DLGqLVgD0kknPGi0mrzi5dg0VIpK+mY9nr/ofWFbYJ3/vqpKpSeKEA5Zs6LFbtV42ljMk2RatCDs
T0Xx2AbZc4bITX8Od8I/jZ8Hknz0aNMvaNQ7WxX3arAQDlvMIO+ONT32m7yLwoEqMETx4Bp7XIsI
3AmoRpFhho82+e+5odicvJ2dTMt8+NnViwgth6OhuykEOjx4hLwkK2wFiwT9I+zJBGxv/4Zv4vtP
7DesGVlnur+19awLpwKK1+dtWQceSWjOnLDlNamIbIdM3iEqZSOycOgvCs78xKx/ZqVYe0HqNYvC
9b8186ciZjq8MNvoq2cUzLtwe6jcZr6KtiRM6ivflrJgeOrLq24IgAEUYlcvQTeuKWkDwx32AfCw
quk8bKvva9Lw2hjPJ9UjydkFMIdQSCyKbHK13PckwZUVC5Jmu7+JX+lCruIkOZtjPfLp2MnUd0BN
PFXj3gqoQKC5CVpU6OhVXCbYvsXLmAMQWE0C5dvrLlxu5jbQmsl03NE6i8h7fr10z9sLesqMNi4N
E9Rjk7VNkpJqhAEb2TGd/fqHYiVBjgiIwI5ulWt2eFtq9KSS0+OV1PeNgf6zyz+wikTi1XX5fOBa
PZIubbrB3fLCQaAwB9M26I2zfY367MKAE3i+Ox6JT5pUPprQILpi6gSRB76j8pz2vi7BzdAJPnSe
uDZVB2k/gJ8uJKURel48EwMGPstsBFjgwZ4IZb75UzN/oaTcEnnal+79IhRqL8C3C4wxFbxEd58L
CzEqyJoZgFtgjjEMu9wkDl76eWLafc+tQs47jZL8jPRhlVdkF0Q1XU38vOIOSZ45t478yEGHvg1a
QlVFf5KLpXQYT9TcnerrRrZJwFQ5mYBqpJ8EmZmN2G5BrAx7UFiiDN5JBvl9ZrDXGVKDLCRn+D8S
nALhyL07Gko7sPmxxA2LfKwjHXP87B093iZsFijA8ijiXRPjmQmNPcwztQsOGt0G0atR5Vr2Wx2R
cjrerDT5bI9Mxygg8/TgUJQ3brlcreAsJGOMcg0xIC3/0vyLu9AZPzkJgK5c7a85tSlvzTIGXDEp
r5gNhulpXzEbBIadowVXqreH5dkORuJ03l52aqQpbnsuLWEqO4+PQ+wkNiqF3VIUoKwN/0F6TiLt
3/HCHK8bnz8YA0nr+QtEVepx099SPfsIGaS+rHKUirj6K/Fx5LlIZuu3ftBmR4wsg6XBD1pn8Vxm
LotZ1oi1aSPM1PKa41Hvo3IMJv+kPL7MYBoQc3B/j3Jn9cLU0AuPJLG1nivGeIzPBbs7+g42F164
NYkq3ekP9zQOeJn2PIQNssfzjyu+F9Jz+2D8M0H0+59qpkBb614nf+9NAOghXbpT7l0SIwWdVzsr
G69wjxHyatfrf3ufewNC3Fwzk1j5bQmWvMSRS9XMUW3DdyW/yNWsNXckHaNXTZ97iRbfOm96KKxt
JbYhGGoSWQvaQ1UGJrj30qx2hONTYGvZ/o1xcLtBc/F07jqZkyq8r7cayTc1J8KZlFBcYipLJrtW
WDxxOv+K7AR0/GPygYNrv1sUDynPO64Hf4IXH4ofJoB8Ps3fIrLbsHtl+yps+1DSagsQcZaJnTvs
Me8AseIJJ2JdImbSGcQ621JjxSekdS1O198fn84BKBXT/h/f3ptkogzYUDYxGclWe6HLaMKFXmxS
FKlRSH1MeliZAoXC1M8X2/IwB4KdsR5xgaI1srSLt8GjohMMfICXLy+zgUib3THkO4qSoDZXBkoF
n7ZzddpiDLHhfVdLn3hMt9bhHMC4Rfj7VNKjF/pInMg6guvEK9IZchG1iur9tLWfHjeWs5eierNr
QISYrMiBpmOUO5J97p4V2tq1OzWKsvtBH0g6je4gzwoWmGwJqaepUbAb79arWd71VM+B0ypNm94k
tz/5AE7UIxuy3z8rU3YsaJjEgtklmxZlZmvV4udcRzh42RGXq+c7KmhSIO0nfgFjVHHKgEL/oRa1
nj9uYM1fBXU03n9nTZ/KHRPJ6SnfeyKqIp3tXAjv+K8eVV6vgkTp5qL5Clv/tXAMecMQf9RvlcsS
50NcEnw84IHUTO9FcpNXuTAq+H92sEDQT2OnUgIpL6LANAayehXPTUZ1PwhFg5MR59w7XIpHv9FW
T3nJA3O1Ynw5J6Ef+bUbRJraVAaO8f24pcU63QWYrgvRkZV41Hlc6CnTByJ/o90YS/ofBhmQyhS1
vLF6/pexcrDQ6nZsl8gO0aUt16MqeFLwTdBufoN62BqgupoJHV773IdX6/Nd9uaScgyPn5XOdtf1
n1emBly1rojYkj2mIW6L0oTa4GclB5OeuoPRXAUURti9CTW+hDTW88KAWB9C45QHd4fT27iyDQAa
+5IN9SD69CN/STjy+AwrHtImNGFF8qAofLATjHdIOwKJj1ZKit1Z+8kTZWWMgW+XdT3B9qLJ13JC
L71BbfYHMtGfpQ+yiunZToCT7ohTGWIwXX+bd3BXWcChE+0B3R7XA1ZMzKoL7/VMRQjUzdwKZsBC
+LUfuMRCn9qXSwJise0LNeuJmCDZ8zIWi6s8ptqrXJui+nmE8IveLtWy7Mk6N2mr01KqHGKfBwOD
4vvD2lJIN1fJX1uHhz4kjF048pYlqpP9faYifd9nt9+WQq3cVBlql5q8fgJQ34rDwlpJfNLxm2MN
1GKgF1H1N1IONebnV3N+C8ol+lZv9kFR97UrO8s0v0V5qaw3VxRQ6+/393E8/JgIQ04Trt4LfsoB
tjsFB9ZMkyKMa2U1bIqXgbssfU0T4Yv9/s7hmWVdBWGHU0qEg4mC9ctnepfjyp72Qa2eYNFS9adp
PZ55nUOIHHN4ViB6XnH6SBFJVnre6Qrc5+7w9b4hRvwDmlKNrt6Z9umdQJp6Eyn5XNVv39qiZKL4
R+wOQVm3LUJLtten60pjQJKep7O4cydetvcaZRtMNfvyYHguqm3vKO1WwwP2ynLSq1epktHOQUXN
5ikLFWO/rj3NeNW/PdMHCvzmnEJ+mXf+/oHjGWMU8pgk04xnZFixaJ8Oih8qymZC9hq/+P3Dmn17
Ebnbqvnk9896gdu0AYIwGY4M2qp/m4m+adwU+GYQ7dy8WV18gRo7Vz2ND+AhfGYPriu6EBocYnT5
wkV7qbz+lK5LYUIBUKGtAnN9BNLgGNbTWqIUqTVjBLPEm1H8eC+ujieZsmb/6cut2KOjYoigDRuY
QgKfx1Ny4xt1R7BbCcgLpo6+Ku2QlXMuHxCK9cGmzcrI8KHNbdPps284qxXoAM0Q+tFv0a90+Ca7
EUBPo9SdwPkXUx0kusGrOSmC9E0qN+Tv1uC9Gy92SAGl2fyfWbnt7qPmBe6J1JvHre3Xw+cRJw53
rfF0vLOqOO8RwmJOZC+CGjvGwJbHZ+HzaYXw3CgdHeoyY38l0A20jh9KxUmEu5qQa3cuC6EfYkGe
QFXnGru9ZpGHYKaEuvKexb3gbSDlex/Iw+mET/d0GS9Isp9fnuxFwqF0cKlOcXyFL7nr/PlOhwGm
nrafnJh8KaQv8HvbNnaA17k876PjxdYsBoFgYm25yM6LsRxImoETT1wx5IzejbkpSf7x2ZE0rJWi
tWdAzvvzmVQy0sxadNbAHex1lCfGLFE91uhGCMaWAPqQ2nOgQRaPYPueXP8MHmCV5pTQmhbxc8s1
wNsQd9zt1Jx/OeMBMisjGMgrdeWygphOARp7Z44k2T4jJYQWi5okB9+a3FTRiEsb9RuGZ4fVUel7
7qJnxLlrxcEfGkEsP+E0jZWt12559gp20dSmsJdWdM2tROMiM2tVA1Plz1n/+sqYYU+nz7QccKaj
hR+JbIddQygFoKu1fi7gdN5GzOr449Dv47qTGRZtHENNW6Lur/WYPZyG0ZUD6lxg6mFdm2WLTVyR
8BMoGa7pbfZfjOfNs989Iii2azX7Q39aZwecooOCa1Zg3KgkheFjIu4BTVErfGLdlz1NJwOYA6vZ
66Fy038roSU3s4O6367mYaGjcSHTGwL4RKHUdg5KFsBCR8v1zpCvAgMu1RmFqP72oEJvSbCDtOEq
jLjy/PHtG1stRHbd0kHr8l2qJaAWDuJDWff5pqnGH0TihHMGjXY6kWMyAeTwpqH2zk4JxwodStq+
WpjBINHBwq5c1S3ax/r3lrHFPqgQZPHNPtGIXFUOyG5T2MbtnJ5s4FLMZpai0R+N19JnUarBwhwi
bLx+fZcZWN+Y18alpvsF3msOnf4GEAMSuI7pSPmngAzWgTf1bgYA0VLGl4RdmoZi/RQv3uKZYirq
XVLPsvqse/qxqcCwgS6r2dJib460mEUw+zWhtFwYSs86P31fEyaD9EimBUs7+a1NT2F9lNlR/k/a
WVFEHcSzvaUc6L/+nxxu4NRsqhTspxATbohncht2Rixe657r9SQEOCpMHn0SzqceyJFNmH1N6b7u
mkhLt+22iFEnNqr6Ezhj6uJpuKZCc7StvpXqFy4tAUlaF5b/O/Iyjdy3ZrRYYf7FmzCS1N93xLki
WSgAxzZOW7TJpvYi+oE1T0E00g4UGMubMbWB7ZpEFnGkdQAt9qGCVPwdyF8oUEYmTVBZLtS6411V
SlLeatu58xR9KVM4tBeXZmN1bj5Cx/NmV4d+vT4hO98g8EcJtoS4U41EnY4t4Xza2shzFaAbOhr4
DlKjCGBzpt0O3+b+oyHWaVhIGvPCHn872YIA+IegCIJ3nMfvDJtE3KyogBf0JJiAOXYcfq+GJZqj
Dk43a+FqJoZYPePO42wWsCZiFkytH8ycq/Kd1nObKSEcueh/XMZZxmtHttLnkOd8YahEpRCdlJB9
sqsiDkakjKOMEU+wJ0K1tbtHwV+qPq4lC3kZmpmgFmNSDluI8ILOkMkBrhzl9PO3/PYI+UJr94n6
0RKBqIaJQ1hCE93G9u+/j8Muau4IMnrM3TdJMaZRf0JlYy/wmIkPAvEtrP4150Qp3UPOvDDJNV7F
OJuFiIBlhZSg5jkHzX/VfJljfXJRtiFioSj2CmdtJQfKpXA5cqLYi1j3er7Tbf0kXihL2jC7q/zh
ncwfrcimRlJX2+P0NIyx+iwJYuOeejNOogDXjfAmzW2qceKHu19yXOyWqgPpVGlWTuYnUpCIzZAO
iqEfNCQBlpQqEXuhQwFSCi/EwpmrCfft4L66QcLatwQwZgM6llAqKTR9Uc2IVV1/xCO+JRuKRfp6
bHIMrYyuBEmRDr/W5sqMBNXDvmvyfn8JFA+7iGVRWYVunOOLM9viFQa2XWX2JymO4Rp0LRZjKNlV
0Xf0uLQnUTdXctvVoX4zTF+5wqAeRxQJYwbrgGc3a5a4XH42LtiX8psYLKhp0FHTyFlH/Nxp/YFA
plTwnHZowWJURy5BLGoqjoPnD1WjaKTtIm6uMXs/pcdi2+rRwxFl+2DcFHG5WA33m5ViJcTtU811
RsoimY5q1Y3WIvjrc2hbiQw8xUNb7iBPsrvYxgYnfuDPk76YrzbOt7XgvEYg9lToViSS50QrU84l
6o0t5BGZuc5I472I3Z34JEE30ycHL6/sW9OkGAdgrpOwGfup1FMcWEkQM7fOCRLg5iqohXbXd2ct
u7qSfagIHGbVXePngQl9TOAZ4DpFKiDTi47Xg66VwAHuD/4R/f6ta6aF3Gz7e7tTrRc4G/KXyj2z
LYZ45EmZrvO8GOtMMrfY95l9GLWL0QBwTu0INea5xnjYknRfEAAVJPihMeJQVyNgZAYI3O4SJ4w2
kD3XJxXWMQwkHSxXOxytSqkmO1G1VXVst/rvfr9qJKHN6vNExXlBmvh+qLflNEwXA9DryrQZiQbM
K+fo8YdtDawGaPpooglPjVJ4lOhJKX6Z23rd/D9LYDLmHvzMuI+Un9HtK8qtZlyjzIrMTvgBIvqF
goiWfAqrKPsQz+r3UO4X8V7PdDMIjeqKlrqsXRwqesOFE99oz6PEQJMKZWRI5+PVPnjjpIYOxCle
AHECaE4ygvi90Jly/L9nGtGh7qWJW8eKZvdZ/MzUxpyHETAAZ8GZBZt+xogLILjrhW9G+wfhVU8X
C/pHdd4zmBuxTtJn4H6Y4l5wM35U877ytUtCxoYdwlOFrxFzpFVI1zV89AneL00Ekzll+zt+viyy
5q4Adj6tfDoLVr/JEL45vp2SFQ1BaA4kXW07Aq+joDDgJQFWqdgSbWb9lau0n+feiCzlF+JPSN/A
9VvpNlZPcxZmwlyjJCZPMi8FOb51Jq7i2SdGPpd+2/aLov5D00x7HH3DWOldtjzaEjS8JzTI6d+l
PLA3wBnYX3il8wyfpuDboPe9Zqj0EpiLahcJdoxQLSMvojvJ/+5C5lWwiC+YlEdj4QlvbCtP9br0
fStoCyeLPb//PFCWJ3QKmOXPfP8qhVijCrX30KxR8LX5jpCOsNPvpuS0+4FO+j+BzqeGRe4Jezzd
1kERnEKUB/8NWJccBBhWDWF7FvmFREkj+RXy1BrHdveJBCBKSbqk0v9q8DptbnW8Jrle2V9Z9j1C
p9DqAd7FQyj7PyXv8z23OudrqlRiDkUZs4wnPLWDMsZGS76atlw9Lkc9v3tBZc9QY0rRhUbuRY/c
jNnCBQ3PW5579jzAThpUeJ8wZRd5qJxcEoHNa0UQ8jGNNO6TNYUO4oYUlg47927HzinC73sEPpw1
ZKEjpMRV4fOKY+zZGKgDIpAemBcDaA/FpTxDt1zS3D6OHK3JnFjECyXxuWWAj7QheCdTabIUnris
mz0+bLzMqq4kawUBJ74cZ+lSRC9OsxMqMguvPMdkosPWaESB612uap+VgJLEd9ToW+GW53YNw8GV
aaoX2sMkkR4X7THls8K/j5xStfE/KO6Rwq3tyvlU6WIXRC6I36urb9aMkXCFIKCtSadJC0eoPh3V
r2NWUTSWrhVgM/njZIuMcilk8snNQJI04x4gbqfuwcPibBXJwP5lVDyHAY/dXG0F1lps3DWdVEY3
+kVlvDp4jjcmouh/SmF2rTGC1TVlIB/LQngyZLCVi5fE/BGvWN8KR6t0EON09oHHpaKs+cJ6ykCJ
MH99GKP3kxsCPPwzKGw76wXECSAvhkfeGU87MhSjtWA7gDt82FtpXC/vMtuq9jpv1nFDywE/L+5z
WmHLGEt2X60WhPtUq2Pp7QlDzMnnMjqhFPMJc3D8zIWxIHAv2mTa+2Za0fE1k02/c2mEkbAEuSK7
Mul1RLGByZj7yB36Oyf6X0J+7AQU6/S67dwp7fruZ9GPBTsT8utM2+HcdX7MlJnfRPFWdLf0/4e+
juzxQRKPKwg+fqoq3mZR/pcFDfrOOkmxNhm1qDgprbrowXLHVTt7IBa0MJfVLRjU3itx5DErzx5o
XLFokTL/zAKvM2lAErNDw1gRb5GkkITseefMgnmzzFY4uLdv7S5Ul//MrtIZgUbKomlNLgFsdPQa
lVaIPA1AhjKm7P7Y9aouciKIQRZtcR9m2O2MNWa13ALU6bErYEG4HmFU1mgKv+PFEwtkIPfw3wP1
EihNDzYEwLJ4Gp1XWs+nlnJ9E0QFVjCXbChTTC89YklHclc4eXaYrjHibE9f67fvImkQj1r0Z0r7
kLqGms6xNpdYiHnIc3bokTk+oWNfvNBvslofRbli8C0COm4Sq6yaF91EKOu1bgY9WZxtjbDBZgCT
NC/6bhSBKmHP9NXHTR8r8PqV9mVn1uRHWQa0n6PT7zxs45N08eQavmY0+6mInAcrzV89ueqnfAqx
vslai0e6nYXcfZZwTq9VoOAF4KrI6a0P2tyLjjuUB7b6l4WzDMhRTFTY3dTXcKqcu6tq31YHqdwO
KA5R4gXm7ZoJGPlcrkvrU8KDXw5khqSCSQ5V+w1FPKaJUwVDQAQvQ3qvxM+nkntTV+K1VFXjxShB
y1bJycx/643FgURb3bYMx37VYuzKwVa+Ma35Q6sjbVsK3JGlnpbhzpUUV0L6UTZ5HCI9yo8BkVe0
2kOL2sNRsqbm6SrGRBOB17sFosEiXc9d71Qe/EsDAKuQRzsT8LSKSgztmxHMIbHalNuuoGnV6IXh
sBR2dNDueB6vVMjyGVr5WIl0211SwUD4FUQuGOnhH0TTB7beqMX2Gl0EPz8gyrLM3iUjFo1Y3I2F
cMKknNpm9mRG8qc/k13Mk3p19L2prWue1iwucendyFaLy2R5NRrUDWvpu6H8H77rEuCwiHtnXavU
Rfb5WaqVJTSY2vc3P3LOEyIHUD4ukj2c3vnh1z0PwY9Dprg4i/0u5QaTHpYCbQOMJXctvi47CtcE
OkaJcAIt+v1u+b4Z87ed/puXH4Z9IkY5toXoqRU72qxzVPGJWDnkyiq3cOMz2jbxAtTUXDF8TFG8
bI2TkqZHk0R6Mus0qG+0rcOCoDEX6M+H+5RmF7gK16+OWKLm4WdG5ZwMUC+IfdRm+3Cr3MngjdmO
dnkdAdS85fsNxi8K8/Kda8Ctn7I44sXJ+GFsYwjCPDGIGwaSEhLWgcLXvguqdW/K6M+qsm7Dnf4v
s0ALlm6N+aM0nzlUseBe/x3alDEJxyFpV2CPjE80WCKTDgzl64KbLVNc72bvkHMYTDHlKg4ywNxb
SwFDe4EiFbZ1RArX/1mk7r/Pb+ED+CPbe37p3dUHgiSHZDDzmKgvN/IK9a2aYvyEkRec8aaoof1g
Pj+nAT1vw25/fQKsSmxqNe5CTXWLtSU+K0aZao4xftSPqEVrZGuyzA26baf9qcrzCTtbllcZfzpG
9yZWeFUXkRrgmWvRV+9gWl9anE5C88Mv85XbSPL+GYWbAAyJ9HCQxnH+loAlY7vPIong7bvTZMyH
YNeBXBEdzzLVdy55e26hF7aNuAOGypyGrHJfNr6g7olYxTncCYoRnOXjhqN35kddiwNUeDb+3QCP
GMtkciha8HUBiR0Gr6hoyFzrqEPifVYiznWpdb+Yzk0LpCmK70kxBflLnhmH1jdqmprX8xJn9I9i
ZOyHvtPkOuZfJ/+In3itdqvZAgELZVDUnlRjd4G7qd9JEVKsSDm5MmEsskBFLVOtbzy3apg3JK8I
4wfGmnuDhxORKM93S1peG2Fp3phWBG/ktEvXOTJO/peVigGsjkCFuH2BVo1VEV6yPvuNPvUq1P9h
nb3uBepLp8HdJ47st2NM9aEKTdoQAe4LCL/qanc1+1jXDzktTZVI6HfWtBEWpKPH2NE12qaTm2Tt
5YKoASXW2+pSVE5nQuAnVKVK7dlSOQ/Q7Ld1fFlCP6JeKkuOzIrHktloPbwnokFVGDpgfnrv0kSd
KFp+LrE6FTyrd2ofSkFLWy8qskZki2jSdxZVUiXlyyishZUWxJi4n07UtwOX+z93FxhjNoJdl22L
ekQrRxik+TH8k2wDL+mpOir7WeG4ZHvyUqyKMq1hoEBnpVDIvKyuwvmGvHRF8biOxo896MDPAfRq
0m9EcX95vua8ZOZ88/bYuP91Yqxtoe6E+F8YLjWYCFWzbIdQ1hBX8ELW994e8yFAcjyZHvwkmGPt
gQeIQxYmXkQ4ItnAlrYftHO0ZIA3g78K7SlkY4O/UhMSgbCQwbXkVAxsibT7sWn9o6tjZ+BVDWqn
YMAx4JZiVAgHa6XsK0zVep3Z9Iid5E+TEkER5iyChJWrpGoatYo8dzrYDRoyqjIfu7op/Fl/WjUk
x0RvK4LCNy/kEVkdP/AO35l69aFjU0x0ricYTozVtFktU+cCm/9FuEy83yy3VUlfK9DQhaOySdn9
JWCrfIeViBDiV6weZ9GSq4U2ZTutZYDw5aBheppIs/4sciXMBNtbDlDBEDsQBY//xTLD/dQ8UfzD
ZtB8aj3VSFI9bKNdyzCIE8y98Zl9pqNLXX8R+E9L7IrDqz0pw72VJb6ZSH3ZPJ/KSiUWWF+7PaPd
msodUOepkSQyqKFKENNe8l2jU7tDpUbDqhRNpiuqHKl8xtjvQUdxQCU5z7JVghGM4iuXCqDtXwdh
e4rPb3PsBfRIEwkqyYLkCPwf1/B46zVQ1txDLT6l9fK4kgPGsjHJahoEGjkDfga1iAb2oeP1wbL7
kkbtEgfZ4gCSy0Nki+AZ0TGBE1GMbVLJWUzdoiWBRI6KJhhAi6O9oqgd0xra4IXDAjhYbrdMxIA/
IZUzxBPklql8xonMuCz2k8AHyMYSvUloHNJMylTRngE/9skxSXKtEF9SLoiSUS44xtHuqSPmdWZZ
n64CmS3imE8cCunGATY3/1q8U/uWnatgblD25Zl7rS8JssFNW4magkJdMnHtHa68819fPp21KWON
UQh+ELZpaKNECr6Xeyk0Ht+ax5bOQ6LlyFgwzk1oQfp5is/tiuNGUl23GQkxOH6MvzLOCqYb0qt+
8uidmGTSBTdQpuqwyIFe3zZyPZsrZRKk4ILTQsw4poBDD/LISo67KXv+n/R/W7ZT3vTc0MTsezKe
exs2xIjCIm/QfMNl6H/nHz1McyEqURx6+VmXdD5mgby9Mo+meUKSl8P/msDJt9jz62TQcgxkLKDY
vvoyfc1YBq9jHJG0AF1DBhtAS3BB96gUqfUEJM/cBzMfFzWKP2Eputzh/llQ3hPfIvHUADsrWLhN
K0qw/cbnTtkA9wRNMxIazIy5Ah5wfN2YCmCnO+YDHkis4KEj/pZWy5iD/iJdeP5gnjCuk9FRHHBU
VbPJqA612qZWu9WsTtpIoh1kUBHP4JQUrMnb0o3rigtJvBVbW8k7rPFcvoT73OknDKY5ExepFG0s
oRerEJt9H3u/nWJeqe799S+QPCKhsjXQrTm9ohHA53WbYGKrwHAAcFd9J6V4TvMkq4T2VPficCXR
OYBQs/rH0nt6cZTsVOC3nFAQLGruPBC9FofrZpu6ohNEg9XqQkAQjuIF+AItw7iAGSA+ni+SXqvo
0TKDt2ZWtOwIecSQPM+GHR8hqmxBb0HVoHNs/jOUJn45EgoeOIycQEwPj9kG81sSpSAHZzAXH5Ni
82L8vBpYWj3PwLuLiWkKw86RgBCiHfhzyz8dX3NH1Kx7DcQzve999vqF0X9kFxSbXU+4qClm0bOo
I1kM4PoFSQJBsIYn5N7mq80r7z7/gqMrGacsXPgxfTPaerabh7jCnKHaTcNmyQwL+aByhdcX9NbD
BbjOSHg23ofmRLgh3NUiiDcaeFcfbOLgTx6wdN9Z8BVCvKMSYhvDYVdkK36q4YfqcF9Q6zD74+hI
jOdSfqPu3nobFg2LfifqIOKtNZ3Z3pzbAP5hxm+XkdKhD0hProYsTspP2JJIN1pLHvpGJp9d7tgb
RTprOI9t4mTakOOJl8LTuTqKajGdLZXuUhOq9zE3htZlq83ROj1xFqWJB8y6yqfcAWGtscOK1VCt
pj8vVpsHXdVqeCgdi97wJ8/EsR06vLx0iGUOVnAZ7q43ODOqZAdBrLrNiS5Q2j5flRyJkXzXVebA
ewspmpN5mJ8Oy407EpsHEX1WvEzdwOTX6btAi8rX/K+ulb0X8nCoq5Cs8oXnoawcplWrnjXZHYrv
rUYLt1WpsElBzDljDnqB9JlfR11VWOr9iv2PHdEEqsQ9jA+Xa2rKMIKgbWsow+v/kp2Yj8D1QtxR
wfDYEwvnnfA2Docu1nxf4o5dBdms6fcP428JDvgsAUujpNhkQPznHtNp+FijrxXoGHoJq+LL5OAB
1Acyt8So8MXK4t1jMtzzoZluZWCwuqDUgAmhrRK8wBdKh+h8OrC4xsIz/Y3YjhBV0Q+HxmZE1ggY
wflzRpMCITwPT2Z1bfXDc0JiylDP69YabDfHC43KpHAw0N5ils9xq+6vqgGxG+82+kZnsKB4Om4e
GMfbo3LsRpTZl5+MaPQdvGMLHBM3jaEv0HMFtSjskgSP+RDFWAkKvmo4XMAo12zqFt/V4yI/+Eo+
+eNe/dO978R+ykuHRylXDwCR8iX0Fnrh43BGjx950Te28RWo05kgSQymDmjy8QHFFvaI1wFAklMy
D4lwaI/J67a5YFrKgFC2FTjUoEuocL1KHJvnCOgO2AlLVMa+z1AOL7+4w1Gj5YG8zfpTX7YSdBpf
Y1kZXtyP9r/XhIk7bFf7tlJZPzQVd+1Aq7iwVgXtDWSe4tSq3lQqclQVf8FCybtTgQEedNjuV86d
QpzKQFZWe9OxYmEbdLjrbbKShjUo9L86/ca28Mk35uXWOh7OtX+O/VKFWmiC+CfDFq00ovqDrYWR
KMzoYiuQzOys2BV52cWGFJ5e33wDIBV+eOL8cMRlRGBZqtMe4VNecQheWc+boVz8PogFYVPI9MM3
xdYpLTulcmkoSBWYW8emPL/aKFa8ulQfUX5tYx5OzyrcWiKRymtSmbsclsz9EbpFXTwX7bffMftb
vnZ7ELRBLp5zK/D1Q8510iAvA0eNGuYFElvL6vUDMYMG/vWxXxL9ZTKkWKxmXnBkmbWYBYXApYfp
DfH6VUIxeGiu0lGbZ8Em4HpV08PrFbfN6EBThL2AWhaEJ/YIq+Kv7BVkZKx+qhCTjO8Sf3yYASz3
ojfE2OofQB+sJnI7O3JZ3TUW0Yo8lj1bQkp1qgoRC/ZjsYTMDEy3NjeXf/2eUJ3x22ACIRNAkdOo
pS2AqoSOlx21fhKhRz6HBQk8rRbfAGAawP7Hh2lwLePVqbAxOdqNGPQ8GD56k7DHWgP1Mjfh6aZq
sDwY0w4YgcX1jT+aaTn9oXOWCxcgRj1KvuyNICyoo8AaBVNyH0BZ2PqFmDSh2S6SOGZq+FwTzpOV
NLwOOEPi7U9r++1rYBS4OcGTVi2KT26MJl5oY1Ic3D5C69KEmy1L9MCrRzqZDIAmpsHYmusNeMzs
vISFSCoPuu+YM7uuDhb/rhcN6YfhBkmq4awt4sP68K1qQUW9YwBgKwHVnnge4v1op0TvcBAqn5qw
fkh7OgCKW/Rv5kiuId7MsS/vILCk6X8MV6S78k83H3LugBOKHdpDF0ylFdS36cUj2/THTqSUSF/C
OKhNkBiC1VK0qtQ8lXJs7mFUnBgE10IwdjEv5FBbgreZ98nti7TRQdZ+wQjAzT6DwdIuNrV4i0L4
PmWoPLik45+3jcX5gqjKJ81uTADb/db2udQ82IIw6JhMNLisBEGOutpyUloIrZIvPTShb/lU3G8U
74RGG6Goxy3jI1RxI54ERhLWU2dCmpOtG9dknM57XFgLAQv5r/mhcMgGckLwnzaZph9czt6zfmIX
cHmDbMnGkVbmh9oKhmlv5BvXzUuqPJCrZ+6hbBz5R8pHWtc6q2AMWZQcZG64za57Y6a92fpTWiO7
xNyjXMYsFhWFu/2CG0VwvHQrQ8JKFQdvZTJ1t9lqC/9Y7ktESuODoOaBoKGZHQHugRWtZPpfsnd1
58Da2xUMkDMcJOSgZCwtCvJ7RaozLfz9FaI50oBc6Eh5QTwgYD8m40vUL1s1RCF2akQCvnMSxQhI
AMgdEJmKUcQHHOFYudVjtDPxVpSAugrLnFiE9x5YzhXiMYuOaWU5Tz/BWFPZCf4m09X/1BLYoVMe
2kY3nUS5Q1nZkBp/g0pnNC5TUzrAzWGBiRlyjn0I7HG0USydl9Gj3N0O0PryW1/ieFtclhcYomxm
J9YnKn6zoOCVJ7LMGl66PqJyQgqbSxpCt2KtvazhNHzdYbf+Z0flsgNqUGQAYyAUACtktobp1vrq
NupOR5UyOGn7jCfNYnGTFWvmrPIDcbpJ2IbOLVqgTSFMQit6f9KzQVWFEVLcySnwaUPNjulSgkSE
DZ3N6HVIUAAbP3+z6VezGw2zkfu8jXJAYkZl2/4o4kKDJJFXBjrpN0QEp9Xs3wm+Q6egtA/bsy9o
pMnqnZRlijqW0tztVzgWKBgn4/DupSLrjvihykhZ9cnPJgilYeefO7Cp6KQ3+eKOwBY3TfKzl9aK
2jTQMcyu9A4WHr0c//u0wsI6GCyANNzvGWLL//tigPGQiQDi1iNmaMOImqD3vqvRsY2K//VEmqAx
uknhECGHBYIxBHINgCNXnXRxsOTJjVMjEwMLjr1H28stDOrFaHmuGOAu+P1aLATwp2hAiHcFKleS
+aKniRpxN34rm2xICATk/4t0GKk0FoM0UUwHdF5wshI8UwU6YPWsZunhi8M8W7jt6Xkxwg74YHH7
+j82kw/GdHYEcLsfhNJUfcpVrpyga5oPPpqJzNeUSYb+zVmXhmGacOkefOvgFk8ck7gk/6h9wo65
u4sqVZFK5Bery98y/zfIwSJX+oUmTlBptWdf8idkWqNNJ5pcDMKnu0l2Z7TC4DztQ2c2TgAKot1/
uFcFNXyTwUuoaOP0quv7vbgEU7OJvaWVyTFYO1EX9Kyo2fkJAk0G/DoJAbHXgRFbPqoproL7ctjU
L4A5cHyVGa8gQrh8jJe2wmcit+uOZfo5fgfEqKVb9ricEQwRVGwBaoBRoUWCE1Nvucj18uvqKvmE
6zmS7dQiC4Mrc9U4q3eQ6u/+V2jvujNQOwsC/EzVxcf6Ch7WkX2J1JSvo8TtCyoANnhAoeZcDzpV
t38/V5NUnpSusjLNp8JWbi5CCFCapOTJtXH/f0b8x740CGqc0JM/4h4pawgnGINnz2lKYnH/4R8i
M1rGMi7baiQbNFjY7LccTAFOMgPqm41OYUMH/dA11ZUTyTnYgy7z2U7n/DPtho9vW6iHrjG1xF6z
YpUbr5at3+Jh3X8K8qGF3pBcteRE1ZTo9UyimSWSCEs5cIbThLNiEpqya8QCyL/1J6KMRYfdAkWi
vpGWkhpJ/7R47BpV6+sCco1qxXDZYk6tSJ7AvERfRK9F80tHrpqHHgtprEDJQ3TE6PNn8iByxcE9
BekJTX/zh/vWr3sIG79Aa1sZjdxM6QwBvmqjqdYt91Tlvy2IlcnD/VzTxZpeUxFeJq4tJ0lxcXR8
g5H/SPPPXRBUS1w9ObZgiujLLCizjgiowmJtwtb0cN9eKWRrTsCTXAMUmDzSR5JFLM4FHmLMAKFM
mDPD2KkBr7teVZYxIema1AOLaOnaPAGClspy5sqo6h+7cqAVYGmaa8ef6b/aC6VnrzWP8rKjNLzK
PjYsn7fGdPVjBqAoEKcB7nEZDPVXgyqzuJnbxsIYzdLKEHcX3NrLxauDWFixeD3jJWHwcpkKWG2Z
cSvdyEvvDeWTqlayLNw0Jg2fj+jop2tHyuPCBC+EaPaBR+g+A+KJAA1Z6EYhJQPrN4pVEiZEfEn9
P+vR5dZyQImyVkh5HiSPxyZhQW1F6RNJDLG4dzQNvGn5kYEfRGQm8WDABSCOiqO9rQDFhFdxWVRg
UuubirRkxjUzE8pioo9bP5NM1KU7Mk0+23vdHhH6O/zo7KqcqNZUFdEB1v9cHvTkW/9zUV31PMaN
uqHqt6y7Hoes/uoZAfWjpcpgc/nhaCxGd3hEnAFyMbZVxLT2Shub3VqlQqq258gvB+VLw/5x4eOk
SljGLMsEfDVKJ5ykIGSaL6RTJFDf9rhrc4UUcWDoa3cUrA1Yj+VaBJ0e/GJap4ho/oopSxdDUbOR
myYJASBXKlEWnBfDr3lh2vGUZMzM37/x1cPbmLtkKiyaL6vXFPxoANbTxUQWkqndaBEdUptAX89B
uPHjW1t6WpxcbsJ67/9gMkAu45lFABl51ACZvTNFRLOGDbWN2mduxJ3JmqHhA1D4x53zmWq6ahZ+
zeU4cmw2ZqZHlVKCdCaYrNHE+I4Y6PHI8eDOUS2pUDcqOfV3HikaAnW+saiSWeU3Hde7waDDwa0p
ZR8zjpxdJso1DEC/708zgfDkCqGfbj/+6CIefxuSDAND7p2g86z8dInsj1ioXhctJk8iFWvkcF/n
sTsH+gOXVIkssEkjwGpr2P9xh6k3IkK9mua0JHXCAmnyLBLCA4CccYFd+A/yS12GH7WpMfpBGZSB
/L7jyeTOIcCRbnH1YN7oz2+RKYlbuel5YU7raLXJEzQrCR7Y1rnQnFUMjoAwf8tHmLBecVc53pWS
ZO7EwOS33vXAr5isaEPJKq/VyepyH90Wj08pkCiWrq13ixDU1Vmh7qJ2zaIO4jcsmTy1UhOAwinq
Sc018KhcaE+29TxLg+h1n1WqQf7hP9xo2TFFUQQO/PaQKT9qb66nF6j4A7oT/E4dnRduuETPJUbq
lyXIsChkgswQ/V96EdzeHKhPPIEaFgXw6OfqAQNHcFmPDtI+iQiCF7Z8FjqYovwLWulq0IBTAUX6
cxAaNI+PbD4phuD3wWYIqZiWYRYIrba5VW7DvuHSm6kkKPNGF37vuJFxQwPYXFzpwzZB3CHPba/9
ZmtdFYQxEZNXjCN3SdrP0dXUKAMzyC2TdE3GOhMCJxHbGRPvGgm09kqEjnpR3ATUMsBD9B3R3Ww8
aupN3ClHYRsGF6niq5ME91uX3FjQl246CWSqWNOSd4Icebxx+NOrCaEQbALPjSrSbeoCVJSi33ry
UNzrAMQKW4/PDSGrltbAHE/MssrLv7yr2joiPQvDkNXP4r2JdXiAl3rzThuhb3Gd97ocrn1zJPsK
24XoXPK05hdJcrxtvAjsz51ioBkp5YAlA9lNOQMxrrVF0ccEOoEFN3V2GsANAfwWcOBRMwo1XNob
E8AE29xAaaKuateFL8+y0izkmXYQMMEyN2tvqDYzJbAirmWRkl7bKvquQgf0/YW9Nb3zTTTqYFCx
mS6AtCzfbxfsqqmwe8NxzgFHt2ycrq0XTClGgbnZfKEY6dtjEYJlC6A6PhLzO9t+ND/npUh5zW9/
f6E8uYunPpTc2EIwiuOOpjpC9X6QEFTNWO3/SMZrt/WAdeLFYKZ3G0smN12Jldk9FpUFNj9BLapt
FaXA4ewiP5aewPqCur2Gg2iNKl1duuHHCHQr/VKNzEKsAF2MKeMSfrEVrihtiCuz3frAhDaa12fW
oeO5I5WL6JHaaB7NATVAIUQwlZXeugA7KfQNOWV7oU1LMMuO0CDnwij+v3QMf2kmogaEFS/9chOj
sZVz9r8ygE6stEPXpqjiXmGV4vJqfSBfF7Z/3YqUcLCSizCoQUv2jTF+s9dpa6o2AXEdLtjbsKUZ
XREEcRREfrObjzST66GKv8rfzTJiHgl4aW3ziCb/aeZiMz7xG6U4n9GCwlNGKOkPbs+Tafz9epOF
xsuCEdLz39wQ9L4OPff3zPHke0HFevgBz0zEj6Lh/fhEKV6G4q8cqLJLDYdisXle9Xg2ckEMvPMy
othUjlK8ox9GRvdi4RtJPF34hR/9+6p7UNBzokC7gY26WBcV5NRxie3kS/gvmmGAzlZnX5nXZbs6
pgaSE5RIHdMB4VfdvuVlX0j+DBtdTsUeUn7CdlEwid9PBIYNuAuGwerfKdSciKN45Mdp0stCv5lA
OtxFOWtXM1Dk2gwjaD0MyMpSYlkd8n8U6WOuzOVusKWb1/1YXoHIAHAidkI8k43aGyMYoMsyMLud
KcTzQWtGccVVLBAtT13dq+6g7qATc6U+2r4PRw2UJ6vwLSes6tAb0agHxwkuwP3hFiAh9NeZU3ph
l/MKHTEix5pFb3zGaXkrB5FHTaTVVUzvoMv/0+Lc5PdwYp2/CJ8COSkP7IhHpnUFaLnXjrRrqgdw
b+Z+H0oxdhe4vfhDhEQkGZWnHSFvFdFGg+xnSUQbFTGh6KpY8P+PilMwXJmDCZHBY9QEyHzUhL4P
32WYt8BzvJ4TynAhFFx8wOEsEyRWQursp/A+hCKvjSPdb3Zhmv189j+63oQ/aGhUnBiByKPXgiis
K/wc8rJzTd234mnE4mHQE5990LtOhsD30Nj3+hWQldOfBw2ffg7YMs6oacEe3b9ojDd0575qTn+y
NLT+lqqi2CvT8kDhfSJK+F7HxGxZOi34S6KsXu71wNGnwvKA8AC88bVr6UjcE6H1pxXb8y6d29Qc
NLzI4NAynCEKqHTX8yx7Gctr+99Ri96BNEuN5AZohrnkcksT9IEMcXe/RQUjbCZwbC/NuJhOS83P
YdCoCuc/wmSgfQFE7Yuz0/u25HKq0EtGUrqr1Dp4+J7XI2H3YZ9l47P4/pBXtF7xFgkj69/NfOhx
5cF9QbLYQ7WaKmtb2QaryUX2pfsPe19XioY4A3aI4FF1yVVkNJJlG9zMrJasJ9gMqlbvZl61qz3o
uUMiFFP36zouYBdPhWNTHde0zywd6Ml18je7dimhvTq+G3EWF9zc3Nf1B8kZn1+rYWyNwoCGHjDS
7RMQb1h3w9Izu8Jqu9IVJudsEP9nxIbwV+3xWsVpl3ekq1EQ/DFgkj6AVPN45QJMe3QSAPi1zpGZ
MNX0a1Hn1dng7N3smIs4ubAcb7xWhmERvH634aILCkqH8enNhMjyticTshcrL1+hnOm1/HvEV1qf
9+i937WTDh9gwzY3P/2YAUai84ss0XC+nDL48aRGI3vdstjcuECY4Pr8PHJBMasQsE1nA7817AUd
Ex0QlX/oaFukIDiE1fhKX8qL8exz/oKPw9GHDsP/qn9NVFXuPbsPOqlRIMUXyjdmsc+k2Xl+k7eN
TnxGnJ+dyHsqvG68Xi5BriVdQ3txAfbIqyU5l1kueZ3+ye0oskNtgg+EGT5Qaf+2wVpIbho4iYFz
bIpqL5Dmnq6gKC0RYD7yFHbixv86uOxkbJSKlpn7vYHBhx3QOAOMP1GMUN2/wCQKcAxlhVBkmD6i
igDsowCOjS7Gx3On3It4a9ZwfLJPUZ3GdAfRXR0fav5YBLthaZV7AcmPL7sEk4zyH4fn6izPv1wz
LhtsmjUpElbhZoSB6OjYKMUy3a8h1enGQWFwnyY9LCQV10frOIqIC8rxi8PMAFYa8OgBzGqukv5l
uiEVwPUSr6ewqzqOiTfSG7Fqd/OOMqkhNSoycCcOtDvrrIBxGKdhqPux32zCP31kcCcStXH7G0L7
4IbqNPpFecZdxj3z95nrcc7U2wjHzo6s2oGFMsiNm8nxAM9UKbc0t0KpZ3prUP2uFDzIsjhjEkyH
flzjhJatLZHcIzezv04HqqJc+bLcZ0aA+DPKoYyKlHEf3LxFOI8GT4M1GhN3Bhj154NZzKfVrqPJ
ubPXansdWjPIm/4Ifb/WO4CRsxIjxfbyi9QrTUt4klj36fcSfCo8VoFmzaJJ02poQLS4lMGIQ+lZ
nLpCmfT4F/mW0uIE/yQ9bqEUSjE1vJHIpfB3mUi6VBXvu4X+4S927C8Z3zSn77Taatx2dAXiGTKf
Q+sbuDA4kut/jNLW/Yfx9hGbUE9TeOgzb5kJJ+hTUMgcA7bQgxW1ORoBCQPH39hbCW9ngZeAHLiQ
YXZd7NUFvIDKHsU1Fq6SJ8lYZzlDNYvlzrqEexedvArVv3Bk30gJKlkf5TahIV4gumXFDfB1vTaE
iVIfktSYkY1iim4UfVg3dO1Z7C8eucM4huOWS9K0R9SYjYQnOBk+FlGOATcQg6YwTKuxIe5yxnaZ
p/7f/fKSViwo44XIRApmxAlOEHu+Wt3/87VjWqgU6lJQ+/QjPjoPKAolpQq4A0PBPGJJ8/tV/uQC
SVot42hRS+5/Ky3391xhF4BOnrpcVLsrjZ233zNUFs6cpfxxtsfEijCOBhYkSwFuiJVdKLdqbXNU
jOt6fyO48vqxuVE6VUKJ0nKvL7wuw2AaQN3XhJ/ZzQyz2/Z3pVbJgkKbwPOVRAcSQhvuHrLe13HB
wcKz6DAnfMHsukRgm0oXxWxKp34DB+qj4HoFOmN3pAGsKmQ5x3svtMTEP+Eidw/wYFeEmGZA51h6
4QcyigNy/FpKr1myNOkKiUAvf/AySVy1xwhUfpDizAnUFHvmzZVF3SYfSFzzagfviW60h1vrKJyu
phEWYh6FYAN7W79o7HtOZK//Y4+EeIPPhAvhInH4r9WGhOVvk1+A5Xt+fWw9Ul5KO9K1hAQHrlBw
ox2ET5+77H5VHT3ZHr8B8plj1ceOk8qAPz2Dy1BcdPWh2N49YLVV1JSKwCXeYOcv6HNEY9RwuGeD
o9PgYLaSqEfPCnQ1D6KbVV3gzm+CDDW+IbnBMiQUxMm86hMj67Dp25k80/CmEkl0LCMy5yFUNV8s
v1wxwa5HlUJQ/PccSVCdAICH1bEdj9Kpu9wpfVNPC+OKkP5J9yTsZgmfbLRj+rTeCRGF1gPJjUih
URrN4WLM79HAbJeo3HkzNwIEcu2Do1So5VxE3963zObSmLLlzVuPjmnX8TUhiUcciD1xzrlGDAQr
tL60hcU1fEixPXup5ndxWxDi/ssQaz9vht+gRP7PpXJm+9K50kfaaGp2xfaHktHe7pUmip4ThJwq
4DzBaciAg8PUUhb/jhelYkM3tri/MwWeKqRJx9dHTsuUPigfkb6mw23/t88UvlVMPGzhCvfxGo6n
Xt1WARUGaT9VXZFNOdyjArF+8MqlSc6ST9BWzKAJH2YTcTVShEWPCTPKOJtjBS26+/uDdbSolG1J
jtnA9hYosdJ2nEQKFGtfkiE53yTuG63d3oWHNDLvXLkOSrSWBbDMMsNcBlKmCZntBxbz+kRe29o6
8yY1MGWQxbeHAvvWtJegd00PZ85k+Jw7B94IKL9kYDvmFpXY+0XXYqhLCYm6YAC+Gz9LPUoImiqC
aWCj5knWnDVJKlMW0Gp5JBKhsmYFBS+GRI+kPAUFJT0LB7LqAd9LvW31XoSKnvKdoVGG7LH8+9sY
PrAkJttZlNPWyAo5WVY+VAEU261xpQUhiWFTdUGZBVWAazXh0fZiYN5L0Et/UT7YZhock74RJ+KN
2F2pdjRrtVzqZFIYACLaTZxOhu36viAoNGotD4sfm5yf57++ch+9PjH/ft8JBZXSX5XE/SrI4/6E
n12YSyvwnmKua5jimcic46ej5Hbh+5myVtx/RhNKp/sAw41pYzf2vDQ0LpXxF9hnlzKE7JFxTri6
ulOybAVWCL8/X8QWIcoTadV7DA/5YyzR1u11OsYtvN/SZEZrS3pOVlyN15i06p0rs+0X0WbkbmKt
oToTIF3cxLgbdFzJqJtd+Kxb1r/9k2wymaUq7eNNGIVVvUzOPUc7ToKnn2v6YddAO2wh2VEqUskl
TGhcFNIsKNVCzkFI8Gzx5xvGoVDcwywV3dJ09/wB0n6Fk9HYuDj5bqzxLVL8iUYUL6eCxrONQ9AH
RpjAWOkzjRly6XVs3LDh4zj+6JGEzFBvA579Z2w/hk/o4V7bQRLkt3zRS2sD/sJyE3h/Lw+3M998
YjS+YQVxEel3I/eXUUW21gMdwq6tDYpBEKtfClvwCca1xng8m0AeROZI2gD7I1zBZhdYKFygHKGi
nW7I3RxUJpDF95tyfDTm9PgtGehGXI8VBTk0WWLPSSCooogLYKIebWPChi7R16U307cDpqSnYBx1
D2dgD2/7vWZtOEw3ZkhhCRlTdboHhUsODrYr0+/bMcQyQYJZBcF19zUGt18aBAH0kFn9d/TnD953
8vk7hdy9O8aswwCkYarJm2s2yKEQPO7b1kiQMogMD905Al4IE7bjdw79arRX6YKPMoAr4axdztGy
wi3O/wdAYl+KcMKPsQtV04B7ldF8oWiNXWvKNP9L4PFyV792CXV7ONapjB4hba8HkmVFD8vINurv
RLLHQygZ2YuqgvwkiXlJkjpnKVIXoPkLufQTripDOZz89jgBAPSdRyzBO78yRUnMp59hd5AINUjq
bCklRwufKjUIJ8NFaUo5IgoR+BZYOYO1P+Hb8Nnb+oPHgngQpbj3iJF33i/+Bjbjrf8N0TsS247y
EtgC0WqpD9h+0ECBHzZLFeOuIvFtvCyDypT/SIi+epkaARmt6hQcvD81O2uFn6jncuR3n0MLq3nY
3Q/8HtGYO7dYu2RJsUHOGl3FsEROg70byj1bAuO6wtwQVIDkEIz4AIXNMOiDZJqwb1dM2Qj43qvk
55yCc2gtwcuAMmYqtaWWJvG/Jio7pXSn0Zbs1f94865B+dGTff1qF+7hkkU9vAbiCQyjfcZyvQTp
2cJsgHgw9tUmMbLyGTzpSMsuFkkIcopExsuDSkKWQv7DvfhMnSrAQWFIwOxefI9/D2aPw0H3hJli
CP4kgkcU1aWZ0qg9bzih2XkXxZ1rgNXNZKqWqzw8wcrfZ25uuyAYHGCua9tJpHJuYpmZLKn17lzj
F5sIfLvKfzwvWj6lMfBDfdnbQq2o6a5YB/qRoTyUoKmtbDoM83dI7St6TIQWK6fazg3F1pM7r5IC
ma3PHlGV59ayCcwm3b4Q6BKMN6nMv3xyQ09QGN1RVP+jgxgyuJHOWvHtTzI66CvshK4+fKspKHIH
aW5/JgsNMFDJIjNkYmh6LFRxNG9neLtqeO4p+YkbcS9/WvLIES2Q6BUQFaqRH8f7aSytzFa+H++/
9JQ4Y71FDHXrO2bwgyc7djcv+Z0Scii9nXd1vWKrDovzddQFvOgynrSSAgS6xgZzxUm+uobLjypb
C6DEAzDHoZWP1Hq/kdRpnhmLJvGF1+ExCIRDcs4f1CslZ+yySBeCH9thzCeoHaCiWkJmwimeyr5j
5c/toaUIEBEKc3THVj2CV3fwgtoVMMHTfKJ0WDQTDkvDEVmi6GiJFz6Nf/Hoc2AUOsL8KqT+kqKX
P7R5MopT4IUMg20sCmE82SRHyIPQM13rLWiEfTOC5cU4VLK+avtQnL7cwC+HDARnsvxbdqaRwLnf
sCNaCt74jSDpIFjnlrkoDyCymbBbzj2eF6anJzltXcgWvfOhZqtx/LSGhoNZCv6r04A9UDXIh8Fc
WjBjAomV0fC2B4Eo5fBrdglb8O41RTykc4o0nY0t1D5KPUS/S/1JZTQ1AXNYm6UPhQXb1MXbTbTK
fXPBxhsyBz3t044COiFyRVxG7xFruQp7rLe1D83SF/MmEcSY2VvydhttTSU9SuRRcbmvNkXIIbdH
LxoDa42s+OkYDMbPVDHrcMmDgl5UrUTAvekhySnNaSyHwN/cBDnOXeleLbe1nfl63Q3B2M0zTmfh
LFc+0rqgP6vAw+93zmOnoVs4p/cac+cEqk5Y8P5IIqjUDXa1EUYQOFNrSeY9BW7KB3xvFxdzSnZg
Y44Fq0JdKNxeQjvSEuL+Ip3e2TgYK5dmMTLd6EAKQBus+AAX9WVATlfRD+nZphhlr3et5b93JFTU
GJCghLRJvDtKppBVTWqIM6my8p5/c+/HkNxCgFrSk0KAyGeqhrJFe8CbHkDhcY2A6P40OzCAXic0
Eab6ovOg8L4zKE+HGP134XnCr7B4Mzev/yxDXbp7WbTdcov0BkvM0WPwTWn/fk/HmFD5QDGummXw
1a6f2gih9pXd27bsQKyQXpnjxpsSAioEE+Da94Y3iObGknrWnxFdH6ePpLeKE2ZYdc2w1efw4Fgq
Z0Tj8MH6pQdGiE0D0zIz8LYgT49/kmF6h2nPCn9koIdz11h5lznCakwI84u6NdFRAnsFuOhtSF9o
lNaTi0ttwI/THPsxQEwlPmVxjKgVLfRAnBVJlU//F+Bi6JZcLJAf5cRLLZi1PW1xmEZgR1xis45O
7R5oTlJnXFhEINqJ9ah1YOD//GhO9lnAX2gBeWP+q5O/V0obcicDS3s9AWHnv9oc5JAJWL9CcoqF
r0rIcS6xlI6jfrYg60+WV06KJ3+dElJKshXP44TMMVu1j2uzhMI6F2jnpeK3mLIqcpxL/BBXzKms
jOCgWZnOvAboi+IXulndxJc32C9CgpFwYn4MmeH97LPBJxDUtrBSyxpkcJzcsSsyUfeqJ0Qm6FzT
fs5PEtG0AepFxPCk9otO7Mnir54ZZnss1IxocWDcQk3TdXcBbABxVOm0T7+lmC5UBjjNRh8fybvh
JG1qnJaYMwJN9/bM4+UY4dzcIZfplTNvaqGXzjtywaV6JZWpP+EGKF4F/JOmRruKXRe2e7YI7PJ0
f00mImY2crkC0ippRGL7/AKfje4dDMCAsS+uJ6bmxWFWjpW8ETShiACWWil5PKGUInMB+971Hz6c
gSKyuvcVs3CjgajtdnRfcBURspeiVZqXIZP6EiBvGXIrHYMwXABnk/HDYt1jTVCGVzwigNvwDsay
kMqoFwvTyTNPGGQzHzaoKuBJhZM8okuX7a8MgnBQ37h3+nTht0kajgPfDZDHDptjIqg7QC5dh5vr
MmCc7N3M6D2BNQ8KK/8HmSXw19VSoKsY5eRsxd0frmxvdQOoiFnDZwKwvcO2CVlCDHHaTpzIOWJe
Sjv68RVWN7rviluhPBqG45TnvMzU04nCMqYr8QloATL+sOwrn2OYuq4yBrBumyf09adjhiCkixqz
ErVInwWvNzxx4cmkVIW3AywPSkld8PbYsDwNWXInsF/Tbs6PUpuIxDLMZwEXKlXmiGUj/njJ0w8Q
XrkBUYG7pvFDHH4a8vlQC4ZIvWdeAgW6fOWEoCUuUpSu8KcwNXnsBsWeTvlstMN2BYbFa3bCKoR0
cRpsWCZtjFupCmSb9ZckETEslJ7h9lNZptoTSPCIbXwx6OF4gmU4Nxntz+jPYVLtEeOKBYqbktIj
sYrhdsPhhsOgrq7lcDd+aDck8rfyMYVnJwVmOJkW4O0Cmh8PEoFlG8PkeSObdNRSitWm9BxuUWbA
eWypX3H4qglxgXWv3dH3ObLqymRL2NX5O7SmMjFbHYnZIbPg6Eqja+IGjEk/yE4DsPzK+MQdS2EH
W7L+TGepxpRTIdzAv82qa+5X9eL2OnL+LbE+aHEEQvw624m39owSasDSFzgbQBhlWQCtlJEI1Oj7
Fj3qzJviAy+B/okS3+1iXUBoeYkGQ7UYkOe10E/R+2gFA1tlXeLDCW380Bf+lYUSIpXsBnqqIKxU
MsyFi7k5h8Ipf8lb6AMV8tiPLoo2hRlQICI9E1Wr+F2k3p3Q/xtIIQ5JpFHX+Lc7xXqYjd19QVxG
FEp93wgwedggqzTQWpVLh/pyxJR6CdmEwVrVXIgHGG37UtrW0UrPMs8rNIS44Ok6/Doko2iSe8RT
NqG4GrBFDbXFdtXLiwyrclYwPVFgmZIAtIVB7w6Ai/J8fvyyaovTyETBLzXXiuvNdZhnIi7W8OiE
I95wCqLfPLbC33bfhYpqZWC4fNDg2mA839PBvZ3YBGo8erKaCbfs62CKqVFYuILRYIRyXbgsqi2y
QCpNUAdNQm8RNiDER7sCeousLADuDmSeKybJP1RrhB3HqGuJ3ALsyO8bpq8FgamzNIWiGhc9Rwmx
m/s6QGdKM+RqTBkJp08kDywl0niE5ef3uzKHXI0FeEP508N9owY5Uf9TGlZC4Z4ZQrWrpuJsCkOY
5eK2Net4oghmjW3MtTcifq+hYs/s3wTAuylnDfQTc8fe0I44C4HVahjTkemfPy3asnkEkrNbK+dN
nyX3p3lv6dK6NueFNCtAekMERdBbt88VCKB537dksr2XylKG03rBhB43ancPEd3v0c+vhPqZvWWQ
X0SCk1uWESVEgCeTT0XfYfmMBJ2Jmp0fN6b5CMjx12kfUuSjpxWM1fTqeZHtLJrqT/yBlVxJYiZ4
KaQ/JSEQSfR5gzGC/XxSIzePJpuojivYw8C9a/9z4j/0AeoOuEnYjfWNgZigzQ6JtjBIU6mx4PLl
QWgFZwWJ2zujhLDw7JcYJlC+Qe36Uef8uNB2Mz5fxQr6cL+QRQfkby2Lam1uAGqVmOqTmB7hyV1Q
PJYnYPIyZcP6qGwjWSqa17GUwOQ8FxWqSpqJUIS2HIrCtEHDy5CxRib5GxdLDpcrXYdJQLOyGT57
ht/RPrqA6gyOuq9GN7ZQpZFgchJVR4CQnoKp8C9dmqkdcxkOg3O2U9pSBJg8OhRyvo79akeGE23p
21f+OuBTNTHvNwo31tmEXEFw045MkTx6NHL3znyCOM9rXAWRX8zibfetObtrzk5CQt+hZu4QPZ/g
Rb9Af81sX8+CaSeL/xv0ghs7gHimSI1XHbmPHFwgu4QgByYEmKh9rbQdZIfdRolUjbaeuykKwi//
wvLY8ynijiDR8nEdsuxRI/Xy4MjeCMHp7Yy/Jy+dKFp9YaMhjEFNpXK+8aYUQWHf6prKojgjAQdq
//Sn46aFRi1fDqNdWkin7qKkrp/yxVHiZdAx6eLp0NOgxQUQQANLx2sAR5upw5Qq7D/N66Pk361g
UIx8UG0P5PO+dPTgsRiHvcZHYuEky4I4Y4gfqEGZwCVlABPm+WNFQ4Oqg7T+rTRYxOsNxO7AVWMW
8FyTdhbIy0zD04TrC9UlflL/fQ6n81tr7p8ODtxVs8iMz71QdUBdCeG7F7znNmZINavMNH78+VrJ
PUsrgN9+C/06Th2gk/n9o7c/2s1o+EwVqoWvB7O21Rd5AGmQwGu9lEFTsyvFSD1q4fKISjpoqcFL
GmUhRu3qhwpCyi3UNgulTw05DyjM4UurmCTtD2YFsrlIJqX+XGUNl6+9XMMv4cdJPXtAsGJezVW7
isyRV+PEfachdhQZfjjcaHgm1vTKA0TH9hQ1VmV2Hol7CXdU70VKH/980Ew+1rFqgoqEawThalZh
0Iu1d/ie33Fwr2ic10jVdJuXpRjhh55SI/EOwgF8xuX9QHhGyPH2s8RLrWesdbmKDwK/1BJsxTMM
LJUKjeI+uRlG9wMaICcSmK2ChzVF5rUd9yzozi4EgHeDHsblTghsDt4bJAo1Vg5rihJQeRTdVIJg
alDBpDSzMKCFGB5Ao76ngKwtU8KGaHOHcQW6rhxZahCmjTr4xVxDSdgwc2XA3p0ZKCXQMpztbE2V
uVvXi7wfdioVNSYBONv0B9a3AkvZVWJARXuQNqC0V0/ATx7obpBS8JdoEZDt0YUxu43RSYsW6jt+
00LFhvwamLkRV/3JlmC3H2ctMCsR+bZ3jexvkY55t8E9s75U/zTcNFik7BT7L7W9pG8HdVgGQ/7l
LNwiBzBrghaSsm4f3l1xaRoaWpJq6WGTa2IpqRSGV1vmnzmmE3pe7Y2Im00xlOrke+gzLroIRVvj
Uav0js4G/shRJoJu1X65pfPdLYjwi5ypBfzOkTG7TTz/Lto1ygNWK3J++m3fzGOgycsOd9p0ew2H
LIOZ2CoSGVsCv92vPDwPjdSZSDaq2iIhlSHTSUZU9iDWI6qp1e/nT3a+f2fQ165PNAhhSArsAZeA
aHXfnlBOgY64/xq448ZoFrFWLINF2KmQtQbxiBSOmB762fMcx+CgA/EzdRp+LlXhDc33jasfSW7g
knZwHLf+C7BIJW1XDrrBg9LYM88j/1dWIMjytVHDiVsCs6t2/NKaYT1pqk88wkrsHbYZdjFFcEGz
vghRdxWkRZK26FZrWPyx9e1OtSECi9ruS/PPoQJRT3gL1snYZxiYOBuSaOvVV+Ha/6chlon6iptp
I4r6TE996DJ7TLmLfWlRwOWeJJDwVQHkDafWfh0PHPy5y9xL9XHgwF2S1ZQidDTnf5YYtbvMaJbE
U/GixrtdR3Oh3qmUvy/pLswwqZlHS6f6Ecpfy3RAQ2/1qhLoBgZwcSXmnaLkstw/sUatDbuze7NZ
8BMZMoxQp+BXmMTaK5BdfvBTScPekg3xtbd+LD2nMUH/ucIsgdR9c+SsTUp7rUNspGgaBL4fUpn/
+nJOcw8ld2/5jvSAJQcm5qEUiu5KLP6RCoxVooHliiNe/zhRXpCDCl/fPj4Oc5zyw38avJgf8nvR
ATUQV8xmcYxG1bn/LS0Yu3BrFnVSdHrc6W58oQ6OncXcYYmaUGeuBgRT7yI9Hvzz7GnW09UAfsji
RBa6OnH+wY0NCPVjr97nSV8LoEo1gIYDZKYv7aFdu1StyPSWB8HzbFFOLD6LjjFOR/dmVJp/lepO
G28USiDKUWlOunDFf2Af4tg8TSqkhwAd7wamAE1dly9k/NmvguGFIfsaDlEGOEZ5T7OvR1KaPlcv
sgV1zcyI7GowbMspjWsmK7QcdbXRefXIFTNYK4VaYJMqsHGHWOmuzaOXpMT2wnuafHngfZ14nGqg
Voq8Pkhy++sE9fhh53Y2zg5iX3kIWppSsF54cHYRtJo/9Z0NJP2+VFVlWxoZRXQIpHOFJhKGDjGX
tQFEDSSrvXek65kD3Bo8p5PVoHBcn95BxG5Y11n5BWpINHYxKopkHZmdQyfFMVn4quaAZoTX8d8x
osALEYAllGkdNg4H1gsEhWDRNf5NcA59c1hsK+V3qLaHICnfLSbyAURWLPnmERnkZ3J61IGAe7b2
hMoPToaSUyutcUvZjNhiYZI+J58EBoz1oe69d+jkYHbzzKN2T+4irHa0wg0wrDn3gHBpqAIO8Suq
OywhUKMhRLMmmjHijU6bAazTulXzW0bOswdUxNMWb1hA8FiSb7V8fO989avOzPJjCBo1bi2ie2If
s6fiV8NR9cRu0Z3UEtlyXKERJV1/i27cEMNBQlvbGe8EgmyrNCgJAIfUyvap7LoebIqyHR68JUFI
3q5/aqqEALRVQkttWnJV5fO0CT53XSLMwpaBTunVAfeTtDPl7Ap68JnJ1tOOTA7uzaOTIORi5ve9
mkGDC3f7ak2di9V7w+TqL4I5J440TNXRaCAkQ5zsiDUsfdvrpaP32YMc5cq3R7HDtgDwcR45Xr1p
OetcDt+y3pSIUY7kX8UC7O5Y1yZtN8G5aXLIJcxzR0DVuL/qS8anzVg4SDxlT3Io94He+alasIIT
swFflILvYV3GPr2UxnfIrPBpAeMgXqcUxxf6v8+dhn+FDhliXE+mEY5JVpqaOpOkcslL+lAzOrpg
0gev4L+/A3yuUNsU0JT7rA9XMy1tEyuz8CbGkzJThHRlk3TS0GVxG1oQlZayZA690Rbi+J7v5WQI
d8TMsRXMpGY/+G7lMZ59VOAjF0Tf0/xo3XbikmkGmA9JHil7BkTcnlccLgOO+743P7ORZCAz7fsS
bASvq3ORbiUMExBBsBIZ/yyaWDfvLRYY+M2YVynG806JPp2oxPm+yu4XdVK//jEsCDkPNFk/kkON
wZGtNkkLhiaP41zlvgw5YvX21lNMuwZV1XVDsunaK5NahNdUMk7m+lickOoHr7bWqNRUpxLzh2l/
D5xxHceETHSAFI4hXWlRBfwf858jOfuU3LPUHEB5wAP3mfx5xvGwfXahQ+YhgMLZUmZpmIcvBmfv
Ndyu62jNS+GrAytqhi+wJ57F63bi+xugPs0CvuOnQ2AdfUUJ6hbwXV51b466gxEgib0ls6C3S9e5
OCP7u0D+1zGAki6vepcgQMnlnBYkPVKf4QWDIuD3TFTEi0IMXvjQ8pJUnGr/UyDqnfCjZXWq8vuG
kDyYNJ2oF7EZ8/H5Lvg6nZ7ImaZoAh1uac0RvEgjgYj5pMwca/AA7zDsNvrkZpkcaaMWtlIJgKIX
JT/+F5LpoaVoCfVvg6dph9SNfpXuoDj9MfHeqHV9dnSfMmEOsTf6aK8Nt4JgHqoFWZR+vfkkrWrA
K57CiNwvaX87+MIJW1vDeZSM8bZFidJfVQLngHnF+VvJDD6eUVyKVN9cra7nbNIUV52xWmoB6JUj
xR0OZ1orHglSXjT2X4NKysRYQpfAdimQ3wJ2E9HWmEJQWvTE/TLym0kHDBd8/edkF2TiMvWp7s4x
hxM6K2/D3Qk8pnL7cE0c29+yS+O95Df0/Aw4PoQT1Pip373YFAzsyOF0QBrYV0uzNQzpeVk9WdqE
bkQHRsUTdnt8DejWFqGX05TGnWyjNEIPj7+MRr++ou0lqQxyioRq16v8GLVKKR1Yjm6fptf+eYfl
eZBu150/vJ7IGY60htPeBPDYF74nYspHTbXfBtgcOWGqzEaXQazY+86gM4LGLKmiQZxJO47ov1lU
W3ba/5o1SF3vDLASN71kiymEk0NzkqSzTDiMwvs4RVz/l50WogBaqL4x3o2h3W/Ez10L1Md43Spp
cJuthahM1oc2cJWgPwmLVaRpgY/1Kr6ESQCHlyE0bVa/t3BB+DqlV2c3uLXW9wT/3MhFjCYaQ56M
gIJGPRoJjyl9EUfXj2frRj8l+tL96t3O+dOjKhcufMawcEmrLfN0Cw74dmkSIV3OktfBWCQVUyMn
LOC1+jbUZsObrf5VJIwrIRuVxL+5FmhBJkt9RUegtV67NoOhAqapUH9GoQVkRIqqEKSISaL9N0Zu
mubVfX9YEkB/13H9JYVozrcCcJRj16oUEvb1old6Pnpize/Y2qlyrc3UUvRy6+s9eTnGTt8p1dKH
SietvyS2zUMHAs0q/yMgUtlvPDyQ6OHZycTu4buvGTsgdyhDGARv8ztxY1m1uWR6NCllapCOhLku
jgnlC4/d5yyhhvlZm8OtwRCDtnJ37XJZL02EMvSd136FTy/XXry1O4ldOU3W8NdpKmx5lXda9TBA
d2MVNl4Zz9xEsSzarjLX4S2Sex2gyPkdq9nIOt0QHDz8LN0Y4uTDuvu3u7E9BMyfiCU+VoZIgLrV
TLN/RGkC9plR92RS0u58aVyBabSKZobZoQMGn9A5N7EVWy/kesVu6iCH4PslFRmQKkgcO2PYHk7R
UCb9jl6HDNc4V4WTyT0HejL+K80sh36rnrxewGElmkd0Z7nMq0wbNgs8zFHgg/gNMbOJLhwsVICz
BgehChpLu8gg8rDVVKYDH1Jl+ru35oihLIP/8MszLyI06h+TN5fmO3GQENSqmVkjOxUIGFprSnhi
FPSkQqbcNE8Fbm+367kXIyxtqQYJc6IpjI6s/lou3mx+e3c7YymEX+oVWnbjckoj1YUIEIGD3bH/
iOUwjpq9d0hDbcxDWPFuE1fzeGARcDm9CgXbLG3SlaY5E8E2XPty+xEpbbHs2xMZiw0IyXqaNhFS
sBiHDp8AMMn+nwvPUJPiFijcTXvoezeLVQK6tUNMnlEyl23OEifesybtLbFhZXI0dq4hvyHABjxF
fObNm0fxaKHTZNwNBN9cq3EFHKTdVMPgNpnQHh/FW7JgR7vsmEYxIYx6HF3FQ7Gao6knoIIr1zLf
fdfT7bYhDhZVPoSKsKKD2C+HyLj+ZPY4OPNxXEWJqzZ8X3ljXpUnEW11Rxxxf5MqphYCWeBZFGVE
7o9El82t9gDOwzOZX9SQtZH0H0ZpIlgx/acVdHuKVR9Jh6r5wP1wE7nRE3kUID9+pKPSaBB4TxNW
tWcwYP+j+qcPCFa6zgdOA1XITpALKtpPM8H7l97D/rOtoE8i8g4OCVU+TktrssXVP3K10pOzxDH6
r8RHweQ3c9ftOamNPX29L/Z0ru6uNJqRbpjTpwLgx/U32D9GDRBHWEvfJkhXrxPYnptThTK4s4Gn
U3wqmd6anrV0bzVTUgns5KXZQ6jsr8Kx/zhL9BGoUY4RrH3DRu4e4Z9rahnR5H1jWkWEMTWmmJ0d
EKacf8aCwKPjFqnD5C70bxdEa/gxu41zBjFajRKHwo78GKGfAHOs5ctFB2bbtHO87rsJiNt/uhm8
KPrXt+HQMR3yDGDEsraoLdMlevVr3kRT/Q2b5/GNqjsldd1Uh9R/ySCbRiJbtOpSHpHh0kCYP3is
TUPqLmUb8kkuvUtFATm4XQZIzAKfqX0ekE+hry0EgWLDA0MonswoBmVJ/sQIDXsPfoDAWOwdr2Rb
N7USslHY4SK+KqpzFTrsFi4pXAwG2iUyWPBslQLlWlVoaMWXxxWdtz1aPCVNmuV1KJtPushnITFT
t4VobWSkhMnn/X53VV18rFdUKNJNSO3JZ+76oDI77F63YktwJpRkV8PoMf3fS4OEMGERP05oZeJn
1XJQnST2sdh5gU5eb2kuFk3hxytQMV2a7bvZhE6VKNIvbP4eqeNdxa18RVSwWiVLBlu/eMgiaYzS
4cuoL3pQ+glAYOc5M9rhE4Bc389+l8M291MGAfVUJkGulGVE+HqgF2qX2NrFpIOoyR1TlGaDjdYR
M7ziMizCSCgzzRcWet19HpJ5H35KQFlf3LtworBKoisjMme/Ez5yKUYX8+CkOs9Bekd7e3nEI3FA
prCQp2M0sU5f8nX6y+YaYR+oHe8KLCZrSZ1wZ+bm6wNocsgS7VetqOQZGnNggC15gWdNfyMsV/tb
mOkO0A1t308h0T9Eo9OxlexADmqnzeaZXYkmO6rVWDMNwzIULPNTjG54SyojCl8omEAreB5Xup/6
Ifc61sDpqqBM2ltxmSSRn490offDhjLVGOCmofKbu0yzoHroQPJEoGnVzzmXl7Lg3sAlSVeF3ukf
7dJTo84ngspM1QEaOdKf1u952G/R8XnkoWzgMkgNb2w6qSobMm5XXAc9aIuMp/NUH9ogwSBUJB/e
0zdxKQAFypZ5SzVkf6xeVfwQkNnyZmQ9BbVHmIP6Ej5334zkHHWpuB9c/ZQgHYKuCVdOkIDRc+fv
NY7xnMBarDTFqYl0fh26x/WyF2WyFoqP31yCgtEnGTK4iFavtc5g4lmJPX3KUY4JEW+rYDLo0oT/
LzBj163oPq9C9AbVwmf1FRTNpN5rECIJLhmz2+kvKPrNfnIw03vUYRb75T0Aqdgoe83SLaC9oSL7
/44BJCWEVG484DpXCmi2MokSsOdnHV5vW796GePgkZcv4HWVvEYPxXhOW0gnwzwHd6wlO4z4eBoh
bIobN0HtE0r2xIY9BinP+1lidM6b1FGUEFsPy9KV6vzdLZqH0fpQ8HzwEJLHPZaaVzxL012ypFct
Xhdp9FBOsoLICIvl7PqEMSBlvbrnrU6yAjo9YHMmiAoqGOx1JXSWHVldSkWShrvyHhL4i8OHiaJV
i38YQNCK1enRCs39d3HM/803xnfQtpxCQCfcwLsvibhNTnaR2txJzEQ0oN/UJsBcxWWFZqCr6jbN
LITUmrYMPwT2yk4M/ahDB9qXnFm1ZHTiXQDUSdQvWql41jRwVaiLyPcjPofEDujbsUP3v9lNeawq
TVacSLLbDc0r+sNARQGKaYC2rvj00tWrbRYEDsFiEt1+2KjtXapTfpQXH/lOt0BmWYN1rtMM2Vqy
fAVW1Q4KumEJFU4nnKg6impi1Inv8+8xLGfWFCOLdvKMdv1WEokA2dtMiXjMYjVoc5LWC8CA0CC2
2tL8ukPhCosAVPqFqqWGayWAcstir1tjpJ2L1/ivDWCetC5jjdX/ims3rwumj/2OxD6K7LAFWIts
5c+yBbcOjnwUWd2o3XGFEx8ZYDPcr1QB5fEiGlMtn6QrA0Dx4vga2vSbNNyeidLbedqaCm5llRKl
fgD/Kvh+rqztStdnP2L8VPcpWEnddzW0Dhs/bbGKMMX+/+yMBZK+vqQ58DrYc1KdRLM+OjOQ6jhS
X7GjIVhCGFSO69duQHZQ9kj8/aZDRXLnxDuYyseX7QU9aEqG2flCR3Ot7siQrTMGrQm578hKUHBN
sLkquvXTOPrn29tx6RAFGzQ9cxuxWWl+W+owGmVrE94cgcoDQXhdFebTPf6iTPY43S0LILYIhfkj
yYcjqQw5YfwntC/Ezanf6i1XLsC/IfxwJXK+WIZvBaymtvQFYMxPUsJqRcx7SBY425bHPpP8fVBM
GshGyJYxcvEiYW1u4nY98MOFMzNvUtWhCDcL5YWYfg9Z5WkXokyfyHHJmAURzeMqCB77ql53MQXi
Iif73lUHkwpSxWNzwyvSdQMR148wp66EJSpSkKF4AJnC6d+IDDYOJ3bkLzBwl5B0vB1ufH20Hcf+
C8IxBpkTsth6jWFGFbF97U3jzqTt/BZHxa4Y6nXbuo97uEojOfCwBOA2swXM96inacWtAFunUbvf
kbOshbnVHgLlIllqOwS5eJjupdlwlTc6FbC4Q67+cRnEr9/O7ladxuuEzWzg88nfcUBn4cHW4EzC
irsk6zP+YkJWdEtec5KFLoaIR/L6PtNDCslUhNmt1BMMZkwJuActvpeOnOtIfKWwF02hmdP6bpi6
nb5U7dcLb/lNJItJYiVpWscs+7bI7D05juJ5uIPPf+cIVRO9JBuR1CBLcVQDlkGZ/ehksrExJ+fi
7ITmNf9c0stYcoZ2hewbJpoQKaqhSjNobJX441nVHKN9ff6xbiM8RkH5BvSLHLIQwWAdnbVOCxKZ
YNh6CJDEDbcDKyRMfqaagegXe9NRP+xREPnnbZhotZ9lh40oA8s8KV4XZyidVppmDCe7mPy6PEkR
GH3MBAgx02cNLlygUdHgMs1shuGohX0ARuDRSRfKxb7bT7DdVb9ilPZL7hNhV2w+I/hQFcBgWJaZ
MYvsrKqwt1LuuRmKqTuqioa4Uvr23IW033UwGOim/tHninBPI3MSoX8IoxtQ3KU01KiMrMz9hDj+
zhYvRHEyCyrMLvEJYc5hYZ2bpeGqHTxmTWnFZ1i6U3CC0tl1k52dGY5bIulawMU8y2+qwyzhBxw/
9JrpuIYMF6e2OGZmaJRBlpQtksR6XAmCT3MPNAnMeay6q1+r0X/Mi3dIda5U8HBEtWUGy9VSs7f2
qKy/piiyxhaB76Hyy1JUzUpTLWm542DYFpl4GMtlUByNNd4KVK/qi1BlIk9kKxclXtCq8cRaTrI5
6bL5HfzPvJ1Rtx67CAhv6FOC1PaQ7mgfqNwyMA+W611D6yLkC5hkKwY//3izLnPCOnV4bhBDmyjy
00ucrJv/OUuKIfNFrNl6iKS7z+3v88gHok7JdrN0D67/0QFIx2mN4R/vk+UqVPfgxLq46YmbxGTi
tphKOrvcf3c+DAvdI8KIPa6eo3s84yUwzG1Rgj8byh+8t8QtzKDjQSrvEIg282FDjC4Sn7gw/TCq
p6osdzVElqIlArzQRlw5quz8jRzNz1aciQKtdftcz4XVuzyUDh4MWfFO1EkLNNubGxFU0Oz2pRNB
e+lxTgjfLHXuBbp2T9RAvOat0iuZpAdueFi4Ws3+b9XfQZrT7A3ihYFzWpXikrwyNyGDIJYT8NpB
ld1K2SrBwbraMPTX16P64VStyGSpUg/v2iHM4hSWYHBw/ORGbwFrFVgHiE09DNsZVDSYKhIVhZ3x
sqEasIPtQ7UJjZRa997Sm6cZW7+isyfqNeSjUU9yjGiWgAEaBQ9ptmYqDNpJqu5pgcxmjXC8+WOT
lEIkvmW+CfpOJxT5s/kGexxHuria2ZyTR6yYD0OS5mMV75q/MXm5F9LFOmPMKZ3FXQCK+lAzMjGF
cMAMTpqviICHy9vY6I92qqUfjLnXV8qVOH4D1X+EpUzbBqymgLeFVSw1oRI6nn84CfVngUZXsVIL
cboj/ePATYcWnWVGMuNTWfaVw2Ki8zbC+4qN2MpyYEP28D7JkJpgYwiDUR6QhzelGyJ5iAXvqmab
rO8nJ6suLf6fR/qM0wH6m1/5wZBwE0strCWk1SgvS8HbOTPpxLfn8HD6lWNzY8wlm7ZEv/HefRER
zQWz6bkfpGnLwDNJCp1VYOpA7AdK/FDVZQ4LfZUhUlY44vZ+7SXTutAdggCul5fquN0TfCy3iwwj
lpBVzYc0k8lnfFcimUhy7eUr7rOpxvtOgXid17Xt0VUzrPihj/ggbDY7DmXfWQvgS6nguWvX4DW5
WmW+mS3++mwO/hvm6fPgzjmUo4TGm0TL13Lh0NPeYEEy7pwfFAtDo5FD2ZurF99Kj+arcTTacvaK
nX9yqfXvYUeipHFVchRhiUrjaBK4if0CYhdIkfelhITaH8NZRyCbiMdtSjDAzkoZgTl9+8/XfAiG
bZGVYnJ65jSE/1LFte9Pfiy3b8Nuy0CJXnAQtF0dyVRWG+w6UuvloJU6zBpJGzKC7BC3CAgqHmBi
mCUSHlCcld8qjyno0N/J1u7TjNjqIBhZ104OgbAY7nWD+HtLMUuojfmla5kP82eu2WS4Xt/mtAo1
FgkrW1/9sSNTB0q0MPuuzhPDOy/6JnKq4ox7NGQ0fBB7MDD7B+DlTn7sS/DbHh8/x5Kobvxh4HyS
UKxUm0DCA9aEBN3JOSN/F0xAdGP4vhukVnfXC7/FvMKC+eI0fSMyELkhxLWLHDOnDwq9JHtwhsiH
c3TEAPOJ/Q2Kd9cG2F25rUkG8Ywk/ma0BCm5SLXW8t5fEsCvVBjoSdOKvrpWMKNUbj4xBdRYnkTO
SIofG4igxfOJX6TbmCYJR7ZwLapDmBQIYoRJxCnpWKMyPB9JYgzBLOO2tFuMNt2msbTK/ZZurDQJ
TqJOE2nD98tlQ3Fw/reAp4jDCo/c33HnLKLYi67XWF8fAtpouQDwFkkr+hzhcpiMuYjpoPqrM8nD
tZ8UzDNUmRvxBxeh9NyAIlRn7tOz66X6rLvQpayTaj9RE9gtGZ6zMYZsVKRqsykYBnj+xrhjl69S
KM9Y/crO1UX7kIK/H5hEiBsFrhPmePTVjbTZWh7FQrYsOPAnPzjC5/KV2pArtkiyE/XjvWE2L5lL
3Mx/TOyRvZnRRSbNrFE0MoqMBHmBc67jgSWD2bgs1Gej1OQzboAmjzWA3EoLxMIjf7mouafd2wmL
cRmFws5Y5iENUm0wBysNa4CacqbG510x8G+vLgP0dBg51D2xNKNc+oxvkfM9yNtaWB2tdXiraXgK
hM/cQyinNoLfz19yELd+0sedkr1wQTTaQQB6erC7ORTSUfpNFONFy190E090D1yTusQ3n0tJdlDB
FXm3RpLi+ndnSakZdwC8ZBBtWH0GvB+F81tZU8ZL/BnA758EZyeEC/DfAv6yzQ62hKXE4tJPCWSr
GfSmIexD6SIR5uvBZ+mkq0Q/yPcj565vvwI1Y8aNv5Av/Qr8yl7Ph1AX8MmnDr/VxD2GZBr41O6s
HmHRhAJ9r8r/A0C0fOcv/W4VgGmawHP4Bvo3zvGXHb6DeKjFNfQPIdAvHIpQa+H8BKWXRjmDIAC9
1hjKCbrFGsMaA4wBG82ZxxPeHN59wZNMsB2UyUZQhrf0oNJZzU+8lGPifBjL79vrWj7GRRwmAUsj
53QmyL/9ntZ6HjWgm4lkGl7Y7TcEOttWi9/aYUFBlHbda/m92RxG5ABPzGfvwCX6Fi8BHKfzakfW
zOlDrftnDskCix+oNLP39awqN8H9smzHf362mxlUKbXB/09lNuxYWs+ASB2rNJzGW4SDGBKwagCe
dVuarGb10qCCVAz+k/VZQk3hONJzgXeJFDtNW0r0q8EKwr4NaazdWeqGyn9tRbgEfddmaiLZwqhF
jpLP42p/GPtwnKK1ydq71PTfnXoryO3sDiOBHHpngUK+Ge85uf8iM3GXDCfcNCygA/eEezzazffh
c3hPdgwo3CdIY8vr10+JkmiiBLVogTUO2BlSOuhZCDXk7lrcs5l8uECSycrtdgXfgK2YktTmC+Mp
mSHxneRRsUUdjGUsmHOPB8nPWOtLMLFHobLbJWdobA74PNYD8hqsjR/ReZyd5IahYsvxvi0ipF2Y
F99g+h/Ml+QFCikUqtxpHKtkHzI6hbc1s5n+xMBURCcKCFNC3vIfY2p+CNi99kIEJOQqPPZc1z2H
O3Dwx0F07JYVTWz/82+kz25HF9/PbGX77Ow/m0pbxTaVNAAQwjQtrb7tDXQ13O5oHGN64Yyxusfw
unMa7zop437UcSsQJXpOIlQ3Cn0Djxjr/V1VC36TG+o1yD51V5O2ahJxVHSv09YJ8fzxv976XGre
wXBVe/Ivv9aXuPZXMVgg0cw1aneEgzNS5UuZkUAU3QiN77OnguQ5PLZFDVN6lh1YDJA7DkYfFSI8
gQUe0vAaDnMgoVB77hn/96zXsAW3dzvzvshZ0+hAMbwM35DIwlWjmyElkAp2RAhbuv39D5k9mVA4
uZhVT4eLaaBFA8QRDWq0cu2+WpRsd9wghwIIsgWBYqKxJm7D6GGrKQsHBFRQ2Yd9sN7bkGuORMwZ
PJ71DpjyeVEizKSzgGyPgLECVEBN55lPrWHe3DjRyWbZJoBlGBW9g4FWwnbIWHTUBv6BYX4KYA2/
9u+e3cYgDjovwpMQBu1ww59Xk4zDR/3y0Vg6OHcxh8kfDffwkxmT89WXnUECDy7UEp4GVchc17bf
vllt4KoBpQ7tPq7jll1R+OGIdrhH3mhKtvAXnjhsn05zriGcd3DPSNL7+Vtrdm0CHHCH9jGzfy0t
0akVGjLJMJM8cV/cuvnW6ThEGuBsLHMNE2Tevn0e5gd1jMGdqg/9pX2O3PmpnIi6qko7mYB/Nsjt
nY0MSk8HfkXybiWUjOCu1M3/mgnIZSEK8UJBxyI8EqHoQ5Xd5AoWKNnwfI0FEQoONqiE7DGKvL01
W8q8hhVp/+veBxagn5rTW1Dt/HyXmRf+qg58nTxuEueWHAmqDsAk0Q1CgAKezwWvDbPLklFTcrnb
+bywggU5hzPvuumqjvFZvitCFFreEq5eAH6uSlF2bl8RdA6Dc5OxMyUO4JlguPCyMf90ASPhV6N0
0Twpj7tAs8fdWZ7aM7j93byp+18B5aE+YlVBFSh14YYcUU33glMf7A6SWVrnJfes/uAnWdb8huG7
9tBwL8f4vVlhev6iG+M1OGraQVuOn35+k9hGfm0N+Ra+Vyhak1Z5nfic++xqoyaU2cxSUiIL57Os
EdPAdZ+iEp2kkuybAMc9Wgma6KdE4CdSaPVpNxLTUqSRzO7BT+XFmsIgjxYNicmjNZCvchjR0Akq
IQ9u2xDu7EskB4ABeui984qrYqvtd4nuhC2jZzJUWvcO1hiol09zr1qASc7F46Wfcsz00caq6lqs
hpaME7pkKT5W9uSt31Cu4NHVbSDXt4d5ebPDis0FxdvmbVhe9QlFiRJRTN2S5mBT1hVCuEE8ms+Z
PeUi1dQfRmJqlqXsdJE3RMiiKpkzu03RuCeUF1xJSx95tpEkL/YZzwY7IPzQTnp/rO8EAGrGqkRm
S7sGhdzd1LcPzmMoQRNo5qYRk9amXODTTWM2jWAohKMIKhAiNXQh3Rmm6t4kDkvSe2w6u5a/Nhhc
WiZSce/3TJ6hZhoCKQHNlCBV4terPcgw8Oojy7FkGWvN4KA/ZW9LO93RxC5At4v8XtOvquzrThYb
Tlx3o0MTAJFyWsHayN4at8KyJ8tf+3VnnhUZ4605NJApPXVLqqXK31MMdQ6GPzHEGEuv8J5QFebV
gxrngAZXlikk7cPfLowRQhoa1qvravRy11LboXxcsBXPmXUC7gbqjJfdG8wIyLeWElsw7uEBUMD9
CYxWq6syWVCvnD6z7AE8liOZNXPZhHGt5jojoOQpcCwBVeoRohfUGxSzWG1O25PAr+InrGVh4o1S
6RbpOmfkf/Kf9LLaucE1cMLwSh/zQdvuQJInDyfXu5q/qOaHyR0L1wgUcaER9fIR5/BiyUZTKd0Z
e96KTw/Cw3xJxGqp1lOMJPcx3W23OQGexPBAkeMuhjFn3Qi9/zxREppzSCZS0Qs7cZckF+seejxK
G3PhUhndobOCVLmj/aHM3naTphV31u1FiWwc8WjYwSinwN/TRLZFrLDmRXkHw2bKKnX8qslfscc5
6yaBAwMItyQecrsB0H40sW1n8lLam9fM/EKGYp7SYLRZcdmPydKe5CakwReJAD+0WVhvtEFr+nuO
4hh8lYhTudxuubJToZlMYpv3jMR2HzOCO5R8bzN62p8d8GNBIHow/3XzPws5PPmyemAru0MQWrWm
2mOiT/sB4EBYkPyxwIftF9AhvUCdtBVThyIYqOtWqnWx7l/aKBBXoRA6eJ4aRCDytaHE877mPiMW
3TusWBeA2n0sJy4dGBHAcT8FnZ1idvedwRfErZ+/XfWTo8MLf1Np5cGUX4IG1NCffxIdt6D0tZmR
O/d/K9+4BHTfoAHnanQy5mrYw+YlGlL2RSah/UtwZgPUuLpxrxDXW4fKwJGs2XK93kVM1ydUxgbB
j9DwSoEtzDn/Y5LO8a5RH1Wozpy2KWhvOjYLCT3t/T8xGC7YMS7/3uUHH/m3H7T7jrSyA+1Ol9nP
xP1CMCsbzekYXs5RrknC0n+PZCsl3Fh857oZNYf2Wzd0b5/X2dpHLbIJoCMgc2qwMVEvHTTl81vn
ANCSXVusevDjRHm3I7UhGjWpLUxdd8BDfG3JeueUhK7gqVLmD9c60whZHqYGlBzLDyGOUumnNwyW
AMM6BeJGYPNnRHHGA+pJGg7ZAGFxGR+mobMLrtxcvUZ5JAwzIryNuU/1voJYX1hTudMPS+wJzcUv
OPXFOQwNukJhLrGL+xl9Yn+Pylyc0MULL+bC/cZkdX2XDoRHtiGDfiU4hOFvaxp4f6yCrmIo5RqP
VUl0lonlaNxHaR9B3DTaaaY+3R0NjUjjxoh3tjffMaqgrCDoRKwbq+ksfpxWn4gStDYVsjB3aofg
jrOnKk25LGxos0BgSeV4ye72AzUHFjke66UNamwZuj3BA/q18EYhaX6xHYuFCgR9WTWzuPkVrDdn
w+76GIkVD9fPYuPRCRyjHcaMfkblq6IelroA3PfgYzKstH6IQegRohnmk3ZEUkAAJwZiwrqafmM4
/IUEAFN2bcWgXQpgiNczH9aQfya89m+qfp5qXLFjRB7I1vYS5x/I3JbhMwbgf7cyPnwkWTFgU0kN
hL9H+l2Sh0L3T3tYjm33DukFWo0dBs3MUXeh4ByoZAcEiPcf1S3XBeRZ85eNqCJ04PDAEsvu+X7W
PfbRCeteU147Lt/yRPMuzGatd75A8yixQE8ao5pp9tqhKK4CyFyoRtXDbcJ21gSze9O8cpVkLF2o
tR8Xq64ZZLtPhHReMmfd+6c+VuqLImbTGnezWrrPKhBV3JXinbb7CZ4iiGFO6GanHyrkyXnY+c3X
1gz1vkgT+J8U6z1GpCFZihApZR5Gk5Y7QWH5hrWQQSgV3gYv7ZA3X5VvFU6VKGL9of20/dprWlQU
lihZ6vs5ZxsvMucNiznDGo0piGygcIlLGp2ui1LUKu+Lhow0s5qykh82Jw/sP43RTAmJFy0XXlLK
BXYPadgsXr19Kt/R0BIm0VvFWBRYO9gsduZ5UIBaAEohes9kyyvGRDQ0KmjTW+1vkuKeQq6VJ94W
XEE0nBxoClIsiKp8zU9SNv1PYq2d1+Ps5PH7DwHOuKzVA98WmyA4DsGoQ/u1rmiQwhXjxdSut/Gc
awlNYwtAGGGeNovnjF3CY+zHALSqa2/8mnAoMLPkfHCudeYCqR1pUEJmjGEHJdQhHba5nHsZAs9y
zxe4ZZCDCLmV/vHsALB5Vd16Bl0CIc+PG/w2oYwsvDKW+8vahwwzd5rJt5Djt6ftXSZsto5RnZPT
kMXqvqHRc75b6BlczvNBrUsT4owc5TZ/YCuC4arcdJNmHwvLyw2zIfGTsCpO+WB93ekgsjK85fuX
n6AuBp3zIy8GYGDEc7T1W+VQ7thDTyRzXkASxeXeMxFSIQXoeY/xtB/jnTkNKXHQXhuq2MyrY6CT
FvnsM31pii/i77I9CYJK2PXzeNX3MIxCYICNH8kMm8h45xWCaiNT+4Ny2YR637tcSAXftFVuAeCU
2qYZ9zfW3XD5Z+6iJWtkFYTl266dS5u3RRydekDFo1vDplHCkoUb0rKLleBnXQ2owLPEJXvYHnCC
doYJv5PEpb4QohY7b5H0W3TWN0GJXb2kZ1K3Pb9U0U14c4bxMerJT1kh/WQQwLARISKINQO5y7FB
K1YTdH4SSm8pqYnBJ5vNevnTxKbHMVtqB/9trLgZTlWeu/gPvWPemu5/jR6vcZoeHhqGxahPLLKi
lplD95AYIsNjYuFBL8lnTxxJ68bOm1wCw/Q/Tq5WzIdNyMxhOW+fdoNdzm69snuhWQsiw/1Wyaso
3Z6pGZm8q/uKDrdV9wdX2P0yCHclaie9TpUn45ykFSFE5+TJ7zKzkvULUtrqiErXhDnjCg4BAKNo
UUf2mbG8HxXhwALZwBkpzB9UbzSfXtSf5y8gMcQ07zarJH+xW3YRmMUEatUD6KXvHYNar69cYybc
nCMHOrZn0cAfwOEO4itokUtIOv9e9R+R6+s4KyRjdvLmWvIwc8RzNnHjsh9NwUz3ZKFrjEUGaDxK
XpOzCMCKYOKvRJSaVDBO1nswXYsMVsn3x9kOmCXr2HnXvCYDghyI8giQ1caqQ+1TbyTldbtfNADT
Km77Eou2EvpP8WrYzTUjJwzG2DELtym71XwQVlnPH/FKxrWUuXtlo2sNT2NleynUsLUrqCnLCK7s
Kv22rOnC2R6Gq5QEsWlX64Ea28CemBy+gk0NCKTOs4IBoPzYG6v40pr5rPpYtqI0m8hXNIs8aPYL
i8hc9W30UlPNhW2XM0/DN1mZjIjvwXePyP8FdwFwOwzyevimBU8UZMArdb4fBiGV/zunf6PTmJN6
gSVXQaMh93a7mX5MVUKjVB4lJExbbesNjNJTFADhbiCJiWGdTSwdGZkM6DY+1mHbjTvRmb/aetPe
2/uB+C5KYlaItAxJf5iK4YzgmSOjg7ZoiP7twC/k9I+3BNCuwezOnDt33wAdtVzjp0rJAm11bBXW
DDrhEjwB/qD8UGDEUPh6L1EXkEEz22+uvs7d6yx40R6lPiv0UfFRgi41BlGX28u3wWKJjtMlyRRm
WGVV/YFm+f3Wu6t3thUmL6tQfOUtvp6K6cFddfyerglsfP1YJXncwruRmBIG+52egr/s9IytOlcs
Or0qZLQ2N9jEK+jsADkP23MtbB1dVIprYWNqpdEtrbqfFIiuYtbCeMcfd2Gd2C2vMLB+vCYTtVOw
rKLXjxjF27Dgtli0H8U6TiKVikzwMR4Jm73wcK5exVvcU5m7Bp111L93r289Ze3P7opw4rEFaVgc
Du2R0sswRaSHcqw93TuNVYyP1733WP7MxbsCaocbDlQBA53ndkAHtj0gGd1fdfpIor+hhq/f5Rrs
9ne/FtofCrVnIONsV/xxeltdhZQcHX9zIuiazKh8uHA/nb/ozyPM5VhW3uBvN16mGzehfgFXvb21
iSz+cemlKA5oaUoEE+2SDyoHwckVu08KRQGl5kCwmobkxXVAsj2vQXd909Wqojk/xnhGdfIjPHzr
6+u0Cm70thhnDR4fwbKOq8eVOAXVftSu+L+qPm3ybof+0BP7QOEaK7zM1QwKEylqFoZWTJU0sNId
M+2ow8aOmG0XJud27i5j8beruu4pNx5dcSxlC0zxAGxfAHmFFsAHL94h/oAZBdPmKJEL7ZLqS22t
L+L9bcXKqXVgu0TExmUceG5dnqkKyWGUkwP0lyeweDLTlKcDc3twfTiP7GXYVtkV+BTCIkET1WWj
Xenj2O6bVTwmp/9V/v0G/INvt8C4HN7X56eAORqv5rc3+j431i9AQcya2/bIXZiFJ8+Us7URbCCA
eq8vVtCdLNV19JRGJocqBHfCeHFCIIZoVP9YLJo+VtDI8BSaZ8EOTkp9OFczZ44CJJaLtTHll/m2
LgnfqBJEdN08PvLChPKGC1lAcn63/ANSxiE4Yo7c/VeDj5TDBLaI4fj+PqA0mYVZlb4CBxzSBM1+
FUBWcE0BUvcrdeEpnU8OMUEFR9xNgZzX0iEkF4KpGD92EWmluqe/usAt1QvzW8VSaXe6lp5R8EXZ
L5DKZAecv8Z3PFi2UZNPy1iTvYTh8hHOlVhpTQ4p48YBswp9ahisnBIdELcjAvuPNVIIuzMG895o
55BI0lJ/U/0EBuvZnJNhrs7KOYx+zWSRTT8Yxy3Ylyhsm1LdHq77bf1gKNyJTuZyUH4BidkILmxD
brqxTSQdPCDM26+hONVDEtXMzrZAD5YVoUV46ASS1dLMVQ/vJgeLgoO6E5+DPvcYCbAisheHQgym
TEiRLbjvlwDSITlSx6mqH/2iNQWiArkSukSKqHLDkvcOck7o7AfWrwjRZyUtLyTL3TMxLUtC0+l4
iifMYfnultI/w0JQfmjJqYga9m2oHweDU9FVtL/bn6alPdqx+Dfr3TPJiuEVW8AlGRgxDicqJOBX
blacKiqnH5nOknShV0KEqV9wu0Zvtu/H1dz8ypTAyiemtQCDnBPcUGcO9CbVtZtltRMLQYv7booU
kj1kuGvx6ucZAuXHydAJQbj2Zfhq+X7KPYsa/HIOqHmqqFS0vBz1I5/qA1lMWbphOY7jiZuF6lZ8
xNZSyR0OjKJAOUmYqD7gqDCedTgxv27UFugF9SVq/8bLblMYnk4Y/QTfo7SoJSxibCGKMe2BhjHG
00lVaIg5FUMy6xSnunS6LTbCrXhc9d97Kb9ly6OJsMujK8opqXPxbxwoQl5upSippxtnRsq5kJPr
jEgbzKNLEEYNy4y0U9fRI6PVFz2v9YUKoGsnISHA4NehvThWNVH5LRN68CdN/Hmc4ZvnjTqY7a0f
TsH7UUU4hP+43r00zvHNpEuwYL5NkPmGWjD9kNICPkB9DksBr/fx0X59/ZQIJJMM/XOnwm51+rG3
BG3XO8oKApzDtam0rspHHHQHPa27TVRO89kGAPrK6gGkVYZaSJHnwdhvSG5M2sLCvlLwrnyHga+z
Un7ypVVznD4m2SsBso7sgZPb89Q+7Zg8WL1ValhdyVAvWy/JoThFcprxvZr8wVFJQlj/9idbf5kV
MsyNkI6jisd0Q8dWGpHsmPaeWCkZ1+wGPKmQ2hl0vfunS2/cuefBK/ElEOaICgAN65NwC/9b/MKU
8WzJwvMoNheHxbuZWltr2IMXXGqEC16NXgW09GvNAtr0/HTAj5C+5Gd94dgr8ur6FYEyIHITnAFU
wa6T8lD7TwDDnRqJTHcPzN/ZTyZCqpm3H8tB8O26MrBfGqN1lRviDxzDAGADxgBVbLq6guvSNjzu
/45sDUeOcNZGL2pNVuMtpkj2wABzXnLaiihViA/8VB3uv3aOuwU06taigPJrbVUm5maYW4VTjL0s
J5kIef21dOoWGu1UBGPjRy/8zG3qMirhPR5IoermZixDPLLxiYwoDHfZqmqJk5hAvktOLppwz/YB
SzpwUxRnPQpleGHJjyiQRZkzdMoC1WH5wRPtLzF/+5mqrPfj5ZJzXeig9eAaqEkVgTw7IhMgvZtp
7kVSu29hF9nTazd5xVrLzj0WKy791z8NuyFnrqTMs+VamwXrW8OHBRu7Szg+Rb0Iu2tCuf4fvu60
OT3I7vecI+ytyQrlL+OVnm6WYZnQSXUWwo9WPW1Ba1WOXiK6wavfDoUsQcjX/Dva6wt3rZ1OXX/s
BDLevQtXTCkSHyZtS9MSmPhjIYfFqkrZRAXMXuv0FhfPYi3Sog+/0LmFMPXMO6L3teugHwnJ3kqI
1S0t8/9U8IUaVL/6BAXKA08SYKmOJC12S4h71a4pJ1pG5K0QyAycVeXe8Gs8t/14/63KqgRtobav
FT+Og11ldesdwQ9vME949TT4a/NTidgyga0fP3aeeXKEqlXRbtHYEQsKIOvvOeBQeLvCiQ4PF3VR
PEl5tLATqPOyFuIOxFMm6hI/pqtF9gTnOHYYIUYKu88FK3Zn8FVbxLcNkQEL8Z0Paerzc0G5qFG3
2KIXsvRo/Ntrp8sxu/DF1rQ74ql6QFhbpPqxNyHXNQgm9hw1ldFd/q7k4WGfc4zUPe1QWz3S08C/
mTPBBaTMddh/sb19H4VC+Qrya7jpJddnufkssKX3tys3Fy592gsbEuMcRyebunstUgCcqzAuolAU
Cm1I/XktzegYNNTUOA+BvdC5ieADG/r8mnGx+etdC0SHrHTshAeYsGRv24wadKe3GHXhcy2BKSYR
N7OGhG0qScbtfTmhtDzzllfIOXFpw6GNmoAsqaCLC4fjnfWmcgU9jrLA2HVBu4tUcgx7zxqjf74e
fc1fZ9pXlu+QMdaMCdy4NtRg8tAMuf7CdDuTbEpUyLhddaC9gJ4ke+pe8Mm5hHg9BXu/IAb7R/ZB
pMWSucrUZP0HEUCWoVd94wy0JMNeBM5KGmf7MiWxp+I0OCaxK9Fw3Dl5CpO1u3xA/EiB7E1GcIg5
XWb0PTXZdr+pmMNIBrtuCQ0YHed7ZVw3xdWSaB19N9HBLaaxD08ntR4GfhvEniLly+UvuGR06Na+
lv/kRQV2beFmx6jwMHeJ3Dm4hWW6r0GdpPWlI92gI9VdnSQacMEkggAG4BtqCkobO33H7f4NsDxz
yU8TxCXTooNkdkOE14KwYUdJcphjFEOe3M+tCiE10CiiPMnjc6JrLVIPGrwp/OyQbcvjX9fH9WS9
Nb0FwkKBzZbwwKKi1zR2Q9bZhaYkMO+LWZdekRyedccqwQ4MCxqlqvqBaigcH4Y8zDbAe0jjxeFM
hkN0ebzDoLLqYfGadKRiIvOtYTEphvRmePAR7vv0Kbj9wP2xMt5ra7X5kVT8HsktM6InuYQvPyda
exICRqt1enr11XBit44j6FC0q7tBfBgTVCzcBKhUwxYA7CjZbuQimUeYjLhlMCvwtPn1ZeITe+b/
VOcLoSX9GfPsjxLxZUVRIAwn4zd8A/Cn30DpUNmhynGJS9KTT/o5ySApLd/9EkJQFjgjhDTT8WOp
LXKBSDUOa1x/vDuoeVlDa8uwD/iZC7m2jgs+a0PqZwBLB0wiuMCBxe3zwenrVpRNSwBXTqACoTzl
2cNpGUOi5EL+olLoQAtVLUgd18ruGskPCVePTMss4UIIMue300qhnvs2/PpTzB4au4ZDu8ZnZj4m
+9ezz1EIqJzqnlYBjBGNTWJYbvqG5BbKjOHy+iG5ozFLIAhf2ZIbwFTNNdW7EGh7uzMWpF6jnDmK
9B036ylGqX6LCBuy9G23kodt6z+xbc4MjvH+ZiV28j72GN110ILJFyzh0oGhGXWIrkDGTyNgaoUE
vogZoqFAxjIQsqWnKgHu1OH+a/azE5/poBAF9uHM+VFrsoMxtuwl51vEABL+ryIPPHqIJJGjqZUk
c7as7kLbh1JrPhNIfdT1ZEmzl6wrcJy2Ml/SoiBkeSctBtIjAJs/0cmk2DAOdw7lvDRXmhkAkhUB
LcocHvyZ3M9ZNKpsZw+/iLfLzdEC47WN7nKvU+pNZBKqAmn/WM9Jtpyt6ioETK89y02rKZwpKIAS
7zeB4qs9N2Rabc8VhWcZq1cBD6G7Uot2Xq755cBJ2fB/0+f+UBvjUbTLG3OCGYb9hViQ3NVjFiVR
fj3uMEdLwMGwHKPMzkPIS02ZkTJPbFeY7+gaIQ8tQCTa+YohMXpUD8k05GAy+Zw4hntcGdcICeMF
atRZwXcsqgwlxOHyxRPR+gYhmqRBqa9tq1HqYu+WLo129grf95mSysSLO+4yOf8E0EFOb7Ub3Ljo
1BCPSMbpCA/WKRaRNYGimLJWMOI3WZ87VGhRjPE1j7joIjBWVg/bA/XSEHu3rKq4ccoMUe7nrn1D
iblcmEy7hi8CBS5IxhxaxQNhrfiPkcPWcwKOyjme+3fiaQP4MDmUYt8YaKmTmjlRZPPeKPcBlYK0
QYpodsZgxv/FuPL42qJY9583QfAp3L3JM/cbSVyPQkFG9TJIVu377YrxOL9iWrfCgYdSlrJB4TDH
oXi7ATvPawvNlKSRr/CItWFg8MYp1+bo08aqi+Ae7gy4RxERdAcGdtyshA2C7pgxhmPlhxIW6N+9
t3QPJKvOPWQys59fT/8LX0mJ4cB/0Oc4/U0qCQtxs4aHtRrzSj7y3QlDmMiPPBFw1dfxvu1Sh1rX
MCmYNRz/VROSQrRhprwz6aX4IXnAej0J/HYbgVBylDotJ6seJCMxaFu2bm+RRg4DQP+f+ySN+3vv
C1E/tHhBP/BJ3eAm+RQHL2t3rFsVz8UZHh7iz/35SZ/D2kIO/gvcX3ijT61M9sVNBC+FnfuYecEJ
iewyOaMQU7FDSUO0dD5dvrExKefkGn6ijNxzQKpsa+inATsHoW/FeSCb4mZx/9euMtYvqOxnCXQw
HZnCVwivC0S8/you86QZ2UPKPXZWq+O2cdPK5oSIWJu5qSoLXDBOlR2iV0AQyhyvLsw6a1ageszu
p89QgEDr0dlF36Vcg9gOTAnSwr7uxPYRWqRfGQstRzXn8In+Spp+hhbZ4V65R+w/iQ+NsXMeCii5
W2QVnQeoV6gPPABpYM6tIh4koynexLnyODGwYW9NyPx+R4RbV2GjRsaC4LwVQ/RVqxNWP4wsWjYS
GvlT93xMH7w9kxDu22HQC2Vub03gN2uz3FQPshP60Nt5DW3FUwcX1ZFhDBeU7yTUHGB0DHBbZYDQ
WJs0pM5rlxqHxB1IPO6cw+w7s19DIkdNCfeQ/OfM5jH7ziY9vbJBphH76u6jrdTDwieSbpyQ4jrA
3LGh89P9NAAhT3Z70tXKvWoV82vPQTZvLY52xwysKF3lWU4QorXX+YmcTBhp3yU/Oirzt4jDY2mm
/WmxigU3oFsIZ07AImb09EXmmltFSDecN7q6V4seXR1+ZO9KNcfF0i21rNqFpiAbpXA0vsw/jv98
q5Opv04fUxRBndfjVtBoQfXKJpvgspaTC6DhwTE70Rc5yehEZZHJGdrk8vYWWVx5PfM1zF+fBqAF
uduksEcLFUeq8j7JyALuC+0EUTalv5LLCXyV12QJzRF1cqdXEPxBvQXYRbzfAFCQcZuD3Ctq/d4W
CXIX16vbnkm3Q0GQu/8pP2LPjOAjhRsVFqOkGIYN1VKgqcPZslxUOxhAuIuL9NgcGsAgzz7u3KYB
hyVQ20ufobgl90zvh5ALYHvhcnEK4zXXXJcOsah9FTIDdpYw2DPrR4YHM3RLVFMNUQJ9OAnBDAMC
kGOIcMFiS+nlO/TO2tKwiuEc5tEU7/lLtQnrA6cdq6HFN8dQzhBvNJK8HbAtKcQTCsDKKBFP8u9L
lACgraWTYN88StdkPKcQ/NqejlAsDT6mFJ79HJyP6f4EQCFsiNc7SHsHsm/1Q3U4jPQFeCqPl29d
DURCSstl9T860od8rA22yIYkT9IdjpvzqwjIw+/UvJ4qep71hi9tvHvKREJBnwMNxVGCK8QS/Hsl
BEZJYfYdPwTy4rORg68FsnLN/QMkrdlti1L1TztQCWit+6pugAXGiu42ziAurkPK+7lvJXg67XhS
Ppl2YqwKn3uNUm6RO2u0jcpcuE9GNhUjQGoarwaqQk/3ujkJXVdeu5eew4fRTi0N38nrKpf+HJJy
ns6HueD8XVkOiZygfe2vEGm3SgtfqGZFVkw+JBLQx7PGdrETONeZn2119krFmL3jU40S0db1Jy/M
ivL9b3g8PVeS/c1pSS8e1JHgqO/61qwIsAarC1MYbbaS8RQBkMEsvg2PXc5K8PkjPGhKkvAgX8Xf
h0NUriJqINqkTsgaxaJdkxdwSMsB7yUZscgffs9xfbrJoV0pYUqy4eIRzXv7qYr5kgYqDtVCmX1l
1X7nMQFd67Q1zWw/BfGPqBRrfD2KCmUC+KL7v+9DYvaggmx0YCDYTcJ87L78JFLqAAtQwc03ilnw
X0PJ3hUUpUsF1twflM++K0Mpqv7zfMzfnIVOJw0eLMIuJRom0i2JzVYndUX4O8It9OMbDWjRLIhh
V7rMAqzWAPIvT6Z8OmdC5kgt+GTxW37rGPyojeYT6Hds9+oqBHG+n/F1xJnXKu0dqff2UkN/Zy2W
SfLNnwVkUsRiP0aMxcQFvYEffpT6DF6iXB9fyzkt5PXSmWO7pj+udwDaeeYSulTPva6+vv+KrvGw
CISnVFBniLVLbngqSDUqUOFAjn3mmNlYjgqOAwtCmdXQD343LUbMcO4YQZsFSuy6WH5fg57hrpfN
wcvX1Ygzx6gRhZJILYPrZVwJqcSz97MWE6DvbPv2DRxXzgu7i0VAM3pQGA9lFIyzpT+TJuqyzxlm
zA4VjEEAbAQX/gy8kfP2F1h40fQSa7DbcFki1+4C+XmcxkBEqXT2gshkcAh+/A+uWnMCi5ecvDx7
p/YASN7nYUqBQB7ekoec98FJqbkuOemo12oBKcJO/avxuTy8rwBoPoUw93rPbAkYDMQsRcc4JeR5
/0tzSlGX8IaLtdna8ASL3UESy7fAaISK7k6+KsEySJv+W9ppnhuQHT4s9H06jDPESVXw5e7I1/t7
k5mMahC8xqf42f56c1uSPQGW+uZk2tIo5BnXWLozf9EMQaIvb6GqhRBcQHU4/Xsi3a6AA8UcdtdK
kHKOXmuUD0GuqJZlS36lN2bSbpNlj2lj9iw2NcFDoIIjtc8pv/E3WG5nyiOW+8qgurKVTtjmlqlN
Nd9vzxXhMONriWHkchcyi4Omzlgv5b1EUhEaIllA6YiqLTE0Z0mpJ3X+3EWUKTcUkM39b1gN4GU/
hlqdwD1apA6TY9COcU3VVlUp76Dn8ZQ/AMmnkurq1ABsYzSYlS+5c4wbbTE5pk5r4bdpqEmceRKW
moHe2L4LGfhuMT2BaCl6V4URC6X7rjqAMtblFUF10vDON+Ze6nig7X3ceoC0PnvKzRFy4R637IsF
J9X518S8Oyhar3Oej1IHvp3Z9LH1FdC31QFGeMwOq+Mr6ij+pefieDfpbXr6e2t+HfFndjTxS3gA
1R/oIF8cNywLGxixp+n3ZbpsAbXRKMMgJuB1JLPgGGOlWSCim+Ui7szpxTFeUvwCKoXGebfii/hT
fHFx9Oz3EkyLV3CPkzXX7fo9ZnVde8k8eoL++3oQRtHh9pBUzyHg0T2AaxSR4h+eAOJuTtgKdW7p
DzVJH4UrcWzB9L+sPh9pcMKohAQKJQ+tB1uNiYqQ7i9JblKWDJqmMoPtpA9fo7rPCULZ5vi468a6
jeHP/bsvtPcTJVr9Pjt0m0wVvMi+ICcfjMakeFQJr1rtoPiqJzJW/TQ95M+PcJ1E8U0/jtPq+QdZ
uCll7sgzC+rJf9fB4UIhuUxMUpoHQZbOCGjp/BbpBIlkj1c7XD/7i6IiSAKKJyINY/7WvGqkz/U+
N8ycxWJKeDk5HxzPrVj0PZnJbQ8aS3KV8dqapzoGfRWuyx4NlYFvm1PgDcx0rArfvLnIDas2kFyt
ybycJGJLtSXKOa8YqWiZo7ePExtxJT2rDyfe/cxPhiSwwKpl1jCeyKfxsl1SOANY22NVdSI1MZ6q
SSfGzZukqOrgPGbTFvp18xMbMd33i90z3VLzH+kdFfn5xNnz3ym7wK1mixBtiihlLm8GHmmsmi/2
6aWQauRRlZ/tr9hYsmwsHK1VKiDiPwB6scMdLDntlZf2ZHUrQTqMhXLZpdOkfdz+ioBFN4/WisGP
f8hVYAOuoYGP/ofcWjXDeskT8o82g5rb+Z3DLvlPh+I2r8YuJSZizvh9HTg7N3XfrKdPQflNHIme
SjrMbrOL6HF6bp0IJDFvGoSmh4WxvNIUTEHEhTWWUW49Z1ErD7IBLeZnxtjZ7gdKeYgLRhVR5DHE
lOuJb+6raq4ycm3GW2PPFR5JPs0W+Q8koijzDrhULtX9fr8v7N/Jr+nX4AH/Qiwj+ohXEsO9hemG
KjrfE2Mam207WJq8ItJv0Vax9mj47O2BiER86amLtNXzAZX35I0qri6HAThoOK4SQ9SYBToTP47M
S80UJ15DEe4KNcpNmQC2ZOMHYTH3n12G44qZQUm88xPKnP+OJUGtyvR+osjjYevewrjhJaPzRBh4
VWw1KT3cEtgeOa7LBEg3kyxk9aJyUFS5zKRj58Mb6ThwPC5JNt5W+D/BNQjO9ycBqIJCiiOIauoW
80ts7FvEjZ7IUfGrzGmtnZfbJ25INwSarWCJNyW3e2L1Tb/FM3SxBddzatJN+HGHQxWBj4tq9Ga1
9lR3fQ95EhSQ5BdXAeqQYdpM21HpfgQOKjvowHdR+94QeGRsNxQyqTpKVKRPdPxMMdKYqCEUWWVm
uIV8mEhJAXJRAEfKou/cFrrczsRw9C8NUyJkJ/dENlp5nauPNYUEfI4k5b1qYn1AC3ydwSJ9o71A
4WZ3LMwAEpkcPXGrWvjGUnCO0zvMO9LlCdBCaDKQ1pXnOVHqDL3GD/gSNaYzW/1k6x5PcKgOW4mh
o4dMJ3asV1hrq0ZC1yJmLA3YBK9OFrxho4gG8sEoBV0IMOdOPrJpCuOIw7SdOpn7D0KW9unPIp1B
w3zoXIDoZc2mudfh3UVDUkd4Qu2BRL7JrhTV6SVxBKYXtFYG+e/XfR6G31m+meQHTKyzrtUV1o/F
NbvIKICOrbHbNCrS383z92CfiVWOqcKF+rLdbCZ7/j9bqc0dEGHdgJHj3nTbvLsqAE4FrZ5nVyFe
YA3RJ56XmMQzKHhin3BxfRE3R6w1eyRb/ImaivliesQXaQb+CHoCHDUAOYgGRLuH4XWRhWPRt5D7
weNAyswlze5QpBii4G1/IfkZeYvMZRloVlZmWid0HPNQgOgnWgpa7/fxT+T6lJlXBA8Gcesg4MwY
i6j6LWH5fRE7XpG8ZkQX4JMkXsqFeEfncxR6Ni6hqGByI22nJ/9p3Y4pPQsvNDxU1n9gBV+SUjmZ
SzgTPRQQWczTVcZDOi+NgLO6zezEL7yMyJsba8FiBY884DP/ddlgM95iUm8mINJfTJ24sVc7Ec9y
2RrgpG5a/+OZ022TnV0iJuAJUOFxUWTD6rXB8niXHDpne2s1bEbRuAeA9e78J+HfvOAjVZs6Brv9
+B/mLbqNALfSZABSf0rHAvKIDuSTFxRvbRI1+1e8dF9Ky2WsxipjcluqfGQZ2g/LF0gPX54vVsIF
eYrM+Y+jgsre+4B0g1Nk6UBO7kfyZxveYSoWY56OiZgjIVdy+xubPZFrt3pHbLtkeBV+OPjSB/tH
B+apf5c/VQ11RWPycFrv+cTO0Dg1C1d9+JKu3gt2/LAwHs9/ql2gkeJzl/TpTBtsca7zTpDepAul
XuWLz4uK2RR2rfkiYx4uaPF/hS+ODcunza7ok/avZq0YeLO2PWgXl3/CWM1Cpyqi1MEqCmE0lMua
ObbKGaKVVWBtxQPyWklkJqjnEHwQrruvWin1VhAqs6jLUreVp2Zm80EJo+Y0dpfY5SgJHHPGac+U
G+/wMExEBuSDJEIdy3fo6dyn0v/DWLdaK60kBy1TYRbjcnHAdgbhvkbGdWOdgnqB79trrwlQozlC
nkSbXniZZUltCinkMLeZfkdoZn3EBfC7XeZSHy9feIVx2fif8KiE/T0O49NsvFRCRxiU5ivovwHD
JKsv4X96WaIaYyBxuYiLD7WE2RFOKnxOgdVCvz5i2bjFd6U+/wXLyMrPE3h+RDSO2XX20kzYB5gn
zTksSWt2I7IB7pAY3YCzjKROtuMm4VQPNDhijG0YL70SBp0MsUIYRVpu25I/0keo7IJJdUHbm78q
xHg3PGhMOTJiuTDP2e5o1WTuyHTURNzHCj8RWcsRaVSV08Zl0G2t7bvOnf30Ho7qoQHCDRX275rE
eM387V89fcfandHMV2z0Ei2btCRjszstWxCJ+Y9d/Yre9u70BIoMs1zPZa1HizveWMWvmMKaj4k9
Le/0CsfF/EAkh0bnz4dr0K3R6JRQJOIz4c9rnLdkY4fQtRJ6m9+j5+mvNtVNHUy6cyWwkbd4jp7H
AGlhal0ae1zJ1yKYB6QKe5x0IHtnFp3UsZYZo09827q/kZRDkapp7K2BucgaSjikZx6K4m0GZRzL
6yv83cvxCPTzxw3OHFdmslDxnoAXM/5gZiIp676xaFbGmU8WGsoL0zCxep1h7FRCSrjH7xZKhCfL
Z0d8q1tLVC7PEKlm2Bf2YEeQzpPTvbsvNRKyAEp6hySxTJ1a0ay7TEh1gDmKr4lOL1jeAFJQJWxj
d/9XEN5nubbwn4hmoLmhyzo3wgINmLy/jeigC5k88hoU/L/ejOxJgEGeqEIeqkgPRvvidTXyWoze
v0wfn2NREUTx0+AUvkGBt10S7idWSO8WcUPh/AKwzhfNkuPBuo96KMzbu1tt+VyZQuedwQvpjjKI
IgWofCcK9rYOz2VIZ5lVXZ71j1/Qx3V8LZ+vSRteQmO4EF8skh0UcqKnhb2u2SfI9O56qJrOWWBu
uQeGqkUnTs6LDUOFVTMxpV7S83EDC047kdGsL4fspQrSLx3xfcOV8yZ13hIRF0q3w7tZeMDslL+V
U3B+HdZxcEJof/s4VZjKhZHFoVmX84CiYYwTEvqzJgRKUsYI4YjWlaiGmOsWuQVEXlXc10MGQGSl
aufohHIv9o8pLtyCac2htHt1kz7PkGkMl1alR8sFMWAR4sLB1y4KUKP2oNDdCGNyynPvyd2U8YJ3
QCd//CHfgALq6B4z0xJ3fYMc5wTUlwD/b8fwKUkF13BOc+trnkKrmYQgu4nUeApmWLedDxzQmSNG
ncDnuTSJ3r5/jsc7VHNZoDA05myLEg3hSb8Mf7xHqzG0ie6V0Fw29adHqD2iePZ5Us4fg29ozPyh
QstAi3W7FWrFR8g4IlKRV6CS2R+7ll0loXIbwehhopLEqhewtpsOyETyQWPYagnmTHUKsykH5OF0
G6xiJGb4f2wdYY+18/Rns4CY/53qzMEUCcHTNN5CCYwq+kiMNI/p6kZmUXLAMBVrOlv9RrkhrmyD
FnPNbcirIMYaUS1911DEL18zUkdY85rNYod4M9T8f12O/+KCK95Z2vrWYbtGBTznSRjcb09fs26+
yT0l7zVYkQTBHTc5G3wEV8hVVCLGLv2O40sligOT0ovPG2w/5kRSLFehYIi2UFCS2sK21O/gIcve
J2XTlUxa5gjfFMAlTPUugbNhERPaKvCFMmDE+zQ9jnktn2NDGi9eN30f50WKpsZU780CeQlwdz6I
YzCBtdUR3gaxpspCJp6Tor5jjjKInTe7iGyc66yLMReQgPHvT/pFzwP58/4ucfuka5nysqc4nQb7
KOxEwMwvA/1QSF5751PtvThv4B/a9cQMUpQImcGnoh9d2ivL64MqxzHrDRsFdGIhfze6f0JTQT4j
v3O1Pxff0hfLPkcAYCqCjQDzOjdua8w9r+QYyy4QF59tpGnZaKfNDCIe8SPryPI5GoRqzBdj3Aw8
jSbTRenRrl/tRnkXVxRDgtR6+2TDPAjAQCMNcGcjlTqATplsra52AmnTgYJqVnaSqDrv2KSTAENc
Kd5Hsog/7Z+eVeUpz08tQRtQ3UUcdkI7cDFasaCYG8RzOJOTVoPGt9IuWSsDDGSfMYf+FSZJtbkn
2Itql9TuqLjSSdQT5z8EuxGlOWZqSOI1Itnko2wHbMIkKM6bUx25bmhk6FwH13uKji3o2RKrNY/s
sWVfo7Bd/13m/na+e/HWqSgzLtxEhDMCh5BGonFXGAQlaaEOK7EoTSzRJ9OTvjGJoAqJtZgmUY2d
VtBlGbp8cH9wi6sWtYaLZ8XZdbXZw+n6mVYZYp0VK98FiW+JmchVaB7ZkDuBlYwHTGWOC1juE+WA
sIqyDQTMKtaHbydFmcm5K1Uhsx1tozij4uVvcEApsuwYJTCCfMxxri4BLW0J25u44shAewlEsnF5
gBQPZIdbh6BGB54eS4o5UpcmXj5XhNK9ujdwdbMrQDjt4jifh0op6zv6ndsjUmAUVOutGUsusLN9
R4cZDI1aQCpM9PlCb4SLwB79s8joDrxkiX7+3+IgQbmecm8xiqkoEXBUJKLPHQelYnlWr/r7jxMD
0EUS9V5VUmiGwcEvXXLXQlcfFQ//PtDyzMR7QM6JkWmtNjr0Eo7Nv0kVW2i/tmvNUSChHS246xsn
vDkZEnIJ5h0c+f6QvgZ0P3XcL2AU/ycp8F11rpew6opc4J0PHO5g/ZEORItcEBW2aUs9gn9fqlDl
JHNE5Y5tVf+sARu7nDg/fYEpQck6zTZz3iwvmThmtsNjlfAxEu3cx57RA1XTaqGYGSVW95d+Pp6H
J723eAWUT7ZBmVNumRNMj4npiv+V55wMPrVCfp7ABd4E8PTf9AdkrCgKHrX7aowxoUrT4y5DoQmd
KNFjvCCgzSBYO9bzg5ncYIR5pO0GApAoSSfqUGOrNmRU8nLc5BtDoIC8dl076mmz6JxeMCH+jBsm
1sJSAuVFLapTw5p2C5EPXWQM5qc87EGaGChNn5npxrvhXKAl85l9U3boXhaWFYfaa4Fwg7CArgOY
pqH8go0nuaCAsmFoSiErXarMd1gMZE1DW4fE816wThWGrR9xQNgjYNX49cPAamdYJsrNzyUcXzar
fuKB5qihl0YQItt97TwInbnXQHhC4rdAaQKo6/99luWx+psUupqHyQJUvwIMKi+Yr+KhLIxTfMTh
QhyFBFIvb4ygTbrdypzOJtu7RxCav45GZMORpkVkjRIBX3BW4xXduG/O/4fVCU8ayoT3lFg3BJsi
FPtKFfjKm5qeo+jXBmjVCrX3nMAcoA6ID8bbkpQvKUSN7ueSIDsUEBKzfKDm8/ERCThjFKcBHHRG
d/ILXNQtd93ncGQCJTLKG3DtMkMAvSLJ/A5GIJxlVq5PFBLyleNaMm/dFDsSqhvgnyfEB3ZsPUd9
LnFo56ixC/KGsyzV9ka0wrV6poPhU+jZUN6eb4fAHEMJjM4JRGKpdd71P4vqHvNgt6+ugs8dp2Rf
8DFTsMwv0IPXMPudHP5C2OLYQ0LUeHj9Lb4BbKpCZJuymQwyXY/as2yS2ILq+TD6L6QHd1sUF7QV
RuhkuJ+NqheGY5FbK2KLbPPcr+P51/9LpNHx+eZBoqP+t0MeUEGKMbqVm/o632GEuMMaiDl+qOe3
KAPjP45yUqCdtQp5T6J59PxMaO1TPxEEnvGT5E+yO3uaZobt+5KchI8wxZecefr2JogE/5ooxAW7
wFVyMujCCLOk7nDAm8nAi00wdnXV3d8HbUGiFiXGC6fVARGRY/gLbSgBCPZ0xa1pE+RkBDHQqGgN
2ROKO4sEaSmUZa4hacLga5z8QIYofaWI/l+TBj01OsONxgC5hQG5vlFLO/ibOBsJzwtawVTtM2Ye
UVcnha76cIOQQP2UnQLcxgTNk1ZEwvpFYDOeDqODHKvhmxgpNMPPt+39kM1upaolkageZ1+VREVy
WMiNaQH06AWwCKCxgSpOLCduaKygLrqQu6wwTe9rENXxRDaf0baTBUm90XP4HBCEjLqiJ4HgU4cZ
n+GTCvoEC2X79qf+BJAGOhZ8hziM/+XuJNEGyMV7QjEszvIv/VQgvsSLQ2uU1hdHJNGzurdMSVc4
lVxOEFITsuY5o4jmP0yZUSwKFf2VgKZKsM56AFco/mL/cd2uCZxvsbD3Kp1e3robIo4toTepBu09
YundU1bH7kq8YlFCTVlbWaEeJGY96mi3B7TrctowGgfetBu6L5h7O4F1dU4qmrS7MEuekZxOiFu6
/WC2d276RZdDPupdKjUWLys2+GLgtHT8wFkYL+b9/BRmxSnI1/rCVw+nkAyVDgM2KQ1zdwfGCutt
bZsfHjvf+reeaPoEZu3fcdYJun9i9GCPPoRtia8i0Ds5Vw0/FutWAls2t5aGsstgAbJY+rE2fmEJ
7DPK3lkHhE+06Jb+Y3/uCqvSiTosP8J7d77QI3o0ZS2BOXRxy1Lh2r/ilzlw3uvElbFLKU8FH5F4
FJr5Q3iLp0sV73+8/EP+K8TrErI3b5PIlRdLhXbtQv+ZDHpz6S3zjc1Nx3L5v5Ic2RluN0HWJkV4
w25JaeO/OLjB1GBEvcLHlo1ktuDQBRaiaDNAZcm2gGrnvX1WS++4yxb/n1PPcq8d5DjmaDVAEQTX
C4+6UDULWG6KBZABaVIeIyVUMZFPxaRyfgjkmiRN1Js/VAmzM8PgVYK+K54egOkbMlqhXvVRjWnX
kdrel6Aada7cgPXJDtb8Ye6ja+jj9ml7qOlCePKbEXrHPLN7WW2bb5sENVHnFXRklcnsWIQ/R583
dtUaQj7OZXn7MjyAs+zAeDW4gMXe7pzHwbb0/w8x0/Fq17ECvl7nrHUJ22cXm9hoVmnx4hBTS1aH
u99a0Ph7c/VbfvnbSNyrpYU5ahkOrpogZdW1JeKZrV+N0AaCbV+STpFinGf8O0P4Akd6AmAJ1cxU
8K9s030yBmQxis4KQp52NOQnjS1rTGvKg1f3IBrW4IGsQ5iHgmh860VxcVwSFR8iPov9/IlyGunK
f/hzrlGcp/Xt0D/VYLC/C/y1vfOZpDolKJDwBIPcAkoWR6QVtc7sHYvBomBq2CMx0e4CQj8d3505
XQozinjmISj/YpCchHNVLcUDCvBgt00UMM7OpamW+G4hsaUwgRyMTfqzO3gprQgtk93AnzKIzLvG
vDNiNomI3X/SIDWLxaLAMy+7OSuGU4TblZHlzVFKDyclEh6AMEDSJqrtWcPHFvzp6huzbMpihCQo
xDUEd0Or8JuMFBDl3iahSAe5xXDECOVMkLze3y7JkrPV54ayBdFHOi8r5r/jayEj92DqgNca4gkw
Isk2EFmFp+XOCT/kAhoYCdQUIwhWD1QNOXl5tnu6X8ydDE90KPido3Q4JRR1cLkLEAC8BQMUKuy5
VP/ZBeO47/PThqdGLp0IYrbOdO3yN7YQdufGFN/pIiZBScaB0wRLHfmfeQ8W9Qgd9DBbYk0rMaet
kXmuYQIBTTmdONUy+3m/lxD0wWFNCE9+r5xSW5RAoqX1ia96ZeJAHEsXBZmiVW06u+C2h22Z1q56
fmjrHOTyvSiS/lmDNYQUa4TATa1KyhDqlOioR8Y8kadnkARqlGvE2fm9M0jitpCjdOK7BaA25rJP
VrXYzko+iFGjaem8GbZ7xQn9n9SsxmT+mOD5Cr0vvwMikX8jOE2z/eYZwL2kAtAa09Pj22J5p6bx
WiN3Y+aL+3fkJeS4DDuZqNxre3Q1Az/t28eOE2dSReh/OUSb3mWTT0DzxuLtLe3zyE1NTE4/+XTx
FUhZ0oJN4unUydzTqu0p9GeQvJGKkfRkj8EJGeY9alw12ciP8r9vfmq3RuPu5GS6aMKO42ok9p//
Pi1iFwkHQZCEJEawuOdGBvDvYCX8bX7oVb/qGFRv4s/22K4WBqY9o290HgKFbR9FmI1srPyH3hCx
T6Td9B9Ch1+ZwPRQz0rD6nFFFiRB56Juq2xrzXON/CKKCDcjGTqqvvpSESpEV/6u5P4mHm+tjeCq
XMkjjr+LtskqiiaLinYbiiMfzOnzZ7cBOWH1G1MY7WR1W5yULTiyJmTX6xrNUYdwYiTrZ7Th9Bij
ubJeK0PG8raeJf+djocxUrwS8r7Ov6sf2roEnrcta2z1sJicXeHql674LP+PesdnR3JeKv2DEHmS
G7hKtHbQwGB8Dux1666hZ5hYk+tKUP4PyID0/fLirxQNRXSqVDoAig78hjBfF7r28DXW/2RxIhc2
cRy//aM/3b0Ur5xuBP/D955+qrO7iqSZQd4Ze0+QXMSstr7RYOf8p8VEStviEL0nJYf3W/T12YwJ
T0Cp60BdiGAURZXS3+GGmHdmAVxVUiM9aX/Cde7uHUWayfQAxGMPFyjQFxD3H1tFh2hk9fJqwBai
dWZDX2Kbb1IWrmWmbpYJ8bxNCuTtheOx2IO0+sMLLsfeYeOwWghS232UTIq4E0yArwxZ35wgZhlF
fTPSt6znftbIc7iEc6wF8yMSDp+G5QJ5Dz2eDr9esTA+OGhUUO8JuhCXDj/V8xQOabSvbs/1qAgo
+LXe/qPLqZAEkfxOS49brQAiXbxgB3LcFPq35C43Zp/m3nppeWbpIgfBayuQ+FvzPGHANkiCdwT0
NH6rGQKQ9avWt0YjI0IMgZN7vH+3BkY+SPJlRZ1ZDcgmZokV3cnxhQitEWcPpf2h8V2w4RAwUHTe
qmhBU2cTtZpBg2HvqYmLAh9Qoad9tO5+wCa8ZWdjUxrlUV4D6hb9ukCKeSRiO4sf8E43469D3thC
/Qmj5khkMsAvJSjB/FZlaLZ1N1nQflk5ICDRxloUH6Ej1TVko3YgBfeSBZDrFedIR5nYE/bZmZ5j
KoM85w4+dlYzKBFTgLZSzgUVS3bXTc/5gNGLkycmXv/rGR7XiQWt6pTa7xOoapx+RGhNW9ONQwF7
DuliPOJkSPTfkROCMK1jamDf6H4CBvyEVaK/jrf/N4qzP0kiZE/3VI0XDWFDw9QGPDHRw51+6dlp
DXQBFd3GBTxnERraXR8iug4QrR4UT3SBLRL9aQmuCKpUSlwhd6Vg2yxEafcmMqtfuh7Oak/spDNn
jJwY4FaCMA24LxDGqxA8XzlzPLhbWW7xohe8VCqx17EIKNGTh6DhjgZlw9MHkPpz276uiO+ny8Cn
1ASTa2fw+IwtuHN4UpcsOmQlviV4GXdrmgGQ+2TxV6JobC6L5qmtDrx0iZrOYiuz6c4ix8hD6k0t
K2o9/tIFlxrUAGXIuN5MVwcv2XHTE7sQTHWD/9fc41gumc9+anbK4Ir2Ukj/zhaHfsctlm+cYGv5
3Fk7kcJpb0Z4exVaeUOmd7Uv4dukDweMmcUx3Oh0LmgHfSYnSuUFbwIrKYWUgpoo7hqsxQB6QmXj
bgO4DrrfWY8RcnF0Rodc1ToIxMqr2IyVHra1JdZ+tTfhXyfT1wtUiy65dpqM9VqrmUioGJuSn4Ig
/Bg5G/bqr5L9C4occCA1p6lt9yUGU+7iWp+fr2P97HXG4njXBxD3s6disrWYCaDD7WVy7cX1q55r
oIejNdP5eFovEGFMVI/mSxpbMUvaza44oM0YjYaNIYmSqQqr1TSRDn+dHk4ntOVO+pc6F0qQ8ttj
LtsbhxExTqxOmRccB1zbddcfiHC73rpM9h/uneAB66GWUMU0rXs2cfRRhUD30C3tlKFsd+dtQmcj
x+blvofQSBUDXGmq5DwG6iVnupVKRivkYLYRbWbTKSgMXTtujN4tPnXAZ+lQyg820gwij433oaww
uAUtCxQHZRBUtHXDzey4As2sAFvCpFNS5Y5/s0AGQC1NxkjxXdHTHj57KFZ85WPQ3TAQwMqcbEd4
LyjU/QkJI+SxLWEdlIgmLOgBKIbGDo1Iti6ocCIYOaueoe9lvPEtfWFVBXt+EJ0phaloDQU3njuU
8G+13pwwmUGhqUTT1hYQhhifThR8gjSGyItRwGotO28igTavsY1u7TYg1wfpFQ8V+PcPfS9IwdKR
qwGHRi8qH+9HXS8Iv08syVVTMASDA4zJ7uj5LnAUJ0cH5+PNgrQMVAsLdSeddfeX5fIn7U5r8nae
tiHTu0084ZBRa+Axuz5Lf4w4C7AYiGCOOEgE9uuQm3I2p0rlAiPQSNfuWXI4+HP8Ho7FM5mHpBGQ
BmTsqX9Bz1TDiOhiaM+AxDoghIk31tZcvfN4z3YTiins645Jyk8bBkj6qI+PJ2PYFd7NXT6gfr0B
6QVhI4UyWjzl4vKtLo1AQMXyl2tvFVc75dPY/UFEd336PvvTMcTOhkG9z+GlkwwzFABkKQ06v87k
MoS/GJP6ZC4Bnusbz4gEvDo/Q5Jg357OOezVGMg1SUh/2iYNUjT1+N7XVb8SV/6Iww8GSbrwYWqc
B1eVuCKSjAwUFOZo1fV17opfhyVE3gRB9xRpEM4k+3lGS1JepV3ZRgBTVHTI5NzioHjZ9r5KLkoz
hQwz4SR21xvBWkX7puETKigobqWvFDNEw9EsLsUKb0s92DwcIGYSB9Ky7NP11NEQkl86Lzvu08TC
7YzM8fLS4GBo2hZYq8cIOMNHasQYBjeMzco6sjLEKJvAB34Hv2EAiIm5pLSpVTFoxkcXauaxVKEU
PfbHwQNn27ywABT8j4m2T/+N3gh+2N196ikoNS+5X6QeyVSbtC7arfPHfBNrCsthZT4v13aeXSyO
pVw028ECf+ox4SNKfJizNX5tJFke0YUykpnyIRlj9HVWAHArV0p0N1raE0IxHSfKaUV600KvF0yp
VXONbGT+sVqIwo0XMxNjOM2TLX8nkrlNiUbN+KpjY+cG4h0H4SkuDX1TPFfWWbZDNRrqeu/DD78k
lNGydBLVKibDBBIrfTJwqpnMVn1pou6akNp/xLEOwQdYdkEpOukG619YJHemp0qXri/UAWvFIfdz
R9x+ObHXkYyAAoywnkeDaiYF6evLa/TG94M/btrXNWAdBv9o/ew5LFOU097sDkcy8dVKMIjb8Hgg
SzHHkqJkrLvJgC3TeBKCuyHd1jI5thBV1DBCoZAfZItQhB9gjCIib9o5sA+jNmdPN38YE89xAwS1
VfggGSCGbLgxYAApESzjfw7lR1OVg7hpFS/0RYwVB/OBfA0t3G0zkBKsdCWQvyPo+ebfWxhcwjZw
AWFEk+/pRtpaWQO/kAvXuLOIkOS6yHFYef48B3rMuHdr3vr5XFQMzxJOt02jybnSPKvOyEp3AWZF
fQ4ucRHGKOl0HpKaXR+m5LPMIWu37dXa9+koPT9m4XZS582EnjLIW94ewTFg/OshRxmq6Ar80Zfd
0vINdD4/JlFuePbn7vDOyxJFrsGsD7WFXESUEXduKVLNGusRqyjHaUyyvrfAMveEMBk+z9ubpLIQ
XAKZj8NCTVg1zebLQrLbfYBmFxzJPBMfxgo7GT4DdYc8muu7+GuKRz06j6QRoQstAudHZ8CVP0TE
3owafQnk+ke2UhGrj/jmfwbgmbbW1yGQ7MbfICpD6aiYlzq+iI/6Hpx06b56ytK2//ZnIQ53dJW+
6PSlKc7AwY++136edVZDhC3PaIgd6lltHQ2d2iPod3O/ijbMrKa76tAZ46QNZisu5pOJJTBucKpq
essRYO0Som6ER5HVhnjcpFwahyUmGZBsZm8pMx9lrJTpPMCSJjASTg+vropyopFs+HDtpwnqKOL1
ryfsGfFZ1h7xdrJe123qty1dFavlla2QSuHwUdNJ1/G0XaMGWCQTSP5jazeW0U9m0sgFdCbEuIFb
jl3tNTQO6EmM/edUsSzl+zbNWxCVxCcF7FA8dQMTPmgrxxUbOnSNvP2JsB/m3Wv6aEByQOqLTCHN
i+wkx2km8MiGH+MI243lnE7ChoVcZIglAe3pcI+8Dw4i84buFy9ysBCrxxGqXZ5DTHe8WBpC4lyd
X7HeeoK6zAxc6cKCQ1tDir6mHINKSr2jCkvQbLE6/Yp61vVmXmfWlPWesqBvvMEnQjouFUFzI4F3
Ms/v8YoGVJBuliFb+ULwBa3Zw/9mpg4aG2lnFGuTQ7fhG97bQIJ+um+Ki2D5P6A7xVDdwQpvxHK6
7GJcx7tniYOMs8P0joE6rEGi5UR+Ww9svV4bKEw8AAgx3t4DKFYr9EtugEpCeNnhhoFoLtSxWvK+
Zcr92ZGvQSXGZbW1bsHVC9P5W1x6OX2IPMjkknJg6mgennpn7saujVOFxRRy2DfMlCqZhOZE2EWH
VwMbcfnXkSviF1LwGIdBD63oJzX/wMUjdzmrz2Cl6RIlCQbXMsSpIfLW2/CPL9dveck90viKAHCg
KZHaJAtEeRQA3eAcEwMihctUadQPZWxRYNiwB7NWXEV+q+r/MYU6fQN+g2Y7x5Nmizs9qTxbKCoX
H2wdQY72Q715X8D3TF8OmNIk+658Dd4xldoSC52xwHjg+86uVK9LMDmmZX8GM9fkVOXjT92tvkUo
DlG1Dwo7UGGPLO7XxXOihabuW+g9e0sqmMY0m9XDNb1xhQiIgRmeHWhdZIG0N4pf7O+/nhYE+cj+
G3J3UV2Gw5lc3i94nfZsDJbgEmY29nKErzKJFgRaQVrSbpBgo4Fg/z9Unw8+abUush55wXPvxnvn
kg3YRR0aReQ0b5ppBSwD4KDKxUYhksrfzZN7cLCuy3UflodYy9yLmsG9WQQNv474JAr9zZniw46d
o91A4cosSGt7zkhs+XVs1W9MFMzNp8KG4oU7PmlJPzskLrhEB6nUKEubi17JH0o+vTBgBVdn+JY7
rWUP5qhGZ9Z8+9e9JPcdHQbWch4mAHyGeZs+ukqkDPj/ZGS3u8WV9/IbAN+RebhA/uy0ebPVcmwg
wP2z1g0PPvV/A8uXUZAs/LssVlMt1IZxvFpsABggrkNw45f/JJPJRtMN67eHxLnf3vIfwrDXJvkZ
WtlqTfP3lyQ03DQcFa+p84FOz2zNLE4SD4bo7avDU/7deaR6kk2cfdx6dzrpWMuiXap6cC3bUNx7
bygQyJqxjNWgulKq6ZjPGS40AiEmLjlCX5fiM/w2DJoXz4LhT7VOwXhuh4R9E2k2xEV+oFZpbDw7
ygDSfmsqFRXZDyvfh+QHRcHuuRaXoLF7PVkpZ4BN/6nsmH2ejFHsqHZGw1tDDv/peKlfMXKLQ+on
ohGNLZFy5/tPjXm/9qvA+afjH0d09vnE5MDkFWZ8gaHPyDhMtk4jV1sI2ZtzjcCgQTNQChxvO03m
drZx2vHVFnnvxfqp6eFZNGg8wQooJgpBt7Du1qzdSdc+UyX/c024kzFWnpXFdicdqmKYCbos3AKR
xfJGnotGmOqS0yVDTwhiRIAIep3KnoLfaYYfCTdNCUKNL68Up6tcseYaPD8T6cw8SXLPQgcimLU4
V9Af6k6bTR/SzV8XpAoq1+7w5nPXCnLCtC7sEEGUfBU32OvUMk4uN62lpCmpYVqN/oNkw09Fu7o2
LcKerkuNZ6NHhgHmFE3Hn8zwwpZ6TeLrXAajJW2nuhuAIdGCLDAtLPPOZL4V2GRGEnoAfZRL/4q9
kENyqMYpcwut8PRaEBFcsbLPLv8J48e5B7eI1Qa2YeBXCdGWmj7tJlxzYbCupDHfFRV4gVXVVr8A
FbgKWfOj2S5oG+eqXtyuLPxaVOmFAEYcwOMEpvXWPfvyAjgLHCEchR9QY1KPPEU1miZByAI3sb/b
yW9igbu9UIwdiTb/kLm/4EZIdv33RDIaw6N/bHVGI0aohK0wk/64TUiJnCT8iI7O43Zth1fZ+4v/
J060eZngqA+RGsr4C312Iw9myosWRG5mVC2JYWJmHUD/qWvrvInB5pm9nZX5u9dBmajeIONkOxYW
+b2lNsdat18K6BWDN5xzyqwT1e8s5AQ22vadSYPNzn1eLlO5iYjaGbKkA+WNeoVkLzeVAU1mBtbg
s7ljkcM18B/pSvRw5dtX5TkOs5eTv9iJQjVSCcbeTeKnRPui6Hj4QTOubcws4HgCmO1HlYtuDACE
ugfO71U3IO8gQQPtsdMvXcQJXBHruXRpQDui/WXXWIkfBl8UBE5Pcxx2Cj3Ew7kQJ1ayfY7Jh4YE
/tv1xSRVud43nHyLsCWgL3K6riHtvWRLR3N9eEPDgknHcJjm9VVncuBDcr9jlf8jiYgjZ6apakuD
q7RQNnUliz8bZtILc65Vv30wrjxoY6mxEiwstK3JumsDjlzRkYw2f9QjELG1vaZWEfsdbvqhv7I0
GgfGx9y0YroWPl3O3Sg63oW4psqE80EtGET3FvbMHJbxpbghl6YNrK3t3HiPTS7SRhJnA+nU7xJg
soCqWPLa7yAMut71jrKvflyu/eX3seIActIveZ12uu+5qLT9Bj1cgZStO2ywPs92C30mAxo7fd/m
URpUWHoHLcQeyatMMpTwMDI/Td2VvxA5ThskE4FyhmMrjqt94jOtNmLdPkKrL8E9IaAW5W0NLxUk
I/BTimIA2U7K/3dZsNHLEzBNv1Gyy48xQ3BBTgx0UudUWSgG7bMPmQNpYmaEDo74kyW5Ga6AlNiI
XYldEmOV8fGtw+uXQvRjJy/nAiz+9yZnvXh13G+gCys1I8um0mKXkgHUgEMo1ev975klBxvKVZyr
999rEZSupyYKM3xDV9eATH3f+YUBf965R1g0I8zC4S03YFqnvp+KQ0B9Gg+L59QRM2/Q2tULwmxT
6DWdY1B+OfaNqqW8GaV5e29OHp+cXYk0ecDOqdvShfoxstpMb/dgYjOygJmg/9RH/e02PKQTSe8F
4CxPf/xFyAGBXMDO5+4eqI0f7TtwUY/l0CFNiVTxgYOxC49MyLPmqWAUjj0s3sgn6g7LcepqbXo+
eZULOri++lBtdiUN6b+1pJ5BepDxG9fIhbyjyfUSPnxHW9FXmqZl/uzprpyZTJSidEgo1hjCh7u2
RM9+vY3epO5R6WCXs4zHqqifSvhyFE2h6+GDEW/fTb5fEo0QkR1Koq3ESQEKaoRw7o2KWKRtrkWX
x+gelCKt4SCr8qt2VQjTmcKbMy8Su9bRcgvY5IBwmuONWc0Hfe6ybb2nTmZKk0nnuxEG1BiK/d6w
P/uUvQR/CZmgPJ4HEMKsTCtsSVvLBsQ/SNyRSEcaxHbeCtnNUxMsfIdCrag9uIe8y/Sjvw71/yz9
e24uqv/kFJWK3XaRFz+ZK21Jgq/UWTcN1G/AYdY8jPqFNc30QLHKUGFZjVGkfhXIMih4m4nZS/ok
l6S0lcTWTQT3yKku37fcJ4HPvTh8LTA74BgCTrtLorBwmN7MUy3PouAJ1vRkxaIamjfcd0gTtWgS
0EcEw0ooMZ1XvGU2al6HbJ4gxvaAp01O6sGRwquwUsytzHzQUoBPxUbJbe2CPeT7R+drK0vGfuXf
QJUZtDarK40TDm1zAOepSu2LOqX9j8rXxqktUEzBf/8OBl2NOBLY/9w4u2tWiLIRsAET6i88Q+8F
iTFdYWdBDLrguk+gyD/U+R/lYLS8JFDQdFVi1ncPC1c9s4kyrLHSeOc9lcnw0mhqkYKhX3iVOrTo
dWHlYOUp3ji1+2Cf5scHLLvL5kylbTDdYHdGGuoNK4Xz6yhVy69E/gNgKYXdnz+y7DeHXWtqDgws
o7qh/QB2z0Ixgkwb88OAd6oM5hYAlDgd4OUqYmSDNSSmlndY3Sc+5Zevzup/G2v4+I0AOWymVaRC
E7USiWrlzKMy3d3ssohr21Yh0XLbM26pXfmZfp5pioDmaDviZjBPLR61zMjjwG2rmD4KCDxgmcIH
J386hWcqSuaJ8pbXgob6Rq/LROUQi9PRQgOG2AWXV39meJdkPG7ndJYiF2jweHrl6FVTqRLRsnHp
hhxU9NT4E7APGT4nqGEg8PgO2rVDasT+iHlgtEmUJcHZjljAOsk4Clx4xGcicO8KFX8nqwhWlLxj
TSxmVf2UgP3TqbXyTNYT821OFxIHd6SXjTg/+/KeH0tUH5HpQ2zwKPbmqE/L5DgJjkev0lMpWTDV
uj236qAXgQh3pjUYn1Ow+V0Klc8gSCvZBsljpoWrHCfRKxChV3oz95RvkWBqfyxfqIebHUnV4Kgh
fd+kDr2r9hdjDVbuAzix8PM3U3xuo81Umtr25A5bxNZmSnfO6Xzk8I/V+2hL4+A90L/Laqx+cB5E
XJX0dwylE1xW4qzGPQ4OcbZ7yaAORcMCwUaxfe5MtHWCJoW6QOqHxVSh/70HmWW3jDxkZMFBKkjO
jxNZk21SwhvsJcY30j2KORxdpMOlqyKAMQsPOFWI4LsdYvHpJxb+YsJ3JkADentJBjDv4M/wCaOM
Tpt7HXqgqjfC1m/7kLPasJ2VjNjB8Wp4sUPA9DN9Dgd6WI5wyvI1/bsuRZMAa4ofMzqKh/5O4IQR
F0cesbaOW5X6u3Pw038KE79kG1nKr5KmvJQ/iFdE/1VqdptlloYcdoUNmEyk78x+YkBMfgb5E0FI
014vhc7AhFm2miz8Gmce5I+kC1GjZS1j7uYUvBheqXo52OfdDMB1KBnON7PSpffiSFHC2Og1TQzA
Jnr6TjfYGV+rJ2OIQKxJFxy5GlUc3ip2o6PhoWc9vJglCRf3C+KWduTifgsrH+4s0USf09KfpHrB
sZD1H6vtjdnJnhtFdBFl/BaTuOYTpV8GkvSAiHy+oEtPe3SeySP9UXjgd36t/latPApY6XZ0K18Z
8yEnicYw694nHmHgeEEU4Xt/czbJasK9gjfb97nkw5FG/fEN/L/e8mi49BxDxLQJwQvBdL06oy1Y
3LDCDiU5fD6LuP7H9Kauo6zujkIgFnmBKRxVosDref1kPavKfk/+4cS9c0gBvqhzzpdmwMNkJqux
aLlUWF/D0hz4+rbL8A6wistXXxJXK0uUYAxo8gbnVyD0iprqNhUMr1fQ0BeWZxbHQWIl12LRmApG
Uit71+6JWKzkQLEo+sdxp7MLVAGydhzAq68hccHpu/ZpPLPsDgCJZ95Gi1zFfpShUI2bvldjiK5t
KqGIqFnMLxFrghIV3MHwLaLbPD1CO3Vo+/Yr2tO8l6+/oRfHXPzDiyQIVGoFUR1ZX9ssyYUMGLt0
Mg0Sm2Q1vfQV6IxDLiVLfUBNSZndFHE0uKSLUPfOIBxtpGGkUDz58pxUtQ+1/h5DYInELMOxtOcp
gEEZFT/BTxYrR2IIEupE4GPZ6DDNcgED5raoymMwt1EMCXFCn+XOGDLKMd5+qVhf+ItkRNgW/wv7
5UZ5HRLNJh3K2tY8V1sVEGGDJdcNSnWUgnJloPFoUJzxci5WYo6nVR72IW/D7yMgJr2olqnZwQtw
cH67t9/AuVAo60QrT9OVfRMzMMlmR4kgZC7JQCm22atEhsSZNxrLyYfILkWNl1fTLCznSJX6lYSa
KSvCtTdjVYN9dCjcpygBvsZOnGsFxUH5DJ46THUvyktC4jabq+mZkoD5iTjzhaZ7ExTuBB9OMBRK
/aVBPQNKQrduPBq8ZRGhhh2payGTPrH88e+2n09iY4P3eyEia7+yFKrJiIiRdPd5q1/1Jq+IyJli
20TsZb1qmoOGgSG0j81/eVtoI3CVgYldfYITmbEWVDgPTEhPnI/n7XJYS0ydMXuNzLFIcSALT4Ff
87FuyNC0YVLqweIYMH+JM9FgL5pb8GijAMUbaSscYkcKlYj0OMMG7bbQKshisaHg31DEIG7ZTKbV
vjMmThr6Tqv4Wmr1fHHKbMr14QD4JLAwjSGWw3JcY9ssyUnl9wsZSaEx7pcxvy2IUIiL7aKJMtiu
Mml7CbLIP4FB21s8MCPeCxqmXM7sCjF8l1e+fd3nPiqzwymxtOWik9oFX71RfiT/XyZ43dYA1YmB
24sIlj9kbRrkYECeOviq2wCC2QogZz58gZo0b6P77dpV8AkB1BTrrdjQ+LBhgomh5htOy4Ijmv3A
velVvo0cN/tqvuw0S/QCoZe7Mg5btqYClpsWZVYNAvCqN3DZLbuumTdq3zV3EfhhThOvFYEyT9+w
hKVH/tRD2/H3UsmrconuCv9mj9c5yndbqE212rrMIS3tlnnM7uRPUhLlMDThKKhhlRqzJXqTqlsm
P1ytittu7ndYd9O4bG5wGMRIXMenW5RRdkaNzj01woIL4ytTXlvHaaDQydzOux/E8sY06UEJUIX6
z69hhcjess/j1ew2WMa7cfcy+2y5cT9mcxjWdnKPXU+9DIxkfV0HTKJqjlL35kxspLmQJeITaauT
/ow6EUoZvChSHg+N8daIFDDhC9AgY8+yPzJqCetEz5TBG0qQpCQmvnR1eH+ZKo5tMqaaTXGmdyBv
mp1WychVFg1ahm8fhMdtfNQJwvxAwFcdPLksHW3+HbKmWG5NirafjgwMKo466aPRxxlRp4FG0Cn9
+B+NK//ootgc0IzRw1kiSm+I2rDr/Kcdqq6fawEls9sw9R0xKIxLp0oO4aeDVnzqqzj3QhevYn4q
CQMygU+7TP3AmNrt2CrUJzexmliGtYlHeFMKutk35zr3FHI+EC1It4VxWExeKXe6sbPF9BY+cejm
QbdA1/6Pm8hiDH14Ptgo1o7/TYk/1kYXapEolPxxiyC3+ldgUUEATysK/O9W1msIeCNCYy36enlX
Q5+dzTxpMm2G1VN63gs0I6FzQ+MoU225gl77+1voJrD6Cz3QiaqzvXyUPjbFScCHehXM1MW483CJ
/mlzY4NIV6TfU1WlxAbSjhh3cloZ2LhYGegVFkp9s7O2tXl84yB/yjeMJwlp4bvA3HhlKCikSURk
4L5meQ6FMO61mNrYmdNZnAQtQ+ZEctIFwOLrVNisS+tGP2dnwzACWFDuQE705LpJSpT9eW0aGKv1
lQyOHuGOJrDIrApvsVgZI/aOj/UKsUaQuDW3d1AqaOJRO2i4V2jLx6GxOY0eDxIpkm/+ovTRPmHp
EeqnVbUrouqH7xwRvV+UhJV9cRcbeUNaTKbXg4Ws5L2Bmz92TcEQKt58vMl+M6u2ovXK3aH872Bu
QJmfxAfNC9tQgFMM9bUeajNjs6yK9i2ONI9b/vmoBhKGtvhgU2/ivvwqg85QIXsXHH2D9TEzoVh8
XQgOZDKekMOVOcFRuFHFu8bQAYbKf5qRP9r66rsbD/f8brA04kiLErnckjZ4TslBralZ9UnMmGGc
Au5s6YnkeWzEIyHu6xR6RjQCNsl2VQUxhGIsoV4HnQppx6nkYZfQZ1qTTP8MTPxxbF8MeDrgTk1d
VsIgHourtdsxD/R9RZo8E9jhi1aPkDtTpCuUMQW+sGVGRfSWcK+S/8lDEZ6x6zvrK2LkoUm5ul5B
1WMUISKQ+jPdGFYxi9ulfz4VCKe1FoOJdcc6H2us2lQzqn6cGCxLuF1xCDjseuZPSsPeics4PzyU
azfm/z+ZGEx1zDolg7Nl79fA+MY5zL/LRBoE9BfMnqIWTCvENmTkvhmC+fBKjwlLAL49ptUNDesh
CQjmZedKsEdbAGJnp+vd2FT3IjOW0ulgPRRdHYVuFJ/Bp/sB0eftokRC4QSwFNcdLgI838Rxvrpz
omhSSz3u0RQD2l2suD4Cch/qiahY9VUo2+sGxrIErMqpAmGy12srZJ0teI39SS2aLuLxQUHSzCAY
KZlaOa+YP++1CVNjYa0Wc/9KODiJmj54MqVbOQi8crT5m6d02f8nf6aSp/9IvUetpMwJlu+MlhnG
0+UWzZW+OwkvWOdmPu7o8neSx1MQVV4YAIwaFf9NvjN2ssyf7wHobZfktiy3tmTRLFv/dacT2t/R
m9Vx+SxlqeKMPHstX+7VuWfURNWWr6i/SMwVAw3sJACrEX/8rBeW4TfpE6WmzvguXDm4G2cDACZj
Zxt7rcCSdD+nK4ciqLxIO/1G5w+pyMPNBSnwsAYHMtFUlzRWHc0jh7u12RGObshlZWf5AKbCcQqq
6eXHOxZn8HKuptlxt0f86gmhAATpqNaaZnwmwmSuBp6anwTZvc1mUpUqPRheoxE/ksP92Yem4F5E
gnsm715cjucOFslkNKAcLjgdlTeSj1G0BVkyfLHi1vk1xMIrszV26+WlNS39O542Ba97ON731SGI
8/01CCSgzSlLCiGop/ktndF5FNPITfglbuOdY5rmHLLVbRkmw8YeiECUoJXkupBeiYs7M3Ypm73l
N+a+gDufpP6tGzxHRVCyGxDUhknspaSDl9ZTPNgpVIF5e1xbIillh2XZJv6d3gzpqJH/IeiAKqQ0
ny/zRnygzrL5+09pe8RR4O0RKom6s9NM3JxdB3pP8193Jw6pZ5IgQ2MGigNRb2teqvVMMIs1j0Bi
vC/1zz34+xEekC9LTXbQV1l6P/AkerIDuj72mlYgyxrQe4hfyGF68JxnyMM6gifFzxuocDLut//N
n7ZvVnbFBQ9yJhBDoxtAYqpeP1nQgkVyM9h7n4zBSDssoTCA6Xa3xrwdLqLTfoU0wtaZ2Vlqebgt
eJyl5tqP2E2HfH/CPQ0sSXpoDqNNhwOAbtumdDZ65VXKC9IAlo6k8onYpuQN1x/QsgBb6eRMbDV/
c93vEwdZS8GGtoyD+WltfgmBOPRaO92KDu6/3hd5UscA168kirFUDv6PKQyfN0v9fgng9N+DvvXw
160w9yaK/IYtoZC3xf694Cnbus6cMo/nGTQDlLHBOPtwKlf78fai4kruWVeYHyCtiMXOHP4RdCi2
b5WOeJRWaRAF7SZbDJaTYqkE157o16pa53hOBcv7KMH0sExG54SpCx9FRzfIM/KBsADkZ1tDKwfT
sjPoGlkiyE9uXS+BevpvTepOrTCpymKrjAzSFvP4sQj00R4YSNi3CBz3az98En//Pgtx6KHnOC4y
155l4XCdLkSXbMl/a8qJ7KTXJtjvoxGyCz0vP21uSTnPx/50AVvXotx4CVA84+AZ6r+o2ao1VdDc
eYB545E5MNi97a82Odr+8AehDdWYYpkFjBKPeTJOhs8Id/ly+KhoPL2EbVWePlJkUT+5n1yCFimu
aPL3JnuspQiCrtkdBr1TTQm0f9RUUU2RpI3K+BAOQm0Df8D3rO2CVgVci3mOY0LKEb8Yi6gEqrt6
5QQswWYFii6FiVCbcvwbkkjegKbQ54nLe++bX6hEIEEtVwyliqlkMfiAGP5r0JDc4FyCCj7pqmrX
ygKw6rUSw2AvhBIDJatFPnfdyJlRhEuumYb6tCyElImmYwZ41cEqzvTkqu0ho/2XMtSOlY1LNfXY
bjhXR8xNZ46/aswzBS4ny6vfhjJg6EYzPFMomfeiAOtdgRloWGz6Sdkb+E7AJ+MFRcuq/RGRQlSW
FIoW8seOIYo7N8Xfrc3dh2GI3JYbREEvRr2REbgnQR/7SUkiWYa2OswVq7/dlrlf72AMjrJziwiE
rh8ZDcf18E/BS/5jajxByuopNe9jCBH4dWQFqMHZ4+RT2yzvQQuDgC2L7Xs5JoqeijlyOBVywpxx
hHN7x4s2/eaELTYhjHAL3wvXWp4iYcE4+Yf1gfsdhJDfPct0iPmASigNqnlq/Q7YH5lPuuWRePHh
rhdPoEtfyQIGo+5ffaUEKb+tJ20AnZPd3KFm+rWqR3eKKDS3mCb4c4CImAzfGCP2eEk3/i3OW3Q7
PDhJxxsPVPCB9sWZTyZBT9mtVph+65U9nyRU1J/8/FxaWAo8KJjIhFG8QPTRveoVLBkKqv0weJ2E
reEgUvZbwy/8+PE45vIWOj1q3YihZiYlaPLc8v7AvhNhZmsfkI+83OGWsApgCvsxjs10Ape/Lp5u
Nb7WK2PVlz1ydF6RTlKRmlWyHJnfp/g2+Sh1QIBGE/kkGkH4tF3cD7pQv6iULBqzgPzvdjMJzciB
OGYwrGVgN8KK4pYELNel/PzqyH2t0h24rT8oSZQBaxdetyQO+e7Dhc2Ez9/LDQz2b48Ot1F7J+LB
GgMgVJqRjTrdFX1qP4mqxYw4GSJ7MA60Ob4SMEuuuJV8n2A1f/h1xqIU6pb/wqkJxj784guPzxYb
0wOZfzCaxdvfIuJU8/QCfKKuQZuMGqEpPaUlpRNzUek0UItxmilxJ2lrCwkQWHwjjUCF4/Sb4OY9
P3/PFbt7AfxXKsVuLZzEIKNtSjJUXndDwx/8KGTiharOIvUfLlV7DkcfOg1sPrznMyiwJ1beALnD
d6tHSOWA2MY6txpHzZ4dAULACKzE0ttNk8V27Hd3bl/CQoLDEEOowxGal9M8E43fhR51xu9hzIrJ
FDG3s16s84CaklGzG7hBfQPOPv12PeXNL2L+Ypy4RzqZigbJi4px5nPo3zoFu8BZUyOJW8+klTIX
a+UnSDJA0Rg/0rVCx/vCLO72PgaegbyN7+tSPMBf9cZJ19SFI12aIp2HhflMbFxheQplPgeUD5Oq
B5Rxvnda1ZOf2UlwwIpK4+D699CkX0PCF/HnQsNkb8kNYy+AS5EWw0DnSvJpBdg+gB/Q2Ccp8oNi
uyR/e8Bf1jm8Rn98ZMkcXOTLEZtGv/vFIM5nv1xD/arvr/mdSBsB+Vs9eAttI+nhMUFnQACAhKOc
TSHfvJQB3fVI+DGMe8wRLMa68WsGoVWvQYUC/Aa5mpnZ+NeKxa5BNvrFooTLIYi1YC0BGU5XHVLQ
y4h8XdgkrDrYFEF8kbo0I+7GQaAVLIpxEcrERRMpUDTneNX54Z0/tk6jKs+wMpKbvffHedA/hqer
yK4+FPI69Vzv57tv1WH7W+sINByr52PkKj76gEkJ2v+dR7vm7ixtZgtJFpe952pxGPnSgZW3Hng2
c2VSkIUy7X1JfuSO93yjhCqK3NgAYIQBnVn9mwsfgW2++cUpwzQt42yt88CMdrGQIT6wvCNhDLsi
lp/8EkP45gxYTl3Gn+0hxgKRnUL+6dYvfpk5F0wp5KQTyF6dWkqJKsBaHMOHz3uzlxbEnGI4vcJU
Db6K7I9gqO/iS9a+/wyekf+OoSJSV3Cchwv2cFk0DKlJ+uu++i1mzAfm39MFPpmNG47WAoNjb5Kj
62ISz4TVZfwRwOjvFmwxRoVUTEmcD8x6YbjtBRiH6x7R3kbw3u+cdSHcvcv0UqGTw28Eu8MHGeWc
EQV02I+Y1/sjDHxfZhhfyUgRaqV59BzL1Koeqc7BERcdI0ZPX9KbiRV7IFTQRp5ZP4aiFMk8tu3C
s7i55K9NL53BX5Vib8ESOM7ZMc/59nnRL2QbHcHAUPHsOm2J5D3nPihFEqhM9HoKbpBq6MjCypTf
PNAmWEGh2RhJ7GM82kVWIPsubEjrAspVbswOSaeAEbKTZpJrib75NHoY+s+bETCy8XPj1/EKPy/D
i78zleXjAxPEnblBE3DeH3jQN81zuR2nKOjrQSdYYTVUP6ndhDbJroHff+hCBTU9+pb+4g0wkWO2
N8l7PCt6KUKKjSnM2Vn1OEqxfeRCljDNHqqQyHuyE9s+02skqiAX3yl77G5OqxvYcFQTzC59Z1Hj
QSM6yz3pH88sdyXgADOBjNQaoBtt0kNSiFrlmRFqfKHx1qV+DPHRnkTjS9i1N1frgokmI+LS8VR0
QKO3e/bFln5U/Dbm/XA6C2ey2TuUxaeIDK72qMh36aLT+OthFdqn26UcY2VyX6mxY2xC3Wtf2Sg9
0forB3fYbgPbFzKK+dRg1ggvJaM/f8HxyCkdmKH/jyHvcs+i5YCARjWMi5rw5lRv6miFuHEHe+tg
l5aROfMM5Q4xANvvK7Z5qZ8hZyWcqWjeYSNVVZNa+B/iTTYmToAHvLZvcsEEegpp5iDUiQHKmekE
EK62Di/4qYBJjv643DD+y1mjM905pff/HHU5wNK+N0WKft32SOFO1SKbzRf9RsxpJYGNOmO04o2r
65ndQINuPjQqgeTWqKbZuGFVc6eabYp/wSLAm9rDsPG80qcGhPnG8mzVUCWoKYQrssQovMOiwCzk
AHOzzOmJGnZSHfrALtZEIbkEy7fPild6nUU8jkI1I1seGC/jTWouf3jyANEdbKLQqcDnfA/3MT3N
QDLK59T4y5dznDPSQmA3EU0MWu2Hgd0kk0aJJTrIcEjZ6MYecy4dV7TSs5ICYwql/91vHkhGfV3M
PAZJUXPWNQ5hrt7IgP5I1054Nf70660nRY1efXO9/pqMuhL39Ho+29ltVGxzxZPYbot6GOSj5a/d
GyojsOC+Ak1Ib9cgO4R22QVaWyC+IQWFbDxMX+nDnCNd5ceQ+e2l/ZnY6gmVFRzNfUmatbg5LR4t
rw1lY6iC8MCYlf8ccbgkBlxk6LTG3FECh6GSGxo7TUe/NAgIP62TjYzHl3T/g8upAVr28JnEvnhF
ESDD9Pb/yafSTrmSSABJQkRFnLdCdIWny08ctYkqiirgxhTLut5reRCh5R03n871Fhs6g2AKbOwV
q/V5rfYWcun7ORIDF8q+mkaBpJHzVK+57EiT8WNZ6Pe5ffb0J1ktduU3IICRsEFvcryceOd0x57W
huHJbaagBIHiqY30wuc9j+je8L7QHzAYAz+aNpm0SXfzzCnqia5OaBz95c43NwhqFHThXytgLAFv
nD1rpHGHHbmAZFt2+IQLPTH82dwf4vAQ5oro8zrBNT/UwxeALR6J/d/PlbE8s6xV2dJB1zQnvhL4
8gpU32ymMGKy1T6IhFAVf2Nihhpyw76yCZv+bLOY7heB/6Vj73qbhB6GLhbFi5kiEt/gH0cINT3U
64zOTJ63GbAJHPZLD9e8g98fKQmri5VKWUtb9pFOwhxnAPNdTSoEmpb9LjenBrpn87TFiQlziYxE
2vOr9HicS2eYZ30Wol0GZq3H15PA2ru8eNnxdQigDv6udoZnWdjcymkCPykpYe7b01wY56ETWZ8D
IdMFe2mlasiM9afB/p41DfzRNdKtkmkWr53Mq0sab235iZ+sdoEahR3fa1HkpCDVcMSAePIdB1jj
8k6u8bQpDsLH+1KlgTC1Y4YjeLhJvCGO67Zz7WhgK+o1nLCtrCDZMVnPnQ/l39fBbz586ODkyUfF
GPaT+xo+7OwsUW0ri6kNucr3K8RO07LzGQu0Uo9E0McF0PZjhHRmYZpgi50VBk5+I1bl3T6TL8zD
GCz5cIAzOGwTowfCEGPlt09tqg6tBOcNED2s0Wkyn4xJz0AE4mDWrkfw/331dZw3+2iw3FHWUA9U
odR4lUOug1GqGn0WPUrS9ZH0q7tpTe/TFj9tjkZZ5PImjHFEdstvQHEkDj5JQ71omkmE6Yq3jVY1
HSu4ZnnvsCQ8w3cV5nw8epRW1iqS8QZP3HJqHLXGkJLr7nzbBExns/3NDbq1CD4wbCONUPm/3Gp1
R5+yfbR8zKfuIVkPNhD0gVS8NWJiSoKm4LdGfENAE7wcu+enE2KrFucVy+AiHbibsb6t/bhJIyER
83ACUAxQb6nRbI79SBZeSQCwU4f40QgIsCZQCd/dHStt2ZuAdef53GUQEw5GExCwsi1172F8jgJ1
HKbqvBFX1uy66/XLb9hEXtkHdPHNex3l2+wmcUNWGt1yvtY/csVF6IfWMEwjNJdYmAJBK2A3hw07
KcMwolvZPFCN78x+zy4If0UR/52U9lKXNQhO7ZNr6cU6tdCbuV3Lwa0qTLnPT7aqLn/fdjHYz/jh
ew1T7xZajjSzHdD6e0yKn5ensh3Gf+BmYfKsGiMsKqMJiK5k6aUTASZDXc3VXjkCmdZsPwtvT2sw
LwjnCG2MaA8t8qG5MF8gPXR0NlwEJeqsA2pOIT+HEZXXU3/Sd7YFaDVCPTNFMzG0gP1+R4qSHNNx
l7QqofTikKrk/Hh1omAwR6OQGiwwIX9nZr9uWVhhe231DeHILMgADvPEQQSzWzzgzfa2uJx1tuxy
l5A5mNOgCPBY7ur+ZBcsUQRTOk4VLQ0NpbpnnvNGvuPN8U16Ebj7ubY6ZOKU8GhL6/jbQ5CghnYh
qMzmhjUhfoLlTq3XZxS3FWpsRitdmEDkEc/Di9M9zi+Wqsot8YMYcv1RfVXmP3gAutWUP7LLEmyo
X3OEDRWJhDqQj70xQgWXuWdUMoRkPe3J35aguIC5iX3JbJTzJrk4NG1PZzs5BW5YcEBawzxdjx0G
rkDi1TVVRb1D9l7oPgk8Y9YpK3bu+/i4mzUlksLgOZMh7S8nE/MIT38CMp0PuiNQVzOdTNVqjwE7
11F9Wad/wKuf/FAIdkmQTzm/qFgvjj78n4kywVTNXEFt2wzGx4JN4/UwsYYDbCCp2wphVsygj7G+
Oz6TeOo5UuaQN5ZtySGkA0gJbhaOSw4zixNsMsbkNgTu4pc5AIYoaFleNH0r6TvaqBh/lYIkissX
tnHDjKLNd+NP8d4BGNMOfpcc425LDWvr23EXsdQmeprNvppa46N47ntCglJftOrGvmfVg+5/9hux
OYWoqDXhCB6Mk3nn8WTL4Ydo2f3c/XN7xtN2jhIlUbqZJRows0NajWM0J6+K0EiBvK/BL7D00rsS
ocwLFyp+8rgMzjw+o5+JZjX/tEa1WIOksNUAPhlkqZ63ULCcl7mbZtQA2UC7x/PzUqxIu7ZhXw7T
hTU5cCAjUs4SKL+Vbi0WT49aEbMQrNLR1uCLdJqxgVu0ygAyCtoRB6Ski1NhH9n/QInL7GmbxS8m
zjNcvlH4EZehivL2OlshAv2FTIzOO572NXgIED69cv9vs4t8FPAhyDagSICUraanF1upS2Ggwgne
JE6GAZNmMdBnwGhxojSGEpaIemNZAGyaZy2Adg4m7OheTonIszxNXDL+xJsHm5D/cQDLzvaP1RYr
6P/o7b1ytWpEPrrjVj46UKK6GWKYn5uAzSjpE8de7qqj4HS3wTPlJluYctaNAd0PZGiq7xjcK7AD
q9jLnRKN2I7Np25isGV4rVegzyHJIQbhMTfwRC7h2UGMlq7xszK0agZP2yaUcSR1H2ZQIb8Y+VTA
bg84DTRiORIv+RU5xcfTvkelUQ9F+HvkHRD/OpOL+nAAbWDC7HeDGTrf/ofRUpgWEw10MJ5sw82t
7yb2p1hC4vI2QUOfyr1qB1NJq0lGcKD4TMKgyhF0xsGK3Rwr4KrtxH9yXZxk66OSU1z1JVNRAu5a
h5n3KTtSSl5CReorxq5FevwYND5Cs6JBfSsQ8vlpmwTtl2fc9qK9+OVj6GM7nFP0pMQRv7rv+6YY
JmxIRifLLxCbAfqpaZOn3FJQMy91h0kcQSLyppsqqBHduqJu5amDZAWUtQjriKdKYpx2l7tgwCfg
2Pizva6zvX56JKaZU/rjenfS30SJESEwYAlGZdPLlO4vSHvuTdsE2TZY2jCXxK5AWhcoNjzL/08V
VN7vRsSvYju0oFEYsfeRkt6i7SkO3tXlkkeSb0ObceibTQ3B0gIIOrrDjO1y14JeqaATFD6XX9QK
WWZoVMkk2oWlDC1qcxY5P5uztzNrrq+SRPgRJqfGWAvvh7uInQCvXTi7J48Nv+BQnFsC0t6bdxCM
uruPQKQyaBoituHPo+zZAVk5a+sEuiqxMvl4IGG6geZCQcRPuq/MhcoIVFjkgU7jdedamIkqcs/e
bIxJmDa9+LqVLp5nvZmmrAFN6qtmWbB3I8XRIwD6lhq0zcNf0QZs3RxLltCXL1JNXFpidgsaciI/
tPrjAO95th21UVIYXjS5NOelXN8LaJLGRSuxurd9msuUq3Zc+y73SIwyYivzc1JmIIqPZVchjiiy
ypEJZvN4MgvYd7x7F+yN/WaGyWJlpkaT9IM2pbA/JPVwYW2/czTbYyUuhwii0KaZvzyvRaKRMZ6U
PMnWXOAlpuf4DOvw3AQ+mQoztaDbWqNJLxSEf4j7+mEyBqFCXWk2CGke7t7Ch6Bbf7SjwajEkjpj
xLlhxbA9UPX7Y6aDqQMcvCWpQ3+Dxx2ZvNknh9lbCHTH4D+gI0xHjmn0U4mezoHlzf223YuqrikR
J9sysc7aUrTNF9z8L/n+zNHRL1Xn5eu3prK85aV7SB5JSQdvlpNxrs6vUd7aoZIHQzlu6kDth39h
+fVgLUmWvbJ2hNAClxW/IMwaTmbu3nreybgGI09qt9D6sa5Ci2eUgf3VJYngv5G+9OIPeP43g4v5
XFRRchKbcf6zcTFy+oCwJGghtTTRb33mcNXUS+QzCj4m6ta2AYYU3CMEcAQZ3YC20wJETF2ssDjF
WGu0m3EG5c3vp0Te6VYHAyfwCWFC9VfZoQr12dhWBRjZGs37JBmbTQnrPoiy43NSWgqYGFc/nxOi
73TmHUI8exS6Vbt/UnB0dPpM/kTn+Bjv68KGjZUjauacPpiZxVm3EPQgQ/zEkDcyP7gKnJy+P43r
IWD+zoGSOog9alqpJWQRTpy8R1immHqMNFTMQriXGABCxq2GH5Ba6f6VHwuNNvpkKvphoDDlHBFy
lQCcyzXU7rvNo4IifLMCkoVzwo606wE2K4pjLbVKDOsoYTHoBD/0YB1MEK6M5c1wUNNqdh3dT72l
YKSbjeV7ninS4VZXjeaTzoRKcSyMuMVRSLKsOIIMS1w1CCnWp8YJtbib4jG9irpS0+qtgoy+EZfY
iupT6TXo5XZ6RSVp5HpfO9LJh24GPXThzSNdZg3ZKgfyjqOyuW4+a2fd50RUzOnRDKJkXOp8qR0m
3Rtoet+dnDBoXawoMfM5tkj0gj6x2HzRfkU+YbtBXvRFLmB9vD0+SuAnXQyoTPxFJ6PfpGKDkW0x
F5NegvsM34bCRHudvZdfRYEhYu2unv5TrNP+Emx34JTRRLbI7ECu1ddGfN+/oG0/fpIH/EVqEe3E
kNF3J57IJaJ8Wu3dkCHlIkNDugj2OD6QOiwmfreMpCmmDej4ShMFHe8++E6NP/ISN2GdomQHh+K+
+z8FG9CKTXWPiHP2klN+hKflK93/RgqOHSYAVH2iuX8vfi67yZszrGbugEFqZAqLAr7iw0v0Mo4d
gBBRZRkP5JnkKEI35n7dKZ+tkoe71BjMgpCYblVnj2wCSz+ZsoN9YKJNNDTXHi8kedn2tqsWoe/5
kfwhJUI6hRivlcpl7MSU1r0u32bqXg47J4fqrQwNxbZxn0CtZD0DQg/AaSIJw/uyWPnjdghZ0T3e
p5c9Oc54qaOxA8TCZtKJ4Mu2vXTXI6owviBgWsrmLRx1FQ1hvfAxuA08Rl21OLXhyWnQKIFcxpAe
b7wQY+dYBPw9OV/qy34URr0oVvFHTz+TBl/J2F6p/NQkI7TOVEL8ONmIfQOAVe5z+u+RnB/Dem9M
po3WkAOxu1A7uyiH6QdtyfTUsWkHRp07XjA0CjO/Dnk9KCawRcz7YRosdhLVYeARCbgmkyPPYisB
6Xfsd4sdXKSp47QRyBY3IaqI/WrP+71heoMm/gF//W6r53kw/Q4enBlo1DjKj8u3GeKH4e0tF+SV
Ez1IliwrFu1qk6MY2rs9alcn7qn9ePfYPIcDxHBl4ISwGm1BH80uH0SdnGbuiRPz/nKPjKAhpE9P
2eVN6UV0TqRSzk9lSKARSErdzTP5aMnd6KYryfPpP3tYYVM0ex0LLNRkHv2SOLLENFcuK69cCd8j
oh3178lQEqUID9N740BBEARDvkoZZGnXcbOr14Sc/sgbmOgKUaOnmA65HsF85ncA6VuD6PnL6B0s
wEwId8wYiN9y6cQrbZ0es9Sz/L5AC8oyNvGzgE+59T8V0J8Be+5ISYwee525w2hcqOuLqJKP5ONf
9WUHMbVmKxtmkzIbzK+XDiaAlqarXiVhk67DhRR86bMPqaphiyj6qn6bgETCpdlb8srFXIcIGToU
6Z3Sz2+aff1rCk15z37Zr7PraecAyHhiksUhSQD2zd2ktIa9ZBzh6wA1uanO+1LaFUuqSoPLBcCn
zQN1574kSi07M0cj7T8p6cnt8KW3EXkQS082Ii5VNVLjeBmXJN3pQJRxTS/3C6EpNtBFNz3nUEVW
I5Z0VdQ4+Hcq5Uk9CKleLxXJtWU5BoWJghDEUlUJp/lGXQ7pxfqSgbdpACau/x8qXvrnn/uJu63f
LnvQxO8M3Six8fnTBnwOpkhutepM5+ZY6yqJYMtAS+gP4z8kqtbvSZnjT9ZW5sAdpJBkS83TX2o0
IvaI/pjZihSSeFp0dGPMm+WA/NgKXYTIaevNSQ2Oe0LlAiOj6ip6HNtJx5IfvneHljJ8fxmdZ5On
u/Tw12cy/7W88vgL7MMIRCAXfdE7Q+gxgIQfHrCHIi+fp3lYvsyId49ipOSpwxF4Wt4vZzm4Sdr+
C/pd/96axif9+5piX4ji0MeJjjNJO9h/AbiPLtXfRCrlPIc81JSQCdnLgPWU7y2TXgwQ/VCBXeki
Ypx1VUwPPZ9FT0/OCxFkwfSjSYYwJ5SLTP/C81f2/9Ju0X4f4McsWYbCBImSqaMv0sQqmIp+pVN0
a+eU7F5NcQUR0euvOx+hziyBO0xt/27nkeogImrn/VQhqRq3wf537GrQJK3EU2xJYAlA4bkD5h2I
FNtW3DsJh7W2kS2+rky4/JFMT6mWeNPkarBINR6Z1p11EgIfhW76jPRsYtWWdppX5x+ebS1p8/Kp
L1grYenuvZ/CHV7GKilnWTpU6HDUlyinFH8tuxwCndGI4BSp9wvhIY1C4vwv/HMBd8kBgoeQY64d
G1mAnZtIF02wK3y7IxzmUBRNgQEW0lUDxRB2Z7qaauzP0SHt2fFCRyf4b7T/LX2qtxWNeRnATN3k
qGrxXepMMhBvGqz7Z2mLQpp4PJeCTTAKmaCPn4twoiBtKJ5ihwB7+bpld68DRTX0/AJA79WhGZdp
9jY/+Ki+6ItsAt3mZ/sls0qZwIp4oQ53wZHetxB7POQK2psbT18HRK9eLBIX+kIyuN4fP9mGuSCP
WtvHlo7I6qEEQa1Dn+OjFl1ehp1bvFEa+msUOAcXOfBX2gDL5IgXOeyrm5aOsAJW/gNafx1ndtD4
yxCg8yAKzVPhpe3j9JzV8XyPcZnHFnVVDIyZE4BaxC8pZBhX52JqsMl3b2SVfcNjonvWjn6J3DFJ
01vr4OSRc/dI0Dac5plSByf25BzRy414UNIJYWhtvBHJpnLDRdm9y3BD/sEjhjoCi9YyQ78yiTrj
olRTcR6z5X8ewORudy66mfH3FeWtRYXs3RSoY3fHj2tBqDwxKSaqSHd3du115JSo8aT0D/oCZlAQ
ccmVoPUQn15cZREvnIwr3L0QJZx54VybJMKITDMjRoKZiX3jeL5pJUi2gKucsx5/wSGyhqUcC4YM
VsZKs8ERYQVpvzFlR6ytX2SoZX+5E3dyoGB8Zb+Uo+SaTQDCPyeTPhG1adOTfngkTPsAfoEn66IR
Q0FZmP/I4geU0HCsBGCJ0w2HGvDxxdV+ZcxsZTGalv2l82liYHmpfaY7A+kcmifT/6JDVUOXT1me
uXI6luhFZFiMy7/bVwfmvuhW4RvYQ32b9ZkjKCstzRUBCTrlMpboZMJbEKRpnhxnAMJbDoyg3VHX
s9oPtPjamMyV2uVGWoOt/cYvLinxWiiybcZ6SnuZFQR0L77Re1FiGw2bmWiNJGaV0O4JTLDSitmt
2Ut1IRrQXED//zsAJ6U0z8WHp3MJZzf680I+5g2LjPM64kWu7H2nnn1DyZNah3yzkZjVWZHUpAo1
j4HY3rCxMLLCHvoDiSmgWYnxwnZZNH1///EC5ItH7w/uH67RV/sUTWJkwRKSe9f+yxfsHyxOQIv2
k+cAy5+Dl2WC4mRZamsbGvRKBb9MwXalArJimcTwXPWhZmsoi1h70OT+iWAuy9EqYuoG8dcuDoWB
a9Lhrf7kctmscmc05Qe4QYzMYDvnD8mDXlHxJnSczoyU5KlSib7QDENPgexYu7zIr5YuijImkOJV
+kcVmO7cEFbiPeuOQcVsXaROmMYSzv6e7fVDzMo81pAOVaz1zqeIQHWhrkRcQKH43KH3uK9E/mhe
KcKP6Qk6Bv4ibbqdRz07vMpo3gPRQFCDAIK6A7Eugu3UXEHeaQb7Us8Ay4L0ZlNT+dLOKSU3d3C7
RnfIh408OraLxB1FlQXo3BDmtQoJlglmUq2xKYCaP5zD95zfzlcTEULhVMYLk+JxpQ5IH6Dk4c1H
4mbl7QlyLID/YZ8I3EkA5k1jM/lBqyF4i26UjYJROuTjB/Du+2WMOttBqkU0lWqZgm91stRQeg6A
PMKlXT1wOI9alZVd/7OH0SLnIqgNU+RVQ7ZQiYJNd1plTCey3nI/EU/n9suDjmChD78ZFjdbq3Mg
h5MVEDbeVtoVHDjHCqR3AR/PI4acp0MQKlHHxzc35sO/1e1jbrzbxJWJ52U3gDeI/0Y7FUHX/Amc
27ebFhgYonzKmgpcAUUeZ0+t5xIvupiSkhrb5/kezNCYQFNhccDIFGU2BTMJjzeNhUDsmtaKepKX
RS5cWkr2f1KHDikNpBAdA/YaagmmWbl3GQ7gP+zAndxbgskprZXwYSRfvw+YL7h3vrxVSBSGVmdm
vje2KCF8wrYQ7UbQzSIbQ4mXzYgC+rU0Vz3FvJ1ACkJJ6JozKYhKnAQkNgycYKCxfKQTShRkNcck
sWy5CZ/KBKo/VoOVLpfq9naKxpVkvdZQry0yU6X80zApc1u2aPZUYLVJuJIM2GoQ9iB+Jv9+95Xp
utyUE8hVqfdC5wd9o2ePJVsyOrj+dsc9t0mIjvvwhVHatgvO/myU78YTMy0SEHyvMb5cHAIpEAbo
K/OYCaC7aw1Z73VhaIF5HTAmjF+ndRR65iefHJDoKfTS1HHJuqUdmm48Ewdz4LSVg9Zi8RJtlrZT
MDGmcqOYKS1Rm93WA4osO6MC5YxlWGAZsA+Q1kNXv8lbZhxEZetox61nNVTyUBw0CtMbe2HC2c/p
SGGlpnSc2ZVxvqwapgWuhZ5bgq/u2YrqP7WwIbXIQG0+Je29PXdwrs7PIKi7GRe6gy/auJTRE/Tm
gKtP2UmB87CmPLMTJEoCbnM30S5fJKS4gUHglViR6k/jl+svHuFVLhTwEodIyfMP8dkdlkaDlaqJ
RDwNoOH8unnsVfz//33UCwmcNw3K9VDXGN4LAodbvfF51KKoG/1bI4YcDChpePyOeZQ/FuiS0UTS
9XwQ3LrRx451RbUPFVXo9T05GeFoe2eI9GeRpmohaIEBss19UohaRAaqTfzmQ8ZKAQVzcZfVRtje
OZsynGRWXVqsqBfQzV6y1ueGOTre1zY8xjExwgsMBiMFJ//QmP5rJJHWGVhUL98HzjpR8djA2XXw
TThGK3VhSufWnz9LqHNyf6ifj+fh5ZKjjJK5TSu7bEOr7zy5ag0zUJXxNAVUpLO51+KaqXMpH+xD
Yh6UoNh0kcQp0WRH4Ozh8RvJeOxoizE6ijUg7rgIpExE5C1Y3ps0zK02+3uGXR+0PQGx5eVXo9xN
32ioLKoa2NvZNAVM1/w9hDc/CyKdKgtmBwu/Uh3qEgHf90xYyN6XH84g4xPV/3npRS4dERKj9ryG
zs06HormxFAirYTTvay99V7rk6PdE+m9LcqgURrC84rkmaq5oGIS01kc1BXh8QwCw7HbJRi6AAIx
XTR1C5+EGBiGzE4P+FQf4//R3U/C2e+tHN5F8aQner7+PQaqH7NF63siADLZtJTRWDLGuCrN0RIf
glnbvWnUzXC+VFWVWo9p9If+Pf1gK1VoDCid8+5CZvyUaPFH8H6K6r5B5AA4wdwHvTBfUK2YffuM
Ths3Ae4D+TAXHYWvyKdQHbyPZEbUT6ztTFjSA1Nx/4p/FAlT9+t60qjlmHiZG62XwmZ8LJZO8WrS
7O+EmzygaHS9sBOjCBOsIAkf81A1VzG00o3PXr0g6qvRQAq+pNNpYGCyEv05rBys4Tl/EQYZicQK
XrnhWrys69zDjmh4SYtEdHiSTUMo3/EqBzlOwHEtyOh+D5aDzsa10Bec4tMSO/N2mrSHF3bmocBa
T4oAwncMGkw65k9fapuFn7xM7lJ1Hnp7KRcesIIZyyeGC4Jy3adAn7Yoa4RipXlETUVrSdH/V+c8
0tLDIhhapI4yJHfHtfEoDTir3YXHNNOuojxEB6/kJ1HNBNVWQk1zBoh+rHal54DQ5Ti3eAK4sSg3
pMBTxIoCB7d4HDEA51AEtvPiCJbByC9yYA39+Re4Ob0MCB9fLW2NJ4gcc6vqfnZKOwns2bBlZaPu
hytFqSf4iJSR7O8/K5axMSIr3/if/dztSPqkeEb+KDNFgtE1iqLQoI2AORqvduvtxzdTvTJxHL2k
3qoVRE6Xy+VXyepc3MEfRThvV/RCl1cHZgmkYxAVcQfhxpOEUGHzoU/ODzb1UnvDJUgAD5KlMEUS
oSYRDuRNjwIxVrZPB2x+k6AxlsuRykXqJDJ2/HGji8sVvXwmmnSokcnTRItfFWqPSZqlJUhqDm9c
9LayfMqfjmF3Z8YOMutD6omsqxsQ/JpDbXUFstiCAsjsTGr9W0PVpm1iY6rBdl0g08UtQE0p2w0a
erUPoshKLbJoX1L+hAmj9ConKHwzQmaDgwg0SOnX4UMm2kA5ghW4JXKqYsZKEr9JJx1I8HdBRJVv
8295/O7pwkSsnm27koaXkNGPiJyiXjkTxubQEzsYVHL3dl5qod4eZUkQDq+BHCuPXsaNj1JLq2lT
WpXHTMkZZqp+NwZqGlK3/8caut4nJMtTahcEL9GStZcXhilIA+EqLx+T7hCIYbJHgIqyKYYnuGux
5hi+IDkfbCmNSyUmMJVDr+MWwEKq8uR1u5R4V/9l9TV1HUe7Fy78NZ+Jf6egU/40h0tWBFeru/ue
yMFr7uCRgUTdPXbyw1B0wwim80agpEN/OwkeL23KnhV/UY315GbL6tmBfEiN9/cUf7PRgq8O77ai
OGvAk1CtPyuaOuE9wScJXvkZ0kE8lp6qCaHtkPJp1CQWQnN/vmORdRVx5SLzwzK0Dn49snNXJdd7
MNTgAs21c6oMlDACOnoyB+amr7kEbAvzE2Q+VYzi975Gv9g3U8gNFAsdxjhwBxq9tlDdWSmM8UmQ
i/5DYxcak0P7R6aixpGVn9lpwj9vmMPURDuiyuUG2p8F2la8eO9Xb1Cj/DGH5q7iq3HZTUKVu4/d
eN/flgbv15tF9v0m3kJQGWU4FXRDf2e8T2Zw79RrGP0v+nWY39oxUNrEDFENbfKNf8kECshgQSHX
XcP40ab1oFWMmRmh+oHPDT665dVMcSaMkzAt/LBGyrxd6Kfb30cnPY2sZw9lLH+2iYjmY41gyWI5
1rm5boyp1uMwSNa2BJsVWq2mHDPe2d2itjFCbm7jNpT+wtpUlO4EEe0iXKFcq2TTm6ia0EhLzbE7
NHKJU/Va89cxZe/ASprnU/rOIRoNA4+SiQFuZUU2GwZfsTlXQvw8w0abC124+EdrRtob7+HXzdiM
xVJ1AhNqfWlhZwiPseKl7wAMxSNvysYHPu4eZD3eobFz7bnoWRIlLyTijMHKdi4y0YJ/iQHDMrTi
6tBPYNGDLmtk0VgLlJhNr0rewlAIEfeoF8fsc6gTiV6+pUCv7GjQkDSDQNQjE62lfCou91lqk02N
17MN8RTMoO8W2/VHcYZF1/aT8r+1B7Dz50eEVyr8ctaQRkLgYaLq4zeGSH9wJVOQgWep3YH5LNIM
EHRp2Am4CUlSajKLDJUHQiLc24v/q3YFTfgGsIKVnadzQbSPkv52fBImMLrRErn6taV7GzbzlkVk
rFuZA3ODgiJQZ8gD24h+ULeDvHIqSpRabz+Q/OZv1SobdWEmnrOLHDYTC8/2HA/OYZaLA2uNxp80
/qhEegAnz0tvQNuulPvUpuEWmPQ3j8f0La186u1TfrkHpYXNtP5iF0hRDZ890PJ8q7Z936tOHyop
u0EPYtAqvfvRPcXjd0/2JRhs23F61FKEpFWnIQDHsYFbOEYA+JSxdIfkorPxMCV9VP9p4PxsF5QA
MKuLfGmxfkEQ8C1N+o8i2ICj/eyuDp6JAs+PJ6Lm4gVGEglDdOvvEWhOWegSqTiBzxOH5KFYOXSm
Ja+f7uU1GrylGB3wVIeGDtZsPEzovVIoHpDI8+uySSFZck/HAOdv0xIfy9mAHMdUG/WwsONJG7Hj
Ns/FGmUNVL9ngCBph5oRQfrFREV7k2OIeWkH9xxaDRmVzCuCiHQu10VN/Tmb0KLTKwxnZs2HjlIs
kWjEaHi85OEDYQ/Vtx37+B5rGJddMaCrFhZOLwuAe66UVbBt4miW+iZRLXqhgVmQe66I/RlunpnK
Ew6dAT4kx6uvTDQnOT6+URgxkEod9vgicrsUIvk9ZihZl3LFq6GVePGFvTYgOY2J8psqAAN182vg
YcgIEPR2WuXZbpk7hgeye0uPPs2IKxzUFA0fRhOQn66t3ffCuM1gs1mgCmIgzKhXPuXxq/ecy6fZ
ZbGRup9+xf1cvezL44nSWi6yyShz/JDDZd0A8FBO+CquMYg57pz45G5zEDf3IFtjqzuOBN9qvhxZ
cgk8axw4ZWSq8FByapM4BgjdALJOGQNclLqi8h8I2Rs8gYmMO3eSFLyAD12lvgXutFlPJOE3IlJg
sF18kaRBsP6iHCm69NNtPOI6YIJtVYClSQ25ip4IhtoVZRj+AhGR5k0rE257czAWZ21sgInh6BTk
ElhwMx/T1yvV9XRjcY17NLDtYuKftRxHGmrZ+OKfj+0gXZIAfpLH4/zpw8YsworD4UxQS+N4DGXS
oHyZG9C8HqqzuXiY05yNCUDNAVgyhaCyGUxh6FYlD8pS07gQoFPAM1+25gPvEs8mOckomVsd7i1Z
wOUMA06jlMhcQT8mdwa6DH55yYHsq7CFPpj+CDf3KyEkm3D8TdMiJ1RXhgA7bA5r6higAAy9L9ze
ZRl/kmILiB1EZXp9zf3tgI2506dnWiNwrOYdzuT79alLY9v3MrjIqyarAJlOSOpVHtFQ+bTDPmAu
e0kISrXizZuaciwJj045EbwndmHq0YHA4rYRXjaTCuxubKT6FyOZgyuo+GXzT7muwW2Txu41MjtM
DIMgLVhyt5SQs2cRrbK/uKGrbtr5aGR2uTIRcGbG4pMRAQALsykt0ABmBANuPWBVgicq1JAYtCSb
kGTlsKAAZFcBky2kUWxuKLv/xCtdU7S6ZqbR06keonPH4H6GSNIErEkR34c0ndxDkN8T3DgMTEWO
vRdArLa/4O545Qn6ZGLXD+mi/mj5coXr5pfslG+f2FiACL9XrkubXCCuAKhEvirwcmZaljuNl4JL
yf9317zMPXaPKeZ1PvkAP8NMRxgdKFJpRBq0e454pACXtKxOJEIc4ga3zmIIukkdxOUmcRUYVsPw
G1UBSvoOXqBXOmqGS7TcIaWHJ1bvek+BOVCGs8Ln5FgQOiy2N8Sf/FxNup2g6tMCtgHRDVgpdJ1L
cFy6be+9yfCwW3pl3KfBSD62/cDXOYqBrLVz9HXqJ+p1FmzbI5tIqJZZO87qcfVoOxACcAY0+3/a
J4NwfZUGgZVhPGmd9BvDgDohgbJD1vyd3VlSdBp8nfe7cjkc5IomOnJF45oWseIiqed1DijTsbbo
79Xem7f9EODeb9uUJJ7w5HjELQ3yJMV8AsUWjTMLBvsZeCjdNHvFPQcDR5dU4LIFG+Uw7z8StPRu
xdQvNxSfMEh6nwaMXZVSyS6uLBtMBmGm+TnjqEoByXVi4AKc2WdVFV7mW92u3RDW5KonDkL8g7is
Nl00zk+fLgNXbq9DhpvnvkRdCd49uH2j9xgB1MKmfxmB9gbJabjbGe/mhg8wLUDlO82ji+0Hu1Bc
uUYoOC+EJBtvPnTeQLlUiDwBF/DzYnGOgV0cPAl+UnLLRqqkbmdcdUIsFjPjuxJQMEiV9gwHlKDU
Nli1nCMDi+riG0IXDIDZfofyHWyN8Q04vE4mRu0Ryq7oSb6z4SzjvgnXn/+dC/5PGK+Z5sdxK23Y
5nOv4II17pKcSDAmaS1EVowoDncGQ3IlY3hkajb7OmaqHQd6C7Dt4ITiREySlAV4XKRYFxXGIrny
g5AsnyVzw58xilmoHq2SYDlXmyFdPMfJFQdh97XcIQ9bv37c+fgdtebphFpx6MTX8VupkOYKdkru
jNOkOYI4udCJMsDoDh1utlq0lz8oiJk1chvxvpA/KGtrifcv8fIH+IVvWu6kP/RpcCDPyI9eEVay
GxiwJBWaatvzwc5FBP/at7l4sKqSSAwU9lOwGSgzy02vy9ObwArOVNXDR5XS0R1bVc4aKoJcVXdL
xXyiQg38Zr98dkTDj0U18xi+eRK9x9Q0cCLh0T3QTgj6YFKwCsDboRCXc3VKbh+yldFR7HPmZq0+
28+pn+B45oePPazwibqMGot5rFVjGlEhrdb4MXTnRxbtP/8LzdC6ok6/OaHdRnCwEbBD0rFba4mB
CwR36JaK8S+uJZDTrJBmxo3Ns+3tiEc+72fh7dGcm0/kB8fEeIR+gcl/yK/zwOoQOQP+cvMvvhJm
8F/3/fIxCxJNpzd8Z1QRJ8TnTGIQM5003iYxiR5KNu+G++b4RWJvvmROQ3vSolZkL3Et4Z8nVqrz
7Kx81AC3A00g8CA8JjhXdDBdeSB+7PQY6cSHqj7M56MIkuqD/KogQnON+mheeQls02+1CAn7XMBG
tRjS4TXgzX9SMhnctcrWH4IRp3+UuHQbF7pblO+GoGzGioYhNHjLx24sLS8GrusuDOJxPekxcRYm
sST7mHnTNZl9/YmF9U8x73SbSwrReBVEmzLp48h/MImIXLlEsDg0mmAh7H548ysukJSxchYaS9IS
GHSY8xidfF4BDlMc0TS752g40hvSgLJmAr60IxbWAGltrVisJjzPsxeOFR46xj5Lj9NnVr/gCOEY
gYa0veNpeGAPUur68lBHCIe3G6kjT70uf3Ziq7o5kF716/KqFjrni0PQOFzs6E7lVRSG8Tk55okz
1dTrpLrrQjkHMgbhB4YY7YpDiIj6CsgjZRo/wImZQSuIEwk31C+VZGZxZwXkfO8mVoi8J9fNEDu0
bVQs4Zm0Cov6DZNBirYZi7er6ywHPKr7QZnsDI5LFpTJZMPoRxwIttnDGg/RRVjkCs6VooEeYQFl
04bwY5L6LkprlETrl1JqVS5vwF74FAnDqjkyEL/ZeKPr5kXKCGGIIBExCLKYZTF4gV1j/AevChHT
HzIr5Ma5iPaxsqt7iZ95KFSFp2ZC5b7eLGgPeohc2VGOCpW7s5VET9vyBG2G7MQcTc0hWQaYmA0q
tu81D4xK3WMyk3LK9JBSGs8QpR66U355ANqOMLrMXG6uq9lF7lbiEjHa1nOYTeRmwpPcnRnXFOCl
CeAT2B0zPu7Hd+ZbQ908+CM4L5gUNsLZKaz9xwlwa0J4JNB7pk0QQNxSfj1L5s0tbz3ZxeYNpehe
sN9yTyrnxoBWgo6Gv6iLFciIBjbf4EBtqoFlZ6K89TUSXmjuQdz7RXD4BLawQiGdxC7HlNmT0j0Z
iRlWWcWICYEw+ww4S2jG7KfgSch+K3X/UVn0lFW0Wr1gwUf26Zfu5v8n51H3/b7wHsSYUO5/tUYG
0DyNHfuBP9rEgFbZWLyV9ep1M3moJcmvBPucgbFTH51fhLJZto1nEPIdfzhYhGoyiYxUUcRaVy3o
Krv3Qmms7eZqDEi45RNTlWA+0s5y5TTA33iXbKG50s9VqsgxDx5GN/SqRuvbLYQ67ipEsKJ5rUV7
uagoYYcGi8B8UfLdHJU2XJfjU57uv/o1ghuTSegm3gizEf/kwwLOnHABgTyNAuC4nUzQli9+GOKc
l1tvgOfBJk9s4NBkpMk+P6NMBIUlNtpGIwe1cqP4+L5YwhqRbCZFNNzaLM1aXSIbwlD52RIzYIaw
NfRCvK9jVOZxqQIkcXqLNjqQNlFeLrLjDZRXRm5n1LVfHaKJFRLf6l9J+MA2zjZ+U1U0VVXVJ4yu
OTUgTTlucQ5z/juTWWpR/YDO6lByVfpDG68qtZLWDBFLPXUCcYdGw1X61g7FOwkBJDVoKytuYSBr
Ln4qKjzrusNeWf4li8mPCzdvrBtFmUP9BEhK95czgJSXUCgxrm1NOAH+3kO4teuy3lzOZ+WpYxTz
lXbOjfP7dWXbLQbDA0+Fh8zCvx+OQnlM5PK2lfxjTNLox1oHcBudbEqVl/eRopFC5y7awKRztwww
GO21SwZNSM3uHrtHqtpJeRaPiRTY/rwpE42LQxpJLMlt6OB09xYX1H1AJqSaFEbbTOJafT5I3hXP
50JkxidtX4gcb1FALtDfEW5yXGkX+gQSU/vEETaSmO/LOsh0zjlACAEu6vWrGWt78k2mOAOPqLBv
iEKP6nbBoZUrG1EApd4U+ikljH8YR1vnvOkp0tWTX0TQY9a6krJU9kjqtDd6fzkHLnLlidiqVc3a
Ax8a2m5KE3Ejta80QEF7kGx03kLIAGOUbAkZEOf7cevMDrEfjTzPk53m8gmUeWlwhZHpugHPnzHG
e4nuiDX93uW81xpWT/d0myxAwdAoLz/UpNfV2xFphiEfMEDf/Dy1kpKUbDkEGud9xcWw6mY9aO6r
cuw/iXUt9AUxRWi7kSyyMmXQYfX/HaC4pjYZa8qtus6xVtW+4Hk5mnlfNaOOruXsxaznsy3A1FaO
g+ihs3acwqCI++lFkElom2UbtG7eCcDWi/kg+QlHcdOkxZCZyRmwniDctt3Ejq9vuesuLmgcO9pn
IYltOfCHfFzVH2BqMPUw/7ZW1rFdD3fMiKdJhq8xoZfJx33naLCufIm/n11SB/xJE82K0ol+njfg
ATcLXOEmBx3cDC8rhUnZ5imx3ZOKlDEEmafl/pRg1pz1MoEDeAtV0jhZOJ7R9mwJA1mBaDsiPxOV
joFltlxGGdYgXE1A12h94ZiJyrNqcKDLwlguPLpxToQeCDoDUzRthOZ22eg9ZyvGs1Ji8zNnUsGI
oQ4XXfP1kvwn4QdwfbMIifAPL6CsfisGKr/Y8RC31jkSALc/H8tXxrmXiJEwDOAFq5vAgr9GnOUu
tsjxI69R4wODtXMTXIEstq7GmoYqhnc1Lisdj8QQBzYeIZre9EouLaUIYnRt3LMS0ePC+tNTLFfB
hFHZDOtIEKwXKUapSjBe5nhhP8JBTQp241G8zd5F3LHy4w7pUowgKPgvxmZqkHw7rdtB5dGErpHK
5W6/iBRJB2oNO+7dusV6ChCQVEWy8IjqFvpVleEbuxM4aV1VsuhP7UO0vA94T3s6lLA3HmzqDI7i
tp0TtYz1yRQeShqlFhuOLG4NB3CzHmm4gNkkYF/PIPQ72ExGnrtAkyGJvFrweyl/PdpZnSezXjwH
V/foLg3myQP5XlP9/17vIvhuFx+HLVLm3lIm7aYnDd3psL1flutsRgql8sEbBsepPSbKVtpme471
QH092NqXh07nZAehKYpulpHErnsqlhrUftuvMGHCGkyjWYH37jGOdYz6wU9+EhTjD/dT6R6mv3Ht
XHGYLtEExJsX1/GOoDh+tBSGXp51KKF6edhhTWFs11GxehgqTKq9oaY3y3EXYfNq3q0+JdDjmhM8
3s9A6jtajoes7ngF1a1qQiYzoEHxdizwtQhQ6YC8rbw56bvYFVJ/YTLkoXYleiljMhqQnvS2mQnX
JRxF2ERxS9/D/BbVYBx7mBMQJlz++i/pLcIErWRdXbrEHUrIN8kRTu7byq7II45XddjP5UVn1HjH
segfS6vX2lNGs0w/Nug+Ac2Xa5Pd5wttMztNjDJLqyQhifmQwj20KS59SVnA/9GaC2ZJuujVl9et
oo2Q8N6nro6Z8z8AqPoXzSN1Zj1RzFqkLkGVfPuz9AfiJ9Q/fcSeBpQKO7gxF6rqTvG8G7HciuzO
JiHo6OOw1XxPfjoGol4HIsaQ743Iu4Q+N9hLFTtUIZ/v2Oi6WIuqumfEcaYzMcN/2qa43wa/V9BV
OqjjxLON7Lt1hp+QngUlSULm7DXvlSdeFbg3zVRmnw18hx8ung/lKx1LiwQHz6cAa8DC4iyOKq4H
rk0Ylt2laozbIS4f3OvdjeaU4AmVn49FfRNkwL7bSXlPQPy3ySiY8AXqf+ERKkfzsok674wOYMBu
VJebiANfbCo0du6vO9GlsGdSJ+hlTV4lj2MkWe9F0W6qX3NZERQ0df5Gs3s/Hdig1AVuvzZpezbW
omnE99mv74IdiRtg9pp0wrhoFkanThZHWvZ/ZypsRP1OLjKe4UGIFpxj8rhYT7SM2c9tA5tTj7Ob
0Qn6OA7oATEEQ/OSnYSuNV0PB4MSC7fCJPm/c78FEi8TjyxaHHUqIXHU7+ZWXjMN/NuqrCXFo3DN
I+td7zNtavkAPCI5l8BBy4UfFyLw5u6ybbpRejR+kUMFzqGnEGdWlrYpEQpV/sSlIQoFLPRIUhIF
EGZrMRVQ83MBIEZ5v8sjt3Cx7BTSdDWihBievh2AA6QVYjuEmi4J8JJ5VRGtLezkYRNCZhmRwl8J
zB2k20cIxbmwM4VJt/mJajBlAXPXai9MHWLBTP53uVA698AFWjmPPTnsK/bM4SrVkGZdV9QAIc7R
gf0pXwTLlpTJfmFBmFscvCPLfhv6+r9AdolDZpsmaLmEEap5/M073pZuRflB4j4N52mIFD74pdhb
NlRSiv4hqLUzDSLASVWji9BpDGcBraJE/PankYGqylXvtkcxVhZ9610HEoOc/xlcrCnoyvBCYQtU
jeeJcOYGu4t81GCAr/LWcIHPuSjMsgWrW9mY8lpvQL1g7VqyfhmJyyOiyKFPlS1CEJRRieV5pD2s
2uMlQkn+WbhOeRlwq0qiKmbgaw1lrVz+xi5jJC2phhQGxANl8jwFixJ0CnGJCcHpWv0rs1iFAQgJ
DB7WQFTfsEHMlcohn5VLQnp0BL8qG2HAvaMufVKoOF20aUGS+OwxhwK8MXOtMfDTYZC392bYlDOz
PyA9/qlFCORh4k0adTdsMV49PKfNI5XQcCStK33a1bA2cTo4jHpPVUXqfuV5BB990cA9n+t3jT2n
+t8GSMY8JK3TCCVFxptu21lRgk4lGycc1nWzLfb6m6/bXTAenOPwVFX3O1l52TjGUlRwL1x50Wes
/oDXYDXduZC+jOFt/4dNt0QUrlKZ3YUikhZikYhBjHBETCTPJ/porjHGNWr2X15ZRVLWRNZc7L7q
WazCY4awYBq150haymU7AgZyBqhi45gDADW5Kj86mUEM4gkdWpM2yOZQ+rhFRC86h1/PdSVfkf4m
14AjwI3whQ7F+foEgP0hzzR7ZOxXaZK6YTAM90MxKh3C/y9tQNvck8UVFbkFsfhmO6O+pEB8RCUZ
MYjmePNUw415Jbj0jlDbVb/LpDW6iL4EA1pbwjU4NCOxCwKxvSCURJsUE/ffZ+RM57Doiop1kS2T
n4v8WM5mYrb/srL+Y/s0hR0x7YKAkdJg2g7TnRpn7zwx2KHd3mWoJZ1hnHmpI+Y76ouH5Hy8nqOn
tSlz7KdnTYutnqt07RPNYPPxprDgAo/BZvJG+549hSJyXKPhxiGUChvRP983nV9p3FzaZQRK3WHN
F3+2vFqFPyiEq0AToahxjaLWsJmjWZTeft9Am0pqryyfD9kzadcd5I9C0oFrU6VqpofoPKo7nyyJ
kuEOn9DlIrkHCDwcbc9Kct6+g2e9/ULiOJQ15DBM15RnFk+HoJ4DX02pdaOW72NkXsV5KNreh7G9
VBwPB6VzydYh1TYcJwpGdJLJOKCb8niyoeSkIs9/vrw31o9VH/81djW0Xsvd+F2NoneGVg10j/LB
IBdp/KPzFHt45fDhdV0vQGB45fnF+4e1Vdy/CJN9MzhIIRXEwIIgjFG9PkQE2egq4sBv7Crx43mR
oYSVR/AA5jvProCWbEzXa8IKoVtPi1+B7TU/WqdTrS8RqHcOl5w/fUPG1s2HCGSUM7kEIbQafAv9
DLxIAauBKTptYzGwUZU533jnFJQ+f9J/38NNXIY9xKFabbvOFyCmWhEGiqV/vC1oxG1MEmg1mt64
nvQbAIi+qBSPRrorj3lu7IzS6OGm6+uDLluLeikICSqMQIjVZS03zGJLNv2GseIr8oKj+UJaxWwI
p8zV5LFxE8UdWzRrvqHB/QEhGo5r3w1QwsabvrxDR8RnN9KH8hvPIckkRsIhnCVim+PF2iecf0CE
SmTalr13ZOBXK3Q5sLaIPQc4OUcTaHnFaURPSkphPAv7PHnFdbmSEPQWchj2KGC2ZAgoasTeKmhf
nt54PAcmdEbw9rA3Dw0L428A59/fcw7HezD75zAcWmY4wdNQZTW/IoGKMqJehkqn+Etf4lwf0ZNU
qWsQdzs+hHkB523+jXXCt1F+TNtECTKXZmaH+KFe3GSUn9LZvpGzVPZyu0sm/tWbBN5Gd1QreNXc
Cf/uLo+d0DykbprKEX9j0rjDWPq5Zd07psUzgIQbX6xbVgL5Linqi4w/c+q3R6R5MOSXryPXdScV
9fbw9l4ni7p6LNiBLC9zWB01F56s1mYIp0EVAwvDHLgXnujYxNEc82M24/i6+yAOlrLsYNMEjFU2
+13GSClztvGytb+dX03PN8zua7qxUV8o2jgsefKJZlM/hLbNbuG1foP6+ypfa6BF/0DVk0JWRr/2
1VEMgEjTbw8r4OUUyXBq4VFdgDptbzn+Trl0GBsEgIJCWUV2t84p80jMsRz+hCekrwDRKp2rtEiu
/IJsUcEU5y7Qni1tfR/ih7uXUPFZZyrVju28D7SLMm8KFXNLpyIH3VA5+bMhyZGi1bq1HTGH9yS5
JtszV3Six05a5DY4J346gXC+SclRTiy2i/hm2i/E/FDLvriblwpk1xT0llDbDL0vmHPqVRbVrIRY
rdd4Rccd4Q22ksR0RB7E66reWpIsBhFKBqRdp9bjlfKZgDGd7iyQFQgxSQxcMqGUX/B3RHoN6r/Q
rGy6IZy04Svrw91tVxNGrsbDkSXHfbdRCwpgXGE2ZKXBDccRjWd0ujIBjWmvkySUdg5wbuy7q5Gd
OpsaTSjN98XMFE6+LFE9Bf+Ug2BiF3wwQ7PNVLiuA1LkxLG2+SIVmM5nIbKC2vTcByViILkxRXS1
dt80IPleGifqgVMFfDyk0mXAW9ZNsSNLNZ6G4616X8RNjKBzh0dpb9Zfo0ULSUtLQHE+IHfu5+ZS
yzxnLPiuthDWBDJH54qqPK7AKg/Mo5K05/7umVhlt0F23j+fwP61j31y9zkdDgX9JZftXvq5uI2y
jFZrRiYtOPNnKiShGZ5bvj0EjFJ6/X0ban5he20ABYOEQrdiLKeAGubbJpj7/2JYulrrJHLBuNqx
x6i+tiB9er9BFoK6ik58bkAM/zA81T/Kz1AvQgwSdEHI/ovJsO7aIvUvPvzykZA1h4/0RBVxNFh5
gE1WGUFVmNGA2wqb/l9XcnjeizYTFl3KyLgV2VOTFHLwiRT5JM3Q8//MgzF7K4D9Z9p+uljd2wQN
ZeoH9s7NzSQm3HQPatypFDW2rIKms3eHcXjy88GwbDfGNAEEHOBOz6LPmPhM5gxu4DL6aLlNWtJf
ad+SLpgwmEkj/zBfBY37iX7pXiIZk795U4lH+4wlHk1w3sxzy7lR0PJgqzl8ZE4fR0y4NUjlzDKj
+VBuF6392aTbp8DiMDTlRb3fSe8ztAnxEQyUdcn5/l7F/DERrzFjUmoNZBwp2+fQqndsdmutHQge
UUfm+vTIIgzXHd4Fp210Z8ABNrUpLmz/+WPU0HqH99ViMu+QkOA8n1tBTSzRxLPW70rl5qWXUxM7
uWj2KEaZ1iTAjpXupoP+uNSifROlqPAWQ6BN8Td66D+zHQ8cPC1d9z6YoHvj0qQlVO1dUu652dKt
pXYFqy/uncgCR2mTFHNyc+Z3JUTjZE2S5ZalvACcor8QQJbnw6CDtVVuF4njVcAsRkYyNjAIitv2
sjuwsKu0BmI+ycB4p1OY+xqlhmIlRIhhmuWiWspec2QlT74F5iqSwfGGZaCsk6jEBiCY6IwMuRtu
NXCp6yKMnjNe8l2wevbwi8jVcS+kLurbOh0FEiL1vzSWRnqKTESfAB6ZAifuoFRH/E8aD6Mx9+jt
2xwnzA9nQi0jzBfxIfccgy2Gi/NriRta2719TQ33pwjsDceTJltLboeAjziV3mPSVShycyvMLJiO
n7wo11BbySm+nixwBhAOs6DuB97rj9ZqX8QcrnjRAWBRob7ijOBSt3XMWvLOmEz/Z1pQPVWFHl8+
fvh7kQ+Qjvw/VZpplEEcdq2gAcZM/w9A2Wo6XzdB7JgGObAIQR2U+Bx1mgPjBVR2NTrKjhWpVcVw
q50NPcYlA0bXxpjQZLGQJCT5pyVMivGPcuabjrWUHj7h+IQG+RcQ2YmxKJSHsArEB1rnCdZH9s7R
eoepOdZTzKfNVcllSvEJhtHkNgqy7ip02gX/Yozzi2x9sI41jLrFrSilBjKS+Hn9HOKBdr0Kc3fL
/vg8rX7+Id5Nx+r9QHtN4C42PYjKhdBEUsDgqFVm8BgCsF6mKeB9ZGRrSU8/PkaKAYjsgLV1g7ax
vYD6+Uzex9pijEIo0KUAy0J7+FImuZ3tok7BBCtBCXYoZ+IDA4HmvMvTOPQm/gKeMKgG0QkDT2LY
36PpiFT/UgC05wWAY4OL6/S1J7dJrhYfs2QZn8VvnOJUECsnsUSg7r5sdboCOOiK6gT4rZWT4uRg
KLcDV3dcPdVYtTzv8vrRmR8nIFWqiwIR3GT23twnCnvaziXTzz9ukMgc66smFKxijbx03pal0ZRI
q8d24wVdFIvI5B0rJrC5027gsPZN4Uk7hVZpxyVssNaQ29jHtjeZydjsv/oy41YpdDc+BdNimDWU
MO4mXMdQD0uaCSZKRGNkhh3V0WOTB6SMTKA5fxas3NHSueLNle5oBmKsbAkyxBKjqp+2j1hwoKa6
8nsRLJ6TXqQ1La1nou4YYmGNAP/GJ4HkrXrSqxFhEUekVVEZof30Inp4OdwGtgdITqhmfjmObssp
H/lKhZ7gYsAJVsYqc6wSWOiE4Q+HS0NApm8yZ8oS3wip7TDDLWj34B+4P0StplltwThiwmdeHryp
sf13OL90wC5xWd6+8FjC8VNpyJJya6Ef7J+fCs3Ylb/AlJ2KZW9RZOwH8jULlIS7Fhuq+dZYNCsp
8M7YQg5zRl8j/PRnncVPkF5LS1PmNe5/9MjLEtSPYWRmIOPSJHroY2poW0iSjJ7HQu4LFOOsWFap
IVWNLs7lQRjMmHLFRhmMKcaOrdC67GGw2y7n2iMAhzY7LLYl8gbjN0251tqwJUoe9b/X7mG+qwJN
LwNk24o7S4hhduI7h9kt0wRSCiebtyQXVI2UixKyJ51KrRv7uB3Lx2rb+zdpxPVtizY2gpmJJ56M
tgRNl19XjUxCLS0+drpixsxyFsvemYNMlyPAhI+RWK7pbP1DtEC9wtMS/xg5XtnbJazgDuIlm20F
GiCPeFCT/2zsy4R+1Cs6YQ4wDDA7h9PwLp+sWl7Se6JK83sE7uXMyVtBKmAaHVNMW4TTcEgVNLyw
SNvnKovM6KYPGgDZ3lAuhaZRFNvaFf2s/7DOQz98nDnTAWl+PXVmq4d1PKMy9PW93XWCr09Onihy
ZxzzGcz4lIqMtxhFoWwl4Z6tGwKmAbvm6WKVJyDiQJV9qVUVdRr7IJ2f+mJ8ENyLoL4qNkpxCFdG
z/1MUKxJE3IlJzZw5m6ZWkY2eXGs4kMawTDRFl6eGwUJXQ3gsN9h7d7BmM+t6qQBFdkP7FU17RpF
WgBujuRL1RkMhs/KCLXp+N5v/FtwyNQOWEeJFB0Ln6D85lFDH5kMEVo7q2xElXHb8q2e0mP3Z612
IELKFs4/ikQo3e6fwUDDGgD8G/571YEYQWftsX7Gebkn/jazKcCeTnIGI5pQqJmNfanQB5p1n2dE
UtPIRSd4J/fCA01RA/87oiMnUCA7+ViErLWqIqjgNJRyiEZThz4MGPT3khxlhOp2eIKR/1ERip49
ew6aO7b5nM9QQ+TfrhyUd/4ZMO1OXt6YYJvGkiYP0r16ns9eOD3Zvlgo93Ze8gQi0TYn8HR7b+95
mlFI+p8RB13H4x2iTZV3juVDViQNSfWgUcmw2S11YDLZm0VsGJWWe+Ery/i1Q6jnrPhf6IORATk8
ZznwGr/EAGCCf52YrCCbrP0ht6naeijt+GkX5lczfmHxfJMKIM4NiVs0ek+VSfqqPbBr9A5U9tWV
lxOjngVggbyOJgJOrj3CkdFoekAXqXnHvoofFmtAfGpt5TNOnD0HOQHhfL2q9AHD7C7FHhqp3Xyu
IqwpbEsLom711Vv+JCB7o8Qqzz2qCmzj58LII1XP2LPdxB3tlaTG2/zUVZhWmQ7h4FgpIBXNJT4d
pTvjWL2HMDb0krm8jKl9EJCXTewxsrC3En/yDKC2VD+GPxvSTHQMT9aXqMCbcYwx8u19MdbVmlim
pZhn1PEhak0YKzpXvZqJV6Fb+0xGt5NrSXwe8S48D1i8rPGkKLc+Kjg6wEEtrVv5GWsLgjZv84PJ
a5dqd82SALz4VPmskD1Q86IAW7HYCVOPSKly2OHD6hbMoOW1hEOCV7N/rNRC0pX3xMZmse0bSroY
hQlQapMAGiz3V5m2jkdEgKBp5YRp3i0HhNSUkfhP2UgXiWQWVSzpxROU7p6DR0PDDuHu59LTlCbx
YV7BRO5fxx2NQJQ9bE8nx5uiz2GavkuJc0zFjx4AUQayAOVoVWESrsUG5dOAGcAsdkPK8KfKrUkV
lKuq3kjfb1jy+itNlKZNMMVsPY14XTL93dXLqu0W83MM2+Xuv1Zt0zs97THT9ma3eEmDRC8zf2wd
Hb39yk3gJZv64wewIANNviDXuu9V7rw+f0KxoGcZjrV1IL5h00NcgDgTYOwZXqzD519SQrjPuY2T
UeVEwD04RRlIdzPeHormB1uVgshu3R1nrBA5zhghBphQpiDF60871sHhEWpHSrjuL5qUQ0LubIXm
aWwNNZhxwnuvX8YREPrGvQtHbYHXgja3ip/pFo/AdXKpiYJx8RQZdr4Uj1wxWLOkBQ7EvVVWkJbo
JA4CqhgEmKt2lGzCxWXpO+oFB5U0HAzGNl3laIu6TaJTXXAMpukJsw/eIHsH8Ff8M5ifY3INvsXB
/ltpw8C4Ae3sVFl/LLxYdLe82LIwkqAwAjoQtSEqooMERsaldx4RDduptCrNYF8COHuXA4qwn889
5zzezf/+OJ7XwPx5sMy4QIjXa41ifiveIOG99gXAqFGkOdpG70y+t1+A0tOpi6kuEAVtr68eP/Ou
yNRPIf7931XhQGscvTQvhpkcMEd6+sty1EWqrEJbCtgPbExIkRfizqwXQewyLg5GXiyv1B4LwVq1
le3zL91Ca30jDODbx7OVGjUCf4vl9Vx+sKdEAjMfiY18NHq2riUTlbWrPzbGhbsFyrNDTfJYVafQ
N6HQipAjWWtIQFfG14U2LX8IA15o3yWimr22RZZI0FjuDuIBRcTbGMSnMwgmNu5QCN1GaX4YitVm
PtaQwZ4QtWbsn+58u0cA8YiABbS+XIya5R8kNKx11hPEnO4M1InjONdhS8QxFPTn5caIERsd368+
mr1frNdC+j1TZiMGtYeTobF+W843lYbV5xD9ot/gv3p9dCXwlcIGokGpd+mQYDV2/uI0RrZfT5gt
v2yEszu5a3UyaRhLo2sXaYZet/kgshVSt7zcw1woBiOC2J4zklEn4G7ycoPVG/SdF/kquH5qlbkR
ghIDJSPprGwQjLVNLty33QYveWTRpc+d0cKMTj39jW29SpgpX91Nhiij5Xw01Zq0cToWJRflaEZl
hjXPXJkAZgBkwxLuNQDgqJcrSLk2eW4mT6J3eIlVmpRN6DDE12DL/nIXPXwvKct/9HtUh9JbyfWJ
xS2gYsbPaMyhxrLAi87EeECEBF3AXNzlD6pUXcfTzE11YwBrK3Hcro3HcAL6ql89lICHVw5f509D
oY3jLMzDtPf+6HI+ahWn5TlaB4EGLjVXRAGgAsKfPYhPPYVK7J0MqKhnDCvx56zxa3tGsfc1ldGW
zE4CVXrTifp2FlYodATFqARMaFoXZMLdUT8VfkespiJ57mUhHntZp4+pulRCKmrMJKgto2OeKb0i
wHNpMGT5N2gnEInK6MjP6fgM/fZtB/isWS1f638gYj3uwMd+Htl19/KQuYANCmTIjhDi1q3iB3mw
9Gt3ASkX7+mGpOnxKJRc5pPrRur2DdtBBHTvUtK5IRfr6kdlzlCaZi/iynzI7DCx3i31Bioq9cbt
Y1fJp2sYEXZvx5Pf3kwRB9NpN+yjALqPkML3PrzZohgNmJj+Y/BPwpHbJQx4ADm0IgtHpE2CAgc1
cp5tB35I0HwL7Zi/tKNmoSRyZszFFkxjMadNUOtrV0b0oXE2W2SczYoo8upWqqUwnrtbdZSMN2Xi
W4vYotyD6d6IN8yjvKevOs5OX8+8tjApTcBjJxPRCxCBH+g2m4IitL8+8rER00RjEkTDqXFiPBdL
0ioj+JiP9iTFG7uKjoILWOLfmGvlBXKp5ufBrQO+Siv7z7FRczokLTnJreTeCowNHBywJI+nPfEi
1eG1h/Dvu6BuSOkSGDCtABuPpXE8l7SKh7Jt09ux5A1WhxNI/HW4bjK1MIKBMt5t02jVwjZj73wi
7kG195PqQttQQbuE6+08VSGVqcySY4yzru86sZPvl2raYeZEf4DNLtQ4A4qTYs3e4kYr8CDLuU9k
I5l245yOOzDISfo0kIRy2IRg3V0x/xLBHk3JPPqDwW5p51kIqVYHuX8BA6Ull2snJ8iAvCnBVglH
sDh+Bv6mLxaOW2qKqqUcSG7ycUEB/juBYkca/wW6Pm1NxrJPjGnoSXFAlvwxNojpKeMEsw5mY40A
tvhNrtBzev5r/C6cNzsuhhKN1jq75vhCK1jgpUYFfS+c/w14kvToWkPMyc0ESbP4PHOqViSu6OQb
LtWH9xLU0jqwKd/OacBf+1TNryW55j8iw0E8snDaIQ+AVXilRJ9VUDYIna0EHTdE4OGVZO6Uf42X
lHLwHSEiue7iF+uIee4FGy5pGdM8w2mc5CC9UvFIv7yPAbJXpPfeeblL0Rixu3bDbRIK/UqcC//W
jLQa/aabwBX08FV8eS/yqI1CaRxvnJ94xPiyhlEojHXwPogsogtsN1J8TDlnf/2rY1TEPzHEZpZR
l/vJsPxECgRAX3++A9ZHTbQkiNz/RQkyQ2ZE3/jY224IijGyrm0bNvX8MZA+U3zKScv/QgnlazE5
vkZVKg6UcxCOw9J1xCZ8HWcsdxHbSs3YI9X2rmiPEEIgAf2am0Vco9pj47PVUNONb63Bt+qOVvDA
gNBVlQHO7c1Pb1QM/jNP7YO/LPSbD8Wvm6AUeCX5SWDaBJaJ67dFjSWP31r8wugBNmZzqeSChsbJ
BOhH4e2m03qIif/4Wt5XnokxjtwWNvRCh6BCwyRDL3sSgsThCd/Uy63EyStIln/Run+7dT6Fdcix
/15N6u3lDjZqO7gD6ecqUI/2lt/Bn491L4rMXdGzMYAc8WZXLAr/cdtkhSTVTG+HPXPCnM61HqeX
STu7b0hnapNW/E7e++lFwsmOUbSJlgitFfnnYxAemzia6Yr9mC7Izx6DCIZl1RssaKEUAmsDZ+QF
pb06M3bAA6VfT03N9LN5oqyjxFGrRTiWsgJzITlyid0NYhnIcOs2LjmyDvoK+2ybvT8rAAUttu6+
/aDDh7QVXok5GCqYctMVmZWpBcXldKqYR42zESWVHIDYvHjpXQzAV0EyU1qw0mISlZA0KnXKhWuj
SdCSrRrnF1nEQLE9iEqTkDLCtw5v0KM30ZPzjsDgWkDFA3mmX6CeZVX32ASep6vTPx2BGBmqImTm
cMd7LFcvsgMFdNs5oowGZlY4etsSG8v4BHhC9CFonBxuQyZCXEkI73z9praoIyN82IS78efiNgZM
pHEuBVK24FtulwpAztGUXnmT+1C76KcABwCRZaOVvJzgw8IiFGN1UAOHD+s7r5/B8m4HhhezaJ/o
KglwOvcJrCVglUmeW+nP2TfzGrG/xkuA2ULb9ZgV0dClSL2heii6rf46s092oYgKDFLy7M2UFvgj
o8zXBtw/f7ZTQC5kI+cQUNtn0go+EyUitzt+FzWAHdWYhW+uky9YqaWZ0V+XGWvuM1k/roY+xT2+
W07DjhgG9ZSJeuepknJdOzN+8nJNGMWLidsl3ogX1Cg4foa6mlpsonQjv2bA98ftjeMJDpc8lw+l
MjXQRnzWOcAinYbzJWpGrGMz0MCLM6JB19FbDKEeT+l4dhJRxplBBYWqjGis8JSZSxQqFsxJRmc4
kscT1ZIzDAnTyx8uB0e2S73rk+jN2rngYZimcAtrgwrNBnpegSZgjuK8Md84UkajZMTF51UjT8Yo
x3ZF57Psf9Ve3HmAdvKHM6FHsju1toio/7cHJLi5Or4FDTRWhr1wS3+v4WkuHQL2VMYFChsqM4Q4
D+3oIDkQNBjNM3VFSK0+5pPKP67pQflTFNNJ9Z3GUmUn6sCNuSICZtZAyioh7oeqznJGlxGljZaC
/ep2BAWxVUNDJOaT0/f2cABkI9wne4pwFGjNZvMyel+td/fNkKRW3ZSw55yUXDf4idDtXm6L164m
n21wUnV+8+MVk909mTj5D8xHiQU84DOac28oPrdKveuW0HwHyBy3YaMXSYNruJCruKbGbEd1bz+6
1Z2apYsJEBdVT8zt/yEshNiRGN2SdmkVFfOBWTluz8DGSHXiZlx29wCX89xZeMx3ntRj3s9std11
jOKufJVb9lfgJpXrL3NqTgjPPZFHkpc/co2wpU6bE7seaEzGqEe4oyU1AKp5SknZejMN0VaEk4lS
pXvoXvUXjhdai2zkrvgwVYulxPRQxz8j+3UEV7wkure4sEQlEP2y0AnQv1GKOfw8MjSfEymqHUFA
pqhke1T9fHgiYJCkWqKUahp3bbJkpeaY1T5gQ4XQQKb4YibCEZU8NavHxjyl5IxCEqpTG/T3oUAg
27ynN8qurXD8fpxf25DbC7J3wjrG7KjUobRXhXh9vpbzDjoGxA7WDdZWbBVEiCXm1yZErARG8iAt
hMV4925arRZuOc1BaKN+q9CjkYNduidB6ibDrhjneJu2NsvTa8QFZcNdmyhm1lmRuVnh9or0UFNi
KOTHzBimbTgHEmxqPVZEiTyzc+c3Kd9eGMnhM9BtABzEgTelj8feYQCd7doYTbwHhBP6XwTP/VAp
CUaz6mzixqkdHKj529/G/luEbXqu2EQrRfhy2qcPV3chzJYMtjO/YGTmYKfTihSWDKDEOmtjAW86
1YpHmhZVKimG5EKZC3LA2J4oULm9Kjwh+iO53OQHwZDLw2833nQsOlgVcSzuGEKO2/vToS0pwqRF
JFuA8xTvCl7vs671wErqVdJuAdUuwazEKs9FT5Y2Pa7/4c4vV9XLQQRpF0KMw3sxZSF8oGW6quvr
Zlnt1rDkw8bLDy5SNCe2RIccHyKNtCgLLMDrNe5M7TJGy9fr3ttCjWg2ZU9gS47NgYIxYKxLMAe/
AJ67JbssnUE5Iqa/SbFylGFydU20LG5SOSLLhPUXzMJb4a1R5J9VoiWoxg6edRw+cunyeeu258w5
68HGnCCZx9RfTA55SCVTYf30wMYU+z8ifw8v/ZKMuLRtJq4lU9gaQrEaNTuAyu6qYWo7CzR2+VQ4
CTyhEYA9b/QRzLUXWR6+o60WGgQakEoG4C2M3ms1ajG8aZpEU4PJOge5nus0+kss/b5lIyWy0Bhp
fvpaTnyBlGRvzdKtU71+SHgGYr8/5TieRCgFxvHZ4sTwKn6Za1jWRVFUwQ6gjX3Oavrbsm88sMMo
FthQ2n8AHLR/S2IH3Yt0MvdQoCVPbUk22/D4ObZyv74MbvrsL7sA1/N0y7RacBN5VG3WS0639kqJ
vK5wSwLz4hpLXzjpRHup8+D2ttqvLgslYg/2QnDwb+ppovvmkwQGUPS7+7572Gw57fSZ793GSIYb
/XrVU0Lgre3y+HMIlMf6EVFgTP6qvdp8hziVbz0GUmNnvl0gyRS1wbeULMK3SYPYf0kcBJwmHWdP
JUuiyFJsqJptl5AVT7i6wsRGcDdB18whnvGUbfsXK+/hNQkQyWyjFbKHWItBaKBKo6A3sQRSfv0r
vm+2tBJbhYLyLszpHIg5SRQjBFvS65j4m8OMdOSNYP3Wj1RVbOBN4G0VP5/tAqTK/T4Exm42bYzD
Lg+jAxES1Dp8M9CKW7QJoynTROHfByLDBTqOyYGjqH1o35Z+VvpJ6kXXn/F/fod9XaGahI/1KuwB
KOrhO03BvaMzEO+OxQmkLxIIfawyUCQKUEUc7ocL8e9+1RDB6WYmV9PntuUoB4tfGjoRl+H8+Rxn
Zf0Vbpr2bdekX/Sqw4nJf28/piGcMOSAo3OC45RGFldK1XwNrKkfYvqIIqW3R/w0O0A00us76KzF
5vb4OXyC7TxC3vJ/qB70bU0Gs6CN196W1h4dMXNRHShbOIVvXxc3sbnAa++4lqLn5Gh5n1phZwQm
Cq5/L5bHb43e6U4Gy3KN1hB+nXeZqSA3ftnHFUmff7ANbGI4NYL72iixaUVDK26i+FJmijVSRgS/
k41Xrr0JBcNOx+h2AX/DlDmuR3rsdx7q0N66C0Dfy7XCn3TWl042SqRh+5uKclE38d5EoG8C3NTM
QYQJclm4YRU2X1bu23jjvy9+pmgqQuKIhs5ApiEveEjn+TXqWuV6gG40KfJENWpS6cEzjy4YnlZa
DKd8ho4jBUJJmJsFRh24x9DEowh2cjYlcL12CbtBRuJo1kVHTQP7QpVK3RM2o5rc8Yf0dpiVmcfC
tMpiFRMVqjcUczSvMB2NH9GleipNDoYCklaWe1EzGsH4Q6QcH8Xcq7hGPkqfoIT6oz9V/otUi4SD
hwNFOek7v00RvugtrZYwTxR1uYUUKzQQjr4QG9z+lCNuiD72+jZu0lHpSYTW7OHjdn+QQ9Sp/n8A
Ttw0xyvXDxQchdM07WtF02nUbbcjOYVR6+wsP08C1E5w54NCG2lMzbum8H4hYtnr6ujOz98bLYR+
9K/yGYmaaq6gz8+o1hj+3Z2e3Y5CT+Kwlq2sgp1MVfP9dFl6ufGOqjijJRfYIg768xVXVwZvvqiu
ZHWDP/nlLJg2d8qkaCFRUWKc4cl5lC+MSCiq/a9DcRVOXdNFszEA3xKwOTi0TQ1C8VHlV2L6BLYU
gsobXxwo60hj74UF8hLkDMYN/fHi6TbKf/GbdNs36o162NmI9zsYcgp5PvKlvNrdq6N0M7PdRB77
dkXdwNrEN8V6Zo7+Msp+XWM/J77m0QN3fUBh9SmLwXZykSHWeTtJD8ZVBC1jHcDlwnP+lqxtJ/Oy
n8Wufjjr87A2oC/tHpl+RvZPE0KDVILIHklRjF2eJ8GcnsMhPf5ny3tgJXATH07l8MItF55nnrDM
O0MZF2rV8BcTxZe3XD2vHE1ao/shxSlXz8QvQ0YB6hcU/KiedYtEFjHMUqTgaIL5yK/JWwmznl1T
E1ECRHfR0brb3AlTo2sHalkL96LWW6ZCGB6aNex+8j+ubxpMV1EmcyXoKINOxxWh0ctvJlaAfmqz
ZAcC+t6r7ks72c6Pa54u+gJJN8up4Qsx1cl2hkbEHkza6VC9Dl+e9vu8lkJ0noZf1Ljk/k5PmwF3
HOcQxHNuzJ1OV2aUX4pej2yviAUf4pnCmufb4qlGMh6PwXFXzqUSo2o0I4BUNLRker5ox4+UTAlA
fV1unpOXkS+cwlptVnL4ax2+Mn9oqcETyN5UiW7Lbck7+pGt0aIwJcVBIp72nVU0n3+5BVNo9JiQ
OPNi9QNRkSRWALmbB8cKlQGJXA+eVUGreAuxIUTUs0rJ6IeXu5CS1/whHydCyVXlELsCR3leZkTY
VQQ3Yvnz0GdtJ/UDb6MQ+Wi/Z/VEG7ez/KOGYkSRi1D/kdkJfkH/dc5jTk9PZZPBxyeH8N4+TqvM
bMFJnxTLT/+eOrEADFo1TjWQ2NuNxUVgTRa42BZz6GFISz9ZtNjH5a+BJA+Hh1SqqSOqCpKlo9PP
WDeUhkh6KxnOmY8sTVtqhKysVd+8yGo2gm4PwacmJaS6hAZDEOJ64urX1RiGJoj7g9dM+dSfU6wX
UdM1/HhtFUYQFJYk2FIBCsyt2NhStpwaX92BuBhpf+JM6hiD8/ifhpY5OGoN1TEZMGFrAWEo3ABT
08SKB5yKeGs3SJnnfwPFi7iI34w+m+rosJVYgTcWCHvqm668kIY5CC8aHOXrz4l9vIE45gyVgWww
g4a7l2xqOH1bZD0agBTlrR7sHMmNnDmPkEAhJ1Zod84YfdR5wROdb7C7wch7Yq4ePSQq3ozmbgxt
MGwG3qv6qvxRKpspZlda6HFB6sRmL8vcKSlNCiFUt48G4JfNnh09u8MAwAWbCAJo+KkotcPQtsdO
4ZVA+tkPax3EzNcZdx0Zqna+yhaGKjDnlgi/MMn8GH6PkRjmiadgS4u1HCglNDWa8uTSR8sgjxE4
RTzBsivC50y1fIZf2AoOA5ATIHAMH5GxdYC4fVwVFYRWiGpGOxxH/+4RO9lxkGkIBa6LJ3qzi05B
ksBcBquRpze3cTEJj0/LiF/DqxLCYJjKgM/hZfP36CXYYWOiDjsZ5UElth8P7Zrp7AxfhoCKIaDK
D/deW0GXS7pY269stNZ8zZlXE0qYQxc8YusNkko4GglNCO6Kulw04iJ3jU2APMDZl+x4e7wSz7n8
fxroISXmaBs+SPMpGMEtd1vWWJm/oEWdV9giQhsoLg1y0ci2S+s51aVLvWsYRyUNzuLTSK2qel/x
mpy+91/EcKFVqmXl3mAOxfCw7riiq3/luwqClpABs9Xo/gMWm8cfXneJ+VWl338ncucNt7EpbJAU
7csI5B3PwqmmxzUkoDnw05haFoZY27FwMP+uRBsTS6voBJ4n7qmhVPJaMBt7KmSqEmQ9ExZcaFAQ
iYtB/kjoglpGrYZsuL9e3sdDJ2oTRVZCs2oidxEA7+tJrxwFzj2cLfOtICwMDxjdR7vqgnKQsQir
xli0TiJ99GYB9Mz34NzQFPd9BLW1QxPpZWgt05XMwwhmg2ptrsn4lqTdoFznNK9PCr1+QL8WDKMw
cclZ/prEJ2GP/kkULYwRvipvhrQXMJToLZzILizoreGHNKSdtR2i6pdscvX2kgSpjPfWIeSRygln
SWyl5HTwWRqhuhwxYzBpefw8lAZ2zZqaCAk21eDeFiPKgDcd6ZqZN3NK+U6qBGYPGvYc1LP2Bin2
ILqSGrgw7VsQqOCfOTb3+r4LCalmX80usENo1QyRa8JF5Qcu5Awbgvk0XB+GQbxzDW2AUErv0VYT
cLWExcIKZ8KJJnyxjD8sozLFO9EQEoGvpOVtNZU2IANDadWw31x2FPhyp0L+cMDFnqJ439uEj4R6
4Bu/t/RT+pv3NVsf7SpEwrMoz3yJzIjenctJiV2ZK/EbonCqP585J4CUDRcIKnn8J8pbmx9bdvdu
bCak/S0Ve/ww3AtgixJ3GyI6N2l6TPTC2ldlbWonD8H/YkKdFGUK69aXnEAYOtpktSpNuU9ROuui
fUrYz7KcruBlIQ5SIb2Y4QxhhLhcN3N7ihWauWewoM89VBfJuggy4sqXCol3eli+bjA83VrHdeTH
OJnrmz4aGV3HiLzdWuPxlkEh3Twuw/vhNxJVxbWEDjc90NWNwIZ4W8F3/rmOMngovQqIFB4PzlKy
D+1MBUVR61syykYIyda3UWO7MK5LUnLYRselBAWbymJpAubpe10SdcqGG4iMlxTispF7RqmAmKKJ
DyrtIX9sW1HSqUlUgNYNSDvdBiKFQDWkw1bVbfqQDHxzWYxFbtLZXkTP3sIR7yP6ffbHEfKKGztT
EzhSdconznvy4X9rQtXn4n9StOqw4KmV0W7biDHZkUvXxL3FtcTr1qvFwmSpVehVq8fN7msjQPI8
CxJLrzN5X3MgJNUzlVbwRK+1T6ES0DO0L94GPA+E80eRHvE5c4q1LfFoUk3P0kDTLx6+p7kZTuUL
px33o7tdx/451J07Bnq2eTwIOasJE/ROdmxbFLOVsK+EUGVBtXAx67z2IVtBYsxyuth53hfca2z4
C2QQgIyBmcgy2BmzHueMWVSqY0UhKBU24ar0CehqcOtJzK94kDnXHYN9OuFFyJGe5JtCeZwTOM63
pcQy1zg79U708LNUvV9QRw8Hs4BzagBafJA48at+vVrrBBP1hRWbpxW/MOrNf6JF3pkMf909tg+V
6g0V9x5QkNtEpyvjQGCMVhHBlVBpBjsbjW/IcT4luxm2HwYZH3/3JnTVqFTg4bh0kz3VlqOgVEAg
64Uwx6FU/BGMUWTaMtkxkiDwD3ZR/JoMx1fZQ3ugvibBQiz1xQG64f7km8YUukdJiF8+0flMS7+p
PjZjBs7Qp3VgK7yKbW3WLWCboVKEQ2I7tLhdxs1TmkEB3IZCcz9yz54WDlm6tkKJvTgdd7P0zlAm
l0MhjELsSqvNHMm7UsPvqNIT0QGJm649qdHKvzynCvPSc4skdllLMFkMhjTv8v/Q5wSk7ofAqkF9
xGDdJkRln1wEhXFMOju2EyuZUWp82xwkhO9yBCzjMgj00XUfITfF/vToJWFFvLy20L2qI823tXPG
me/QkbQOkV6DZe9JZtcECdVUC5tx6xpRuQrHK1/iCt17xJ7jqakdPid2HCIAdPvdIVMkL9IrLr5v
MdREaQcu4jj9d8hIOSaYytYYpLVhadqb9pyyrVglQfICJ8Cv6Sl6mFkDgxHoYCbe3T2+SzQ278qJ
WIgWQd27jYmA9ibPjF7yS43Gi9BRIDIuzPKVf5ryecZcgOT1wm8jCWPiTO42+GbQHqpa/7Gb/b7Q
yTFCVwCc9Kuy7xQ6hSzT6cv44igSzAlRh/Xrq0I7HzeZCInQDgswFX2KliyNJHvv1DM2zkDOjt0Y
2ytiKaLGlA7SIjfXzsu7IC8rsoO8MoptGbG6SaSXNdS8B0WwdAeZdOIaDe/ipmDrKcY+3vY250Ej
BCMicmZeoouaRhhgGEMkj4VYP36dijJQQcs8cJlVedLW36Fq+Fqng709ezBxE5u6DKgwCYg5z2pt
KwD5EfZCMZK+vu5LxREYLNLO2N/KVCNdr2UnIJ1vDZmVnGFRcA8YiK9dKsAYvtLVHbnPtDv293iO
r5/SOciSH84n/gsyj1cCeT0vqqRF10oMcCVRWfRpLXXfw2Q3t2L376eWKGfePtm4FO1O6UvbsRak
YYpx2SezdKm8s/vcWtA0zCzLsk25XTr+kwKduEDChjaNON1QRFlrHxOjRoYY077mdgqQsRmIFBdi
UjWeAtjjUEkdvaILhCIgdX4eW2cmnbNnJwNLEQtUhl/lY5AJxJa78UwR9RDZPCJKcuhMZsV1MV4T
0WNvBL+zpnpMrvN4qDHmTt0DmVoHyCMlSewuQVQGtkoFNt+A3gjBQghKd9YeyJyc7Io/pHCHShMp
G4D4J2/Q7Q8BbXaFihUu1P624l5n3Ms/LNKHNHbMglx+MRTan+uGjo8KKdZku6MW/iYbvn5J/mOU
CstSBFnf5WOLbrCgfR4J5pICzJYY86MAEHpWwgPxv4qVyJg7AGTdGcUhZMYEQn+MuIPXDBPzDyNU
xQaS86B969Ad4WV2DMQpkprnOFcRvfQC9nihZN0cdqEa5np4PR+4i02Wc8SRVDxLQlpPi9CJDARo
KfoPTotPUYfl8vIrf+xauYwV+cNtn+Zs+2KG6L22r4L62h0J5ZfXaXqUHg87Bp/t1xPV56rbJuIi
XtSUgzODTjHX6oR3UhIGj9zMD+q++horA+B+yQtp+ewVFrIPaxBO0cHch+eEpnwu+/SebbxxC7BX
wR168UNYTt0cUwRHd8Z5JzSFKNS5NSwMhiO2kUJBWmbSJ/QCU09fn8fN5yxrxq6rjHFgeqv8wmDa
fNKSq+5+bPlxgvnWkOHc4CIJcmDdjfFARlV7yoqVNO7ty1ZPdXGdEPq4AssQ5+YaVRJITOstZh8F
62EwbEYojS/QU0yLg1U64sbTzGGK2vtvMF2wT5Klnf1I0E2cJn3zj1Q/Bx67P2M6exkNnz89K3O7
iz0CkFRXpi47smA9BInk3M9I4EmFOdkYy2K6Cj7PP+n0nYMSLUMoqzgFxTZTkxxENLi9LVSer+FB
a37C7tD3WzhfWJ6DxqGGjSnfEvmTsw4HA9zA3WRr5XE8uCV368RA9CgNqeCgALxyw/ramcLyFDLK
ahNAGmZO5aOlB9xSJORgVs36xDh8EGoYGtAgK5NSoczj+g4OhY1rVGRffhJxXUQNSDlX7SlKzNfw
G86hMcHNu4TOXpr9S0vRBPhTzYU8X8BhyjpZc8HMcQpMERqOoXr8b6z0KZtjm1FcGtjwk2qaGSnn
awpaXDRrJk/eUWtbrjvx6tcDNxn3A3/JqlpOSZcJxn6qomHjzET3JiMMIsTpSYqI49ppTFYpE+V6
uUatdFKNC1LxsaEKGbt2iYzeDvBzbupGD6bYO35QZPyPiC/gt2piJLPZynmtDi+0G605w2wnrR5u
MvEatZrKBJRWW1FAysQ9Sy0XBM8YhBkDRYtoQCqLOPHrxDikl7W5ak6cn2RGvqqAJilAyn7JSTUJ
3Oh3iwSWi9lmI+Qn/rnfnOKGdyXRsm8b3GLC/q9IiIkxi8MpwdLSAsR5FZkQTxAGmOT/LhAjBoYf
7/VLPYPhpTW9/IbjPwbCwtHua8DyMMZJItou1tZvjYhZ1gVUIqBvsvhfoX/FDvaJpk+oUPjTF88p
+qIc9dZ5/+yYCwmbd6GApAezbEsQD5iUrKA16tUiU63Pd8hwcwG9wLPZV8waRWMqBNOhAEeU/c0I
bkeXmXK3b3MBu64BuhGtMttG33vR64C1Cxn0TKRdn21Ju8aoasBiYBMdYH7VWj7kTGmeLko8jTsg
XvF2/HyBInpk+Bw8TIjDgXnb2qxrZQZfYRgHruz6ZlQctix0X3tdlcyr18np4BPC17ohz+sJ411F
/RnTV255tqZwKbkjxexVVbH9UA3rC81mKeOtXeDXiG6UzuC+Zk5PhlsubNSMdAQ6z/NVkvWiSvVz
dFXjBkIZWCQRIer7Pfgq+I2GcEnL+7NhpCnyXkKZBTWit/Pc5t+KpRY84dwC6EUR8Seo58CGP5su
qCMR+B4sC9o6wvyg/7gGziTx2nwXY7uHxR0Dncbafo/PTQb+WM8Wcl1b9yhUjc9ZcbjGOylz7uZq
ewl8XqqJgd6p6A7He7ujiRXl2JtuSMdbB2jtRxj+4pA2+ScThuuAQV5uhb4aGV38xxy3mjFwNNRv
FeRTpaPjtVnO88OY+7CVnpMRK1fVFOE6Tbd5IA+B274o5GPAg60/yxUPoNS66OMKrgVJHdDb7nyg
0nK5fE8aFAnXfBMENEXuIW7p6Cd79XfMzc29fNtfbPjAzpCRb/ABDWcyFeF2AvX6CqLgGfMUSEsE
DpvR+BEH3t1hLodOm86b9jB8HHaK5vnyJT4P17Ii9G/CDdc32TUkYmltH2mMknrzKqYtTCkOEd0A
0uEJLDUbODKHOTkUOGtwSiZxVzz7BLQK0ujX5vKVx1AgANTNhrpXhTjgIYnZBUQjKItdi9enzywt
yW8hW6gcdt6GhOl7yHo+m6e5Et48osqyVVlGXx+15PWwVlsd14WqP8fTIkRgEvwvxn9GZZnJDoKd
paP5/N8VBJyzOQ+x4/MuP+o8YHO/rI4kffiYMh543fuJLghcdMJ89VF2NX4H2pVHnd34NhboEkRC
WuPjd44DTT80OAq0gEx180MWb/oIaphwAkTxd0ZfIagfgUHjj1j4k7wzODoiEpcerByCVSKo3WvK
4asxqq6IigadVEIzfO2IsWI9EC9P1KJ1I+ZatKRlAevbai8St9545d6tfLQmXWUXPYZDz/Rgxf3p
YBjpXsCmlFayZw933YjEh4Djg+J56N40Rxt5/Bb1laxQjYd7eRPPKIapjWvMpzhBlyDSpFdQbJkG
g64XYUC8L51XM2P078nafhUi9zdgqIrIaSUxxwdrxaNX1SRnViYnVk55bhQiT+15su23bjJXSb4p
hOpB1NruGZRRf4SVM6eMGqpJ3eUpXFzmB26hIPjPbr/R5s8FXCoFi49bGavED5xi/clLtM8k79h/
vUg3S8PhZlmX6tYzbsKIYEJmsr2fMzq3Hj+50SyZFK6w6LnDVdHDw85yTcV9T0FmRTWn/i2hJF5b
5FMLfnTTSqNbGZLaiASUQKQgAxHNc2kT0e1vlniZNAI6BoCQZd3jaXqo35sUXLEX4bbAeLq3Xz1X
qgtHApt+qX9EGHWtOJi4J0amZuKRCaC3DyOaZAByHjYB5kkxgjsgk1tkCEiusCq1dY768FPJuEsj
RCodGv2LHOz26KVegBJk/w/x6kimRaR28q/5kjBuf6Op9nB9mizbT10ZhzM2bsQqzbIg1ofYCA57
xMHV2eCLL2N4i9hd/iWIQLnWUqXdq7ZvmZAknIcp5lZGyn3fAMBij8pyvOs649H57IRwUVj3hvJx
/RLCesGKW1FWmt9uPmsIoX1CFExNW/3tsi2blUTnbW2Ubboj7CefnyAx2rRsX4ojEZzxk4zznZ0s
69u5Tv4zG97HImVs+T/hbRL15Y+dap7P7pBM4BGIW75+HmL7UoE9ETBnfDAnM5ufLt9bTFf3r0Xy
FCakrBLtgpuU6zszmJWm/OqUBB3m1HvYGq+tSH5e/frY6dVPSJm3UYIkqFwEyCShScYrnbgQqAai
60tb6wkRP2QHed/O1lk1mvr78P3hG/ql++wRkncE8+Df8GcaxkeU6V0bLzZ8Z9Qs8MeM3q1gMr3z
tHsbSBLzvIej1p7k84zk/YNE383tAGKy9fI34xaO2JrcdZNJFE6U71lxfjSET1gAYkouVg3xJtHT
HN2lkJc4keywHB9t/BC/clzg7dmIRHzi2JnBeTYphYxGipfrhZfl+pSolgtxZ1cxuKs4Quf5qTDj
GCVNwVeuJnwF8LF430dKxP7140rfZcn2cnLkkbRmJVUSuAqxW7kC2vdIPsA3lu3qkT/vXBkrczsF
u7+ylmGtCXakxZCXp//7dsjSwc+JQIF07YO83sZ/nkgrzQym56X+2h/sg3Dj95SbLgyg96TkojgN
J6ivGoQXohDWm5bG9DIBVEH6Nl4NurIwcp/ilif5oRhNZgFHv9A16XzKdoCePo1XNpzVF4fdwwmJ
roYPBos66om52LSomNcm9Wljgpjs5k/WQK24bUKRgOFKxaw5C7QdqeRxhftmomf+Xt7otTdeWyxm
nFu7binXK7htZ2N+i5ouzk5zdlNxAgmW5HjJeJahc/SnJF31bkY9NTzwLUnPDhA4Xp+8zCEMA7ZU
5gItW//GptrAPlrSEoksAVpeZYNLdPVvtSQ0uSiJwWDpyMaoCtCbzgd6GaSNrCS9x5KOtSIXe0W+
OsMnk0GyaKBRIAc8L2s8B45oZciQx9OD+XM1W243G6orkVq7GLgJ/jqzP2mxh60y2PJyok8CzW8v
+ch/9IhWngu3ZZvbQiuk61sIo2J2m5VnlWVgTlqL+INEZ6dd4f59MiijcnunMubzQQ9uh9FtTAxP
nzrO4XUl5rHojfyKips3T3TdAkLuxw7Z1lRPyfK8j7XR++sIYg2BuhA8NiQbFgoLwd2/ut29sfHL
jIUr2k8wWtyRyXyurmBZGoru0Zu9hl5yDs0lTKP4NYcpx6fc1LycvunwJYkoI/qh3Y8Yvp/CxI03
pA5tLd5B75erkVcGXp9LRF7FSwdcBwK0UJeQbK3zdn1e2bcnxyuSpYC105PO8nyfRhnZ/ppppdIu
Lv19WUMu2K7GBuDSrv/J1IURBjnGgrcTj4IwFBFWR9Q+gmZ//jPrZy0a4GnsBNB6z1Nv2wS7q6eM
3XeMB/LByj3Y5RdrePpKUp+yIvshGBJ/SVfbCyc+p8/fNinMTH+g5uZSNANFW/ZN4d6H3+LKt2uc
DwloCEYVt3bVwiOcXVVLAuTBuB1LFEsw9R3Q/I8yy4+pOXdYaMY5mUorOc73hpcNVpX9pmM4n9Id
5aA5lEPx8ewwfe2wAQ5LuYP7vTHKJD2KnyYyShBit6OIPx0uZ/uu+DoVhPCC1u0Esqq+yVo9Rwqy
Mys+cjNoZDQV8vmKX5eRP1LRTawlCqweiGyj3WuLjiCIs0rtpTpNO2t2M3FCV2+1zK6WkrsA4a5V
RjRBuiartljn+UiWCntZMi/U6zCfR2X1aXUaFiRbhRUcILUpLPXIALpNDhrBAsE3ILp55HWMnBoX
B+eetC6GdYFSnHNSFrixVblqoSZBWwgqc7qguD3vadG5jwRox2HysF2EY8DWaHcf9hZ4qQ9pRUaW
kZCI/MZ338WQKM6FPZ87QLVNVztzkPMN4qB+NUcjvonsMY5qWAkwee2aGLcrzjREPzpL6pKGHh+6
UmH1u/cSiuO+Jiyl7BxSBqBJWaazOa8E89bO8IJ9I81zXWJDNfbVt6Hv/OKiZ5QwPucxibg6npUQ
/aX/Ga70L00iwF54dflcFQW5P8auL1ZO0QiCBwzf3Gt3IC85a1DuN8Xh+YoAcJCxmUIvlnX2zD5f
6g5aazow0e8D2IPwPuOVuVZl4yZ0XzB0AWL5muotiIYm70YZOTaS7b/oEgqxQx8x060B6aGdT4j6
Ozwbb6FH4bd+h3ifl1V1J1Zmpe2xKLPf2Jx5Xihc8hoIB31/gfpeVqU23qthN53O/zZoCB5Q9U+D
zIMp7TDBXnN61sVgu35t1M5SCDTjrLO5om5FOZXTlXSajv3C9sH6k10GsVxfCGRGOnowdOlC4iLc
Zzq36GVciyMkWwyWV3Mu5ikiHGZpOZ/obw3hhTdLpPAcqL9/45NzZZEikQUMdcphsSsPO3nwGxma
26w7wRcEI6X/fVMG8ltt+XCyDDnvwyWlxyhDxFvER2hiAx7fBN8WKmnHTG6ulM1YEzq7Hah1RQhy
0MqojfNkmBBR+Lp9UraifGWb55luGse2oVQnouiYpZfZedJihQuQ6TjCSFnVf1dWus3PJadfTISW
2M0Ikib6QIUqfEjZAE9eKQFItc4rK0fEpie8YZJ1Mz1e1x/Tn27w5l2ges3BkiWtSRKSKZ8w+3I5
uT3+lC3MS2o78hi5kSsFLt8n9aEc+3Oi5SOpY9ZXcsu3iK8Rc004J8RWW8i1AIAtUM9pMcj7Xgni
Pm/LWChnp9UIrt+jK9fh/Nv6KHGG4AfIttktpdZw9kf4+EIVp+rh3DyggjSu5TlChJ5qbneDG274
7MYTCa98lm/l8xwtihNwIPr6L5jd7OpcTIO7ka2S0q++Dhv5am3EuJ15JwtMURaCxHM7Ad0zEFI/
/Q3UzGXMeAprHtZdnZqMFdUH+Ls97GGgDnsI0YCLkTWGkuNufj1BwpvecWL7/zQw0bXDGZaYbaoR
eNbO1VXch4ihNeIFvtSsgVg3MexXE//OSvocxp88s/+FTqDRtXlp+l8jfTVoq7ddwN2yHan+vDHz
GFFBtbNQoFmUTl0jbCxHjCG3sWid2y/AioK0CCU6V31zGyZ36tOaRmgfrt0dSnKUmpv4v4gMzntL
mULLgBqhEmSYXejTJ9QYWn6i8/QrOQ4jInVC+EKuZCrj0dOeVPNbX/Kbv/pp9EEyJ/pF1Wn5ZdGA
au/HW46/oIXPA6dBl3ck6Ejw5HG9y6DtOTEmxDlAHoER7+ZoVG8IEKwVQcxeYtqSI3C+reTHi1Fy
sM4YU9pBILBrZuZtDhyxtPtcn9ujVaKhhK9pbM/P50f22Q6pQUhhx9IlAgZGwHPrZUYcdwu8oGon
91muk4RzRF0dLcP3HnBXaevHg7w83QwABNUWxOGfNOQrQC5E1ukst/yc4BaZ09G8DJ7DTisLFOQG
XgBxRfpGsh7zSn0KNbzq3oQVusBi2NwNNfOiIlgwm14ozY23kS+RWd8v642ePsoqzVpXHqVvYwKP
S3mfDNaVuWEQW3E3U8bxf74nv2rjBuFo0GRYTBNUhNgyJjkHgrMaBi+QLAkvqlwixam5Dt5wyxgg
KzkitukZcKEIyFbsE6WRoVbw28qtc5iCUybgDnUn8cyCeJFhw4BAsmdAId4mSx4A5Cfua3ucOJp5
LH1tnKzQke5PtYkls+rAF974wj8OgbRzreeAc4jGpNRHxWEdLijgaadeC2NUEAtEUp7F/B42p9Xf
MiRLlRW9YHfgHqcLf02tS0AxXGKbrslCY/jcwbvwAjlpLCzFLRP959xHl5XVYqcP/LJubbZUvV1Y
TXBnBceeWWHkliZ0Pb7Z9ASjD4Vja6Yy9fea+ZghyXAaKDVxf2q3EYq9iXm2u4yPoKS9qwJo0FsH
sRthbAoiy/ej5Tj8MbZrxOCpAglxkIPjS0tzqhCV9BiVK+353Mi48alIMeZrmHaOBX4nPYSAGqGb
7lS/NF/4SNg4iGtnpBTmqvkrivj+5OT0j/13HQyCsjDDHqCs24Kj2pxRt1Po4OdlJ2441mGnnlOO
ZTWAIKV/80Sg8iewqUgDSxpu7iFe0Keu3Xa9SJYJ8UFWn8VpiJIN+DkotDucWDg5GJv4cu5daQ+Y
LDOSe2qImL/oqf6nfHexeJ4Drsaqyc/92owBT17iutwTHKZBGXcjJpv1HPdo+fPoVt4MGOpZfHkY
kZSnVrM1mHKOAqoeWRu7A9F4nH6JZdZ3sMqtahfkGLwwJ7X9iyAKB19HhobTRDea6+kxJbjyhBh/
D6u4GSgkXTkLq3u4fHHM0V88b1RacA6SrwriJa/Mt1M+KWysLB/NcSkYxsW0+3/ZHRnphsCPB1bo
gmzTZBUQN3+ucpfGg8JxhlAhaj5/efxVsb6iHzInzUvMoq3GDfYIJE8WlRPvj5RhYpzOfHM3j48W
AdFqeWIxx9eOYvbY2ABtYr2zTT2xwUY1FjGaM6jFz8NsJY+MhZHPULiurO/7CbPD4D7U6kTyhCeU
ROPKZWrI/JF3oOTmDdr2gug37z5bFzfHgGPK6Td2cTdTXZCh/U3bKTLXHzSebwXnouParQj1+ghO
Ot+eokQb2Sob0JPwHyBGyTdokMG1UvupCivld03fbnJKa+avA67us61JTunjBFpQBhTmrVKObXLW
5isMDtRZH455yah/uVheyqAl+/KGQeTN3VIDQ1k6dXDiANINkQhnv4MqgeCUjXOutlgfjLF8J5+U
fTuA7S0Uhc2Z9hmchXrY97/FdoBtTGynOtkFRj0uVbbVLCZC9bjZJ+7jTPC68/QciW5tNkx3gBHf
GtQ8BVRN6OOCoZ/RuDB+9AzBeu9IiRtXHszLUxCNrcBi7IBBGh54EjlunF71FDwRLUFw24dXR9lT
E0cL/3Nw59ev3RR1meclf0jScJlOT8HHxOiQseLBtWV2c/fNeEt9xET7MwxRm9Y4QcSMTHdv8QBw
WLZUXIdfSmvuxRyX5LpIHWwJZ4xOBtvmzzvlzsJgcr4BJo27WdK++LrZozx+wCAQg3GRG3HYpoP2
P5tUqcl5v3/0kFxU0f6VFz0VtY8sL3PRQktM1mvis0pyQOpeWe8BFDf3mU8xqHjEn450cRLh51h4
0ke5IuqHsdgZiRMSLE+2bD6ay1L4PQRqbFkw55Yj/msrTfQ+Yv2ivVBD5GKRET9RVsWDS0XtFpkf
5zoOSXIykGyxxeTlZwHfLYcM9KHFOIQ3v6+Efn6HLJ8zvPHoy0/b/LjqsrMhKV6kHKuLjUFMplFB
ehd0qTC56+8kL3XpaQ6PGI0v3aIEu1/YfaI9ap24vB52h/tEfXMB8hyMn1QnrXd8xyggD56kzUdl
BjM8Tnq3jGzVR2kPSbGeipNkDgnd+orrXnUlrNAQuu1VQMFoC9rcEf3te3rGOS44uZzH9Xu+//4q
iQ72SieJveJ3QY9AT3RKo7xYHecinmFMoCp4QovkaxH0VvWwkb7Qb+4tCCZ2bqmwO0p/u+SXZTBG
P+9K+k3gYBqXalVqSW19tMyQpzZwQWsRAXaSSbCzhCuN5pRn5ZqyaiSyV2EtrMd/Eng1st/qsU2J
Ftl7fuFWb4UzK5SIFg9oUIDbYf6PdmCiipFRehNd56uAhiDm/13Ywe4IRDLOz5INKaujl4cQcXLr
XiApMR6aE59J0p/9hozFxh8BAe/MNBmev8vCQt4dFUm1DEWW5UdOYRsCelJvPQE7N3+3e31ECR/1
hCd/yKq/KiLFyHld32FWOlVE0ITUJRc9kH+E+QvUsq2iwEl6vJ2NSHXqSJdeVepgsgon2QFt8Q31
ba14s5jIGQ502lw3bqtxBKvsfZzM0/6WYIh2RacsVrXAyAiFSnQR6qJLPZBhCysgFL2kMxBpOSrH
IPMTqiO72FfCdtoJLAbBjfbwKg+mWQHY65nMpCaK2H4kxXyiDpdnNP4AF4DEWm5iAZeOio0DtSto
J6HcvTWDfTTQW0IxCi3F4Vb0Z3hCjMYg3TKs6QAqua4oxGTaPaqSfW8vQDK40YsqbF0blulAJYzZ
kAjI6Wf2iAviwB0svtJ2/WgzBqDkDf9olXoQtSc2sO6pjAlJqfvWST/4LZxxyUCtIguvHFxs3wCT
K0XelqWtbHwJHTnoByFS/Sy03LRiEBcnGlszkffxFdrp9DF6oko/XQ6J5FeQjA82lCglzSFbTrLU
BvASQoIpdJU2VJDpQGrbOpw/ujrO9YpWNfJHk4vK47AB+0Z8XcAMD8EqrFu2tDV5KyV1do3BD2hE
D9VDSNy9zJjN+T9sVQ65KmLGsYYujnETUIbS6eTl3gzpfhqfJP0b8OBiBr4VMx8xcQYblNHXjzI6
gGMFBkNjenYm5QEVFNAKQs+PXu+4l536qW9qEso4iVN3/GxRYb1NinLJap057e4FHg45P3pWegrK
Ej8nUD6rWN2HTDCMKCel+TExrUV+UnJTx6DAJBtqA/pV069/rJHz4lWP8o1TC00LB34n/x+FkQLZ
QYJqyllho6/VisOICCBJ6Q3QqcCeF69pbbQpqU0G79ThkfQ52HNjtiGujvVVlhHgeftC4Dnc8w0c
+LhaCiKarip/zyzKAuITVkT+OgNb4UvbCIfJsmuj+Dk4AVB5rNTFOXIbZOV6b1hT2w8YqMRQCCsr
yQi5EoV/E+FJCoMw/O2cI9tFOrKPDa2IKn94+qnLpxVnkIFjmeWN14jCxPsBzOMfxFM96W9k6NOd
blyTpFqyvQlhkcrAw9bun1AmCY+ufQtLxVBfsHoKLUI3LUVOBve+9H5KMbwM3ldG6dTcaRypKsi0
uWS7+PeiNo0xBQtmPmWplOn+sl4CR77K/x+UKk0X2OgHqEvimDai2/CGZ6+TrnbxbEpXfrnQve3z
eYZcTdvHt6b22qCdEQwOfTOs7HGuSwPS/4Vc2y3fwXDkkSPF3idGTy89f3mpSBMtdRjIKf1vhh1f
hQwMCqk5+D9BiDPFHwNAuhrBUbFH3MU6qid7zRbWntUvOgjOTE8wIbk5BaEf+YxuSzuydp0ays6e
BXO0LWONZ52Sn6in02lkAxz5slZEUk8oY//Yt1MkYAS6tS29RLTPLckpQBUGLvHOeXcSPo+D2Tqn
Bw9nU49NPRtURaEu4PxbpK2RqKh5iWnBuBvlqQ1biWyAwjtXHimaiE1Ij9jQOnELxkb8w/iYqIua
MGFsX0NKp5PiC4m6yS4zQBj4Ku80vxNKEJT0seTdJtrBJHPWNKZuC3UK2w4mJAiiskGyOXYiNowd
aeXpCO7iW1Lw8YGo7p7oo1arEhWLKLcJnCe471xAlQFlQmjcXhu6F6s60+sfGGYBaKgQT6zLHAr0
2ZaYgpnmzVV0TNeIbas+cZU/rf/SDGIhfJf9+y2foDxifpdWrlqdcyeXRoZl2eFhulIN5vxk5fQB
Knk/j5LuvEAV23oL3uZktleZVDsTfvULucgA1B5zJa2/7TTss3NwjR5v7v4llmZNwerZtIHwSZ/2
3TO8BiPfrGe3Xd67XwF8aUXHoxLRaIdtiB+asvKbKz/84jexe1JJcPoAu0EI1BZTXGBYho0rzHCT
8Fy9YGKe/wgdzbDMyD1pKXrN7PjBjO7XGrBfV49KTZwthcsKyzbPF3wQ2SVOm6B1lgxJDKO+zCps
7TVddRCzYVtbwJbGaj/HP9I2y5xAIb5VQvHzmnTuGDVJm6+M1x1nDgcvq3ZuTekHPxIn0o7BQmQV
Gw92eSzXxRqD8m6xhp+jgf7jN8/12KJ5C+yNgCYiv/FNQz98X/U9RZgsBK4JMDDqHAiCXP1u4JT9
Ga6WwmS5fTZ+Ffas+8lUKv55sc1eRLqhbK/VN0g2U/nI7igALAg2lToNqfk3ns0QLXcSfin9HJkP
RViI7kchkaiiQoV3m17zYlZx+iEcySeBU8xPdj83yOcvtk1vhC6Nmz0iP1lXz7aOfs0Q9kocQvj+
FDArBnhotdYKvQnhzLyrd48y3TDQaatGYxh5tyRvNa3tlNvWvcKyyb3oTNQTgAw5IJO2FjXxvYDs
z/D0xYGnzeXtSMhYjT9JYcWXnyj0lXgEr8CpsZ1dnFdaFbcNwK9Xqp2rCN9QxIHW+laWetUfPh5J
j3BMkbaL6+gIHSNeXt1znSj910+rO4Nx7iKnMor/nsRUp7bGM4zBJCJN7OqSQghyhGNla2j203nA
lWT2PfE7yA6OCrpzF0OV73sOxs7Qex7pBQzEnI1QKk6qoVsRv2HRthaNARzZzA3CvAR0Idv7mR6d
0Ft+jnmDLatC6UGjFxLEQT1z7sIV8SObe9UU7GDRa4+jnkQwGHCstKEkisQtmLsxhL/IhOejULfm
g5DxAZzggISYc0I1bMsPFYBdZCd+4Vqd6JQhf8JMTrXkresVUHffPslvmPdk3EBbScTWQEv5dKi8
woAPKm+LER5A7a+5L16mI67tUgK/iAswkxNc5QAqlmMTGj6q5x87f5bw3whUV8SZlbPi0NM8kyVQ
U0U80E/mhPUBMGARMpQAZcCd+Jm/GpfcOKnc/I9LVUWFz6R/d9rx0FT81nX6ZqC4AnPepRUlTD9C
U1Dkk+P8uqM997jUSBFmo80CEy7gulOwGehl/ZfGzVdG0vkMcOnC80BW+FRK66aVflnPrJ6UfsJh
pr1mHLuHE3yDnNg/o0dczTfM7H9ZzzNrAuggRay9Da4DToQy4WDjrWIp6Nvl9Br07pDGfPsuJd7q
Qa8aMWqyeWmpXihtNIPFtx31JfmW9kw9cVLEEKrb1SyQVyG2waf6vrE2nV5lZ/6y9Z23vpwrxYXP
Ptp/FCfA6a21PcAV48G1u301syeEhQlur/KReU7kIyEzxg1vyaB4d9CBlxFS2zuJ6LdGhjTlzl1y
K8OKhaurLDz4jMHDsnRiQgmPKMimWfewVjdYj2reikLRVNaY/WlGJcgAiJoOApg77NAgw1phJad9
xHHasCF6+2egZ7QNtX+TF1JXBbixG6jYdNE2tLuVU+PXsTU/FkpqppFkTmILkawgIerVZ6+JVtUL
9MvbRZzLek0KM7O6wWYxkL/dXX5mQSdNY3FQpKp8Y7gpHAjMIndYzokz9rnC4lLxFAM9itNtWY/r
3N9KMCwFfiZ/VMRCMzlUIdzCScRgpzUsif2oVeH4ZL+icBuSOZDfogPaep8WQ2FQqsgEDIc4ZSjN
PK77u7ornPJ+moshR//+Oi7PsAdeuMvFbwiZfRP0cGRC78W1QHsJoSHoZRa9fFLYT1UNF6OujjpZ
dS8Pk7tn9x2vjBbOE5bFqnu1gmcbTBJKpg/VcaeJ+0rSr11zNMTI819YEMyS/D8ydbnImCnsxJ9Q
PzUrufD+JOkVUWsUZkwiqBMdla6j8Ue0I1bz1TbDDUa93+Anc6IOFwhvK2ik1qIPZTT5hgMkhqwS
ypoJ+RU3wI8csZLbYNRJLTMJN6IavvRnVzAopQaREyIA/Amu/xvCOlb1Edo+TweKA9LHcb/Zo+iY
I3nVgC3J3TJUk+tdRUKRxyYylV+qyXxFFEyCugBnF6ZT7t2x8UBkvurEJuLi2+Qx2c+nRxmSuM8s
RFOrBxqrdN5EKGA8CGPRfLnJvVrSbILThBEIAUbpCXRQ0s65i4Vg0jwiga5DIaJvGXcYMACAkEHe
XKHWgfCgFmrv7vhN/v7zlU0lD+Fs1/ju6jn3ZU949xnaW5PddpNwoZVFVdublvHDelwDmSVMA1UI
HpGl5GUFrlRuRfBByNJ3Ny0ML06zW3A/BzhSV3PKDH6GqWYw9QQhVos0RaKbeJVBkDGK+oL3ug/V
1+r3jn8no6qN+rgaPPk/AB4Znx5ZQYhMNN7tQGdqaxrdg4ZIQkAZl+ervm9YwrLf2tuywzWSaC8i
Q15stGmOZHKo5ppj4gsXJvaDAGatbsqeDUqxa0mu6EJ85k1YCnvDqUNiyz4LxPDBoto4eQ7juqG/
3nyL706zECSNvCx8wARQDp/XrIptAzjM5pbrTuBixz2TqNVZ19YSxSD4a+XRd7cJ7buaawKvqgJ+
napwE0Ugj8DOQnr1zRlK/E6ofM3uCBslbHmokji9F3Yh4hjFh9mTEbr59EeqXpqqJowHisB2ikUR
hCXAhtqnYjZy3O9OPN+uAYHiGl1kX5QkEyxvov8TEsCoyTdk4qbrysyvnns6mTlM6y15W3wuVLmf
mBUf5/WWq1Q9Gkzp3BuEN714E42n+SDkZ70me0tAq13pFHS+m1wTjcx/5TzriUZnGrngJQ0b/ZEK
Uu7DL4OHkY5Rpg6A7vQxMeDqOFM6F0sgt/733DsBhzPWL51oKky1FwRgG2eUZbgPGE61ZbdET49O
Um/Mg/fi1pihahCacthkc4/n7iwpofMa08QMa6A8iEmT9NPh9qbyVGW6xOxGFI57/mVimwZjL9G0
M/xRrHhd/yEPQ1loUX3PXWdbVNZ7MyIKVjkOfdHakaaGf89YWG9Oq0ficMHrRi6lSW69ao5wmdex
PqrzJ5Yoki5d7kkOyuDQ9+RVwSH6uyfpKKZijGqWEX9/pM++zjg+1tMh0BggGQYTXUB0bPA6SNCf
R88cEF3CRtZnsGDXLa6Danhi4MQcBf5xH47zd+CYn4fyhPwd13ZMrzqSoNIXV9zwiGEdtgTZKYin
gbRSb6O8WL/RlnyuGrTpSYEFerEiitigp/TdsgNEKBwgZmDcv0GVP0or6c3Jl1x3QIVUH9AfX5/0
aeg1P02ZTKjBKMWFN5altVxlciaRW7SJIslsTdhY60rAjw7bvG4EanjrtheuQ4KL7a4JJRGfa3Ig
CJIxf6UN0Fqa3PojCycPWKF8JgMR2TwLAbki9WQvUCXQFMXKxm91WyvAOFx7w37QhVYJ0XOW/y5w
Kj15iTvyMaH4j/So47XthF45Dr3vzw5qBkz4bmg2TPBhAigi0qnjsbbxE+tX/cBqniK2iYEW73/H
N2PPt9sL7up4R8umcW1d+FVUY/qMECItpowYfP+4PLq4YrX64X+Q3xYYZ7V/cH+KMhmZQU6xh0oR
Rei/Hx7+3YQUkCTAqxNtjpit6sc652i6vsYP6tvgnBIZhrkpifdUEUwM2e7QQVN4ho3doQwFdPMH
WuaZwNE/mT707ttOEbP7mMZV1Z6qJAMxaAGNW8ZMjDbdHT3hjdgT50Y2ltduT857wruQPEOFFdHo
ErzWd8EVpsQuwDte7qMAvrgDvEjjGqyfcP7wilUZLsh7aRXtkzoxPuNw4UURVopTlFpNckyJfadG
UhbwuB5FtsF2+SBTlzRwnfz2sdzgsQkTAlWSkAZoOgSobedZYLJzd9EtqBZAs7jG0Haz4iEUT+9A
QD4SPSEtBQ8Wk6CWsTIG1hLizNhVFVbCFb+NyA0d713V5DlOzTOHSn2ssn7E2/N0c/EwUrwx89zi
eR8avrfTj2ZMFF5+Iap1JEvSPIm5e/k8CeHWOgekgTGxxT/Va7Hc1z/EJ4vB0IQLERmYNDj5A0vu
a84evFW3RSCSUqhbCRvKUwvadDNfskjh0Cekmbo+DtQoRCa9m1hN7snFXg6Oi5RIkKd2miKh9IPJ
W/ub2ULgCrpD9feqi3uNyHryAhxigFM13WiEiSS8yvGt6+2L20hKsQcj91SMz4oMwEUsR8HUrLyy
NcoKYxGHHSFgqn+fSFI9a/eFV17qg6kTYRLgux0pVqEmMJJWSIn+aryjP73j1ty/j+Af8JUj4ESr
kP88qIIg4eZnCXuYPKGPHvuFNurvGrVqiOcQJSCdQkklleV8GxOsxnJxsiiSr+7JmoMTxGG9X3Iu
BYzT6hMwOLaG0vT2QRQKGU5GcmacMSJEny+46D1xMBgp24rMssk5Pu5si1inTWMbyJ23Vudb0E0N
DY8NTS+mruV9RLUkjP+PltQGBhWc3veYcTv39926v2suihr2IK/L6V8RHO3sejL2dZDgTOP8LKLP
//dWzHlUd6eqWLsUZcKzPSQnkh2zXg9UHD08HTnPbBNHmOdwBi/GlEV2Jou980NJWQ4vdbdn8aPO
jCWv9OQ10pRXdApU+jU4Ya7J/ugM+QcHmiITd8qG9bf9Z4O/U09EwXoyt6N/Ohyi0ZBtG6qujV2B
YIEzqCrQVxTaA8lExrK4K1mddG79qVSnkRW0pzjTWAkBAZzvM2C/BqnBNg8XB0S1f42JeShu2wuL
ULjDCoJ88yAhEPOTYoyXvgzmuEYCMkjWQ1dGjj9/qICDJaBRDVc5OzCcOQRPiX1y792WqyNMcDIU
ZY/4JMPniZb+8YLwHn3wiwEj97SjvWGUPxFDlGbmf7CLtg0ijcgDInvGyvlZYK/GMo1xRHWvGSeq
dydNOhSPIn9c14tJDCAGQtbbm4EE9fpMPVvlnfYscA9mOetlnphdbhyltaYOtG0M4aHMn2RLUXm5
+sOUFPuCmVn9Nu+fW88HQP1PAsxcERYAHueXflc+wDROenTatYZGGMXomxMoamHW8YnIoF45C7hj
PkpITj3yj/paTbByHQbA0zv2yQcwaVc7MW1Cn1yn5VVkLxeq4FklTTu8TG2/CEkQDo0UnoVvQJqa
dDlQQctN7oiLuH1fgILu3EhSGPo19DfhG99ygAhHjINFdESKLJhO1hsUuiO1d10EiYz+1CiERUPZ
B5YbZ0KfnEK4m4T2Cb0ogSTSSr4amcLAURqaq7oND/VoNAT1V3lZ/nwAhM02AuUnGiMJAXjAaDyU
uOZ9VQ9/GdnRS6y9xXKcFC/TnGtUkXtHZjHOCjNebj9b76qo2vBJ03b72H3deeqDsInTX39Adp05
VVg84jmUqxmxKs1xPwfqJE/JbmzcTEHlb/jHNJsunLLXRa5Jl6IzdTUW6SAOZairmvkhhD0CFKSQ
NpwkWHeHvaxzp1BLpk9vNrRId/d0ZJqrUJcAliV4CHgZ+uIt5I8ZklCRS7KBt2sN6Gtb896sx9q9
UPCSAeVWTaXaZm+exxHK9VDPiqe7n9GvxAfrlP6sev08UE94EkK2Yx28J4hdq3qSX2MS3uPo6lGV
Fp1qR5erEihejP/HQVDeofrPlpNI/rZzrEazQqiM1VKxdUh7grOnQS3on3yb7/UdtjXS0HFfDXcT
DKlrve6LmLTZNSfPpY6+MioCmzeMFMY6ygXUfR3PB5bUeDk0IT9dPRJe/Tv525s5PCfIct367/Uj
BcCkDqgUNksoyrU6/az01TaiNkZKFS8aGEE4XO/N6yXDTmrWVy2pDoaZGKHhU7rWnOuHjW27k2VA
/Ylgsk77BfKkQ/mZqHQSABztwybAnlk0XXSWdyQMMY6r2uvEGN95122gtQhuI9QoURvaJtnr4OnQ
aPzHdO3QWav+WObvdcYkQE2Cr9MCoZgKDpaqibsASvxz1fl7cdJp/x4ydp9OBMqcSeGYjx+aCZ2V
/wYWOD6VH6/LwGCK5/1Lu6NlBf4nSvUiFnAOd6+G4cApMrJBrLDWPBf0ZgUepDfVLFjzOIolNWyi
skrKgd4tMG4sB0hywDIJMJWFGVGRQxNrpd230cQJg8YlFskfdEmSLGI7kRmNYoZoQ4ot1RkqI8Bv
fLjmBvhnY8051NzpT5mijEPsHP2C13QOkNlz4/oPedCPPIhonnaXjl5KT4ba6J06CQus4C5OqhdU
L2+KTwRM6fPk1l7f6fcVq49XcVsCNuU32pnaIoOUToYw1woN/AhSTj/mnFeb5U6hLysOeY+AsB9v
QfXc6IkoU6Jdx7bSnuTI28WD6fjGxchsrE1wI6JN0Yi4D+z7cdwV8KcKe/YydA5hv3i/EF7wkRSG
uVcnIFIKukz+zUpcEVnRAfWyqbnUdRuhgvgofd4Qrt28FBgVYtMwLAg7HoI8QJSdh97b2UFr3phI
dxPUnHRJ/5xMH0Vj2P67zkhEkO2uVaS7SRTAtB7AdbCIgOb1I5+ut5Kkq7nBeEIMrFwHChPCCK48
FuUiKzki5D2H75MNpyLzaAp6Wf0jc9zv3uQcoYo23Mh69vFzDGb5hxyFetsM7Ell1G8vaSFswjqq
n52OGMk/6IsSeYY0AP1ahcfcTtdgCWYj697t+xOP4siCObY4ZC9UeeheUArz+/xOnfrlvWAEfST7
u1Uqc1IpXn5RCD9kmSGplqND11Y3ZavDZlyDXRKJ7tHUbzUJr4wyziI/KDrHkqvzYhGRbzfM/6iu
XEAtueensx+onlzo9ZeoHN9C12TPxPZlFXxYxyIfSKp9o90Zl2JQUPv4mYe8G5E8ZZXXb4hg2ZSO
Cgaa9pPMLx90snlb+lu5AzoRfoT2FO4e0MrGR3QP/1Mx9A9JxhOoqRffmMa8H73OJgyae3xNAIWW
6D2a8TXqgT0AluaB68n5nXl4qicYMQvlVgzxVmftqdKXw1WhURoc9de0HSwgD6yGRRpj6IW9F7t8
muTrn7sLX6HhVK7JjavSGm/Lre3gVrQ5reIcIUiz5f+pp6bZd3SJPyRWJqrxFFNDbSbkLE8sEjTx
8Je0i5o0r94kdkrxvkHHYbYmb0C/WvdLWIQ71vkQGWzo1QM1cPSRe3L98/eflOI7/JnBGDlvCoco
AoxyF4wVtcOsWo0CHfBKfO2Y8L1eOUEukcPMjtmzbJ366lyFUl7mBeScb//gxpvin92kuNneaXED
dr20pb7G8Job3tHE8/0NtUBtp9sGhEecizjsIG9wVYKvRo7y5x7g6K242AVMK9ia2Jyb5qbsAwCo
c5/iFtmRKLwiDtUOQCz3z46VjXgPc5bexNex2SW0n4MDXVMwMKv1BKUXH1Yu+mnCCoU5yISd54TC
8gT7R/0VQtRPhegUeZ0QjNxynXkyrk9Isk8aDfzgzd+IaLppZEItDGSaGWFVrpbjB5peoYmzuzW/
2jEBSGW7mAbSS/gwBv5IblmWWZshSDClREAmaPlng1eZ/+AeRzHCsoa3VO0wKrQ72Il8Y0XXN+02
yREJ7NusS5efS7bxPHUTZlTgq6zAwS2N+AUudWdA0SwMVqQ1B7QPvf3V+Dz55sOixm/PXqZn9aAK
VBlb1IreB9wc+KuvYlFduSi1yPeQF7MLLeZOd3D3My5F4k75vfn7EHQp35SLVldHNTxGj1jFv8hX
buKTQTXBfiggtazK6Y5NdnvS2oiGNfMTTEJgDfEunfzMxhitf8LtOS3Jx5nReakPV1fpM971+kUw
tA+8qdmQxUSUZqbUGBWdJDTXG6HSEt1lNHkNa4oiAP+Ggs9/rZzj+9cvIhk7NeiWBvzQy3k6KBSl
XVT737vo/1Q58wSStcXj1QMACVl9bCXpdS+msP7pf8WkYQ7BSUtxmzIpXwpey7PwWt08vnOTiDJk
/1ck1mYDs5dyFfkz4368Nff9TZ+6lbPT96fqGl25Oz75cubsiKOuGYtKJZHTrRCkXK4IySYJvraA
R17dQ9I1KDdhprWWH5kox8kdVOAxlqoC6N6GQd+SlbAk6CUD5qIpAd9I5MI3qS+ISRohgkfqLUGN
OV4GA0Iz/jZrd0+VQMxkQs6IucyG5Nj38B5sAGnnnUIDyRvdPFLTFzXHeSxIUsbvAJTqhAonocq+
7A/JjjWxS2AHS76EVAEgJUfWieZVQC/c4+KYoeoYV4VzbUgFW3vpidZ7hXqPIWt3rn7Iu5jqrg7d
6SnWwOm+zwHjUruDLmfMdLMAEV4ZHfgb5YrGzKQBR/BJdPCNVwb/hTnHsrLsOiP3powTRwkuZY2h
BtVB2BePCpJ6eM/rh7I6jYYPT0WWagsdTIeI2pdQydqghxMbY9QKUpq8M6EOqnL95fCMRg6OgAQY
4rSZBEwY4koc/4isRrDc+XF9OFhpfrxZnK3UHqZbXXSfud1Z9jDAilpaFjDQPfKR7GKx76HwWSoA
/+1Cxg8kC9Wb/9ygJ5QD3WxS+HxSIh0vylLRTjTTRZPHJ+RHRwkDB/y7xxn87v/JUwlOUIJUrHHp
GZjSHIMl2EdfahEm+kJkJUf5zF97pJOtfEF6wFwaKJRxFjBrecLm8MuYj/u9ffgLMVn+3kNELFS8
6q6LkB2ALIQgH2ehw3ajzA3G3lnKUnJ0ndLvO5mNhY4e0Cg/0UTHQs9x/L9Tu1PtRQnPHluIqi5N
EfFMbVGHkBOa84OKrU1Fi0sZhTrDTZfIEZVNC60JU+UuqDTiCBW6bT0C/9Qyq946coJXymIyQvaK
LXnoQgGR69TJlZ1dv3GAndlKsWtJ1LiOgGZgZPEmPQiCdHMWUsX2MGqKhsZUWEuUFs9TRAnP28uF
mq8XLt7u+LBqUTBkmy6iMQfYbShbN0w6B0V7S6q//TkjzTnYbUuonaGuFkmjJqPcR7vmLGrIbcD9
Z3LI1SbS1Sg4C7n9hCRIZOPjUxNSu52SoX0IPGGbHAeiwNbui8rlGl6h4Ei/cuvKB7WbcSIJ2DCS
qIdHO+Qqe3Acd7i/NpsidIIYZsNDaL4lqQ1C32qALIgPXIu92PuXuv/8aHk/wkPKPiKQJaWffi2d
wOYuZk0sx339/+rlE/tH/qpNhE+GQGxSk6PVNnV0q1nMF5xVSG+6feY0YgAp7SGC9PHs7OVxzVYc
irk5XEr53gJJqfDLecC8vMyPIMlDu9pBAsTF78Ov9pEKV+74UAPjRWIAIrfHLIjthq4iEz6POHIl
eOkM+KyEIRM8UI+2W+wQS57keNblowYdEVqKD19kkXUtnzLUqO3m+GnXBcLeh9XIg73hDtH/reJZ
K5NVy18pQ8+RFnf3TEBLrDW7CUlzoR1y8jafbLujG5HlSbYLIz0+DBorY0a2Hca2hebdDv0tR070
O0t7QiwROl5qQrkR6eHdWAFEBPjZOMXnfa95jTyd3bCEG7X4S6iMOtKS/4oro61/QBJNToAJPrfP
/qIBcSnU9MHEc3mlAUtiJ77q6HSYndUg+XqN004qQqyxk2U/kgOY0PNcg+gW9nWoTIhEU2CRj2OH
4E/tKbJQgqe2DZlXFeCYZ7OsgKM+hLeKinGt57vzeyEX7rp+em6Yww4/yJuymBFDZUjmyq8GuutS
qwSasxrq3+t+fTJUrdVH96MihuJgvwF6+OtjGuYFyn/ADlflrFqcHJxUt8Gw6LqnGkcfkU6ffzeu
7XsHJG8/PAOYPRcQ23Zp27UsSIbNtsOGFPoxkHfyQtZdfn97b6FibNORYcZYn8NAj3S0OuMFBxwA
zJBdCMaVteaLBU1l3IKa3AaNqubQrJI8ikOK3MlWNeEv0txNgEExWZkWQXG8u/sW8j99yYPT5QYY
780U4oElXnnv46mSpq2HtoZ06bzQ09v6uGPfrag1kOOwaEgKrTy56IsSY4oa8IWRJqXC7X9bslAD
pv7oopY1IowmnnkmfLx9uZnwooUCwi27VvFsQGkDMCRfbi5jegu2uG39KfxoTVhk5g0BQz9eDqEY
+cXvCd1h7W0i9+/RrbqorZOxCnteTY3qD+UC99/DJGOAC/ltrXcjz2UK2muqomYqoCn3lrjmHTis
IGklHwQkpOVpCngs5iTToO7vl9s+3ruSr1yu/jhppLr7cOAMDF3tt4N+ibTnbxSAOvXRkgAs5+dx
p0vsBSySalpgQnbzpnARtfVXr3SZFwwS/ygf066sGTI9B4kxz0UR1SqSm/Drd037YufQ+NcWtAce
HgFJrAaVOePIoMs7oV/pbRVCLwRBu50nQlGb8vR+aQyXLMfv97sEFunplDN0LLoqO6S/j5+ff8WB
ngQ890uyMgwEUFby6LpP1n+vJb3w7PcaatdHXhmXBEGsR8A3Y7An13Z9TO7afFNw/WQfDkec3rC9
z0XZrfNP16moOaAtOzD+VK4+1EF2CNS8wEoYwkipDmacpGYXsB2eFRJlTewO3I9V+lRCz/313Z85
ZCb0HahB3DuQThReRkkJRxiPLCvLwP3O0syxUPl93gGSnGAXbWs3DPglh2iGBiVlWCX3iMQNPuST
P+3dPiO6LCnmr/254s4KmooKzNoienFC67RMIAjP2kda5GoRCuNAr0JJNdQsTlVbh6OduYarcpI+
4yo7QyuWNsPRVqvbxEr9lXgAD4ADPRWDOIjnagM9YxZHQktlq1nJUsJLxNfxlKBapWTlTNTTypNa
5/TpNj2SZXsIbrUEkaMoJPRzQ6DMK5tRWfLKNoqeQQdtdbKViKzUpwd0D1/BLi9HFJdizmYAH5Tp
f7NYqQSRVI34xIp07uk4iUUgxMyDWgizJ5RY6+0PDzVPpxlHZgaK+pAbzcwS3lYAy6/UEks8lUOs
C68zB5IrARGalP04eHyFxq47SwuFHubhuKJ55oZGPP71DoMWexhzOtjIBaJeaagbqb8CGJhWUc3t
iCQa8eI2xf8LLfKu+uQHRMi51GNEk7vCv0kuPVvXrXJTZF4tLsSAB/rWVZqCcQpZZ8hi007gVg3L
fVGPZiIIdp1F39DYzgif/R4SQKKhTZmnK7uLtkOCxfhw11mX9fyKSVR9bks0qk5nHyXQWcA37dg8
yA0BP+nvPi6KSDTPk9+k4L/v4xRweCbIqwdnv/E7JHzH4/QeXEp7w16lIvNfwxeVszjkRgZOSv5d
1ve7mdZwOiFDSMGFTGU2qnmnyzCaNR7ctwEkRl3MCsHzi8xA72GyxeJTGC3rsv6/4WbBVRiuMbiI
qMVyEdF5RedfsBKGhm6iLYrr1XvBPat8n9uW9+k+Evz0yaKyLR1yZEZkxrSc/YHgOHbMuek4AtzD
2+I2jFdgZMBLbVfCdalGikymcRzz4udjZuDFklw+3V9wxaYdy9ROUVlqzwPTB8Tz+CFtO7j9j5Bs
7CYAzUA50M6lre25jcja4rG0cL7HqDX7NKPpkp75VEgzu9giXzfuLNqI2Z/9RDgBmi4oDh7f8YAq
/zMX/roXgpC+uZuDK7SoHO2LD7N01qDpjN4AzObMRacc5FUkLL71tVcrCjur4hvNHVstNrB93LIc
aL0TXclHh2Ws9/hybEpam+boFNZooADMo1dyVXMKayAm8iZJQqOI6Um103jo1/Ha5fXXio0nxEmN
j7T8sXi1YsEhSuh3LGGsVsOZVHLmCuqS1gUjHC2wS2X22FmWxrEG5DSiKKhBFdT/YnP9MD8X8NA5
SDGaaPpWfOGuSokZNaf3eup1jN5L7f6yYNbLGGmZuvl5mvmVqcaFOsUpux8tgrP2jWAZcOkLjSdw
odweBN1GOQimtM8OkLcr0SZ/C9OUlrouHzQ6wUMIHdNR3bAHte2M1jRf6UHrwiaRfo3WiUQqenc8
V3w6A47XbGRuZCj8E0dDUE92K1DoWCk3AEDoxHyVT6Xe0bUuCatGZWavV9Y+VmdD+Q9+afoo0rb1
3q3JFg/iNdq96PVeaepDlke6kQ6PBH2g+L7jdjiKzvrvPUuAShySJoFmu+Zu7VNfpAmEIq2qyiXG
m8B68ef3p6K/VeBTDMFiQ4MyMvsy1TYV8tjwWuOnYkhRFEIEG++q/7StwxpuzOHvIpjG5rmHNL81
0muQ9sH3XY6XruMaWRe9LyTdAzcnMmzAWsUGs6A6xivccxUz67WdtLEiRZPudy9YxAGqrjgpqnQL
+Hoqje6hS7TDuDJ00MVmcvx8aRcYeQ1E4Dto6AGi9x6iyukPXBgRNoQS767ne50ZEwpF3ui/d7IN
ovofUy+Dq4omGi95rQNUQJ3EvoC0sAUo49rYOJvz/8Zv/yr9+7anVsaAjVltCFr9MiMln/WJLimZ
j4uCRIIVP5vKKqfppVFdsyPzY+iAL91ipL90XGP7i83jCtTYZ3A8WSsb+ZTnfNsqHOMoRJg2Ys18
6Sn1Ogpc9qpIFLrporRzqIQoou8JBdWwwh9rySCv2wSf5OSq0vV5zwGzMUdxdIJqc0IJ41RBsnlr
L+LCe4b3EPBSbF1mLlg1/lBl9+iZ4X9/+vsZSSj3RCsHumNbwJDaVSHgzXC4sZAChZ4ByLCuHfam
n6XDcQPf33OBIo1OJZXtMY6EP4I50C7KCiHisuC0XD1KmJovrjzOmZKzA7vNKGxTYdOVtkH5Om8w
kAHqSbzycW9p4LRGRRB+WrCj8L2bqOzUJIPp7OIs2O/Tgs/LNLWMWr+Su2OmYTbI9MC/XP8Y8cHX
JzN9iMBguC5aGxMEbkvFObSN3RJwSoZfh237m8QivtMGe0x5JY7xEsMB2IhCOKMtWK7/IE4udxfJ
Q23PJkj2urqdrFfzFyLyLrnMRSq9gNFPQNml4cjaYyiY4y9Zuc0Y3TgFZtWTPpMPHtJrejKU44Cb
IgjM6ziKbrA/0hYMxslunvLnZaD9HCv9LFChIGU3wlStX6NLvLA+5rr568yDqq/LhEeoPBJDg7vl
jerZ3Yvbn9QrZwCwyKvx7T9cZGcsMToSDrDzyKpo2hq8eADZlyYb1KSefcIvzwetLjCIQZeBUtNA
y79ztzLxCpN6yW3WWA5TH4LO//XiNjBuZTlwZtOiX//XoPBgbsHI4c46ol+n9pX/9Mbc/vQlcyid
sWtn6dnXjImFlQnpi8WR6SwLAFigiIg4eLdCI0uaqyzuRWmuXSWmGQunu4dNZaRycsvtgWHvEFs8
vtikWuImEaxNeabP5afFatbH4zX40hJ26dZUqCqwC47wSUlpI650HIz8L6bwhPuSpbWlUmV+HhVz
GI6Mgp5QvzuAKMFIhRM9WOb8LX77YitgsRDtpo1r3Nd5kMhrdc6jzCfDlneXXoDU4iF162zHidGK
YG/8nE6oNV2jKxvjLIZeWEfuziQF5xxOyzImw2b8Ki+mzuEEOWE8NMaUhaiXK+uAmbpAHP5EoHgR
+YSH7YRqvadq/ZRjBYBj8g/78xJhZw55W7dyEfxdpWd3bqBW/QObLbERsAJ5l+TS58D9cswOCX/K
TmQLgQXohcMVAPWMTVEdEO8rR8i5O0n1e7vmf1SLdJIGmc6ruXL/hnnRhz6xabxB7D1ETwMtd3AF
+2tD1ZiNVP/MQLDtLdd7HLY2Vteh2mxZl+KLc+0XwBQhyopgMaZa5YQ1kJoUotUss5u03mRR8SPv
3wf53t2qmx3IOHXB6t2jKaibXkf+FVfSxhOmfAROVXwmKSmEY9/htgiuSg5a7RvXQ0NvZHltV8Qp
o8iZ3I7R/HD3Tkm7OEb+2TZnzQ0I/ZNBuidQ4xjivNYy8H9PmFBF5Qt086tj/gJqOHcW9Pypijvs
L8X4sksukV5z6wuvLnO6hsmk/k8Rzk4tatvP9iCT2t643vH3DFp/JUTUKzhDJfDMA2Ud0BQFfpQM
VFO9eBkuHP1MG3V0Z4WaR31KOFC3+SvbdGBnmwFupNp95fyn6gWkN0PGaFXVngZI1NuctVzWa6LH
t/ZjeMMnv/NIsiQaoCKoA+QUTqrzfT5F/2sHu2gL5vhd2DnlgvcCrhVpMmedRWZiY8lqVBm5pX24
9z1eK/+qRLEayCQOyns9MZztGtrj7qUXBNWDhpKwMy0/hkPQ81qkTwEetdHEaQHKkkCs+Qkvggkd
afS10qo5PZVFBJanmT4hA91br4vGTyWHmsgeMxHQzlbTGYfxqDHkRnFkY3PVpx5AwavO8JbRtCa5
+Pss85Fp2T4ggfhbBctvOKbcFSPhF+Dr/5PC4AaV/GM0F/Ws4nLe+8z/z/EtYQHnr2xbxVoKoeKZ
kFgz2yQB5zX7turd5iGxgWdABpK9nzuJgTFhefPRORa8XKDZuL6dXygIiyO8CBZ8bSM87JFugdcH
Hi30ptQJRVYrthucGC7J2rDgC5G3j7ASEmQh5K9VXZDuxfxt1X8GO+s1xqV7FQ3h2zUnAA6RN2zz
CfZ8d2tH6GlAfWi3bjIRhPVUi9QhGRvkNW9uABEkF1HKHD0zXGBsnAt27huLrWOHWQElzBD894O3
1UG0PQUMnDxM5+cIJOZY0cnILx9t4saNY3p3vrQcItX+nqwLnjBNK7k5nfOV1PsiKiH6kA4zFWTh
h5SVplsvQ4fyZn9K7ixucbCXsnCcqNKzU7GBLypn8jho26JBq6Y/WRNiYiWm1KRAnKijiROnGYyO
76r5tmkUy7b9pcXr6PNSY0hrc1g+L/OcaD1MiPmD0MBn8IwT8slfJt3S/DViGWF64XQPs95fB39y
6Xt29hqUjWiziN115wDfxTrivkNKOeSaHpM88b3qeEfgilh4G9oZ7wAIZnhCAs+dxDpN47qdC8Zu
/aU35+mVd7amBRSPwljre19okjFxdACLy3Y5HY3bc74uWlIlAZZG8Lvj02FGRJKRfByrBqtgOxth
EjCJsWaoQ7aUBSL2lJMB2B9VUz6dcVqjNqarpT+LW4d5qvLzpWqIEuK60dkicMGsqCRk74+g+DmZ
G2ahcnKp5WgGGx2ft8sIvJBbj7yypUulOzgpGyrGpwpYMzStHuSJthM+fW/R60hbajoEgC3nzL/W
YDolYGzSusUJ6gp94cccDxcnIr8D9M0cah8FUuqGoJftYZqeistWNeMbTLPXECatSCUrKj7+noo6
er3wN3dlrfqikUKo2nCZqMyXlzJnwg6OnFZOs4JW1+7vxquj5pYgoPTKEQNa53vXPsGOveIhA7CP
tDt4K+H/ZlWIYK4wrDeV07tiKT7KGkBDGu0yw4Cke4efvBwoaB9cv/orGshKBZvPdFFs/ZePWYFq
9bKSrxDz5yw6RHOMM8XCcIP8glKeAyyS/FuLvbNHwqVDk7tM9VTR5Y82bVC3XbL4MKTMCQ7AG+oI
RjEWIopgPhpiowfeHjrZnUQ9UD82nW3zjPWsDneWaGFgh/y+twqepDvNkjSF7vsQ8vZZ7tZ3AlrT
bA79f5L4y61FYEtxbMlPTiK0kkifZYDEDwtErWEcKPAHjRrKUD7wyqj7XSbxNdz8xptZK3IkjcVe
RwF408S4nshwMQP1jX+Q4f8q6ZjF91UCGZOQ4bJpG0QQqAjn0r/YUWXvlLqFGlO5F3y/GakCijYT
ptDCDqtLOESg3Aa130j2PjpwEfYGTzOge5BbrMENS8vEw+loLEByDSlE6DF8EmbpO3jiB7tk7njI
4cQYskWz00UvCdItytC+Ux6vQMXOmsVJN9PhmmfexctxsCo0MH4CzTUIYZhZnq1YVM36ht3VNhcd
Ff0sSiPc07WWgnFjVh7CmqAsBbRukaKKlIDOcIF4tpxJTaasKrxISuonwJ4L0VikfVfU97eXrJf0
OlLdkmrPej5RwzdAQ+5zgAhOpPpV4c7gcysS4tjsgwBvEzy/g6hKzwXmaZCrsnm3/KPcAFixtxzh
6nHBiRd8R1a9W592fjRr9PCdygEWdXl3cWsfQ2KwsT0c1GRD6LPRASfSr9wgZPcqwIwCv6indqDN
9JBNJabDKGGSVLEjI1xMGSd1YkDFLgPNkOc6zS/TDAZPbUQIAS6IlcKkcVcj/HvE7i/BVGq76uZX
KoWSmtxnQiJ62FS+mmbKuEyDqU5e2NqB/QMZPjwUeqT25G/UUXgDIonWVITvRvRfoTj9Ov2rS6D2
0N3EWDhWR35lDW5Ed+jmtc2cmhdYQwu2sUc7nYgS+KN/dqZ0e8+w+g68nylkHoCTbB0lEo7aUcv+
0vZJEgnhQFAfZmljYt0X+UDHdrP4QYpZ0Xj9ggTNJ1dCD99mbgEHgQ+fXf6KcfnIeiLFaDwfL2t+
HmWSQuXjsKs3/+dhvKzTe/mENtQyj0xvMkHndKJGF2k55cJfLBLm5pH0Ea1FVt/aCmGiPP563kAH
+cnSyYcxfII9BjPtX59W8214v1GQXWQZSMQdLdtYi4GIqcJalsh00/2NzJgh6Z0xIB7j0Bo/t+Gd
mMC8OV8pSBuvY7BGm49sS+qy5yUyuC2osKoNbOtZfU49AByN/atEQNMB5KVqoEbI9l1JsTCyRzKB
lTMikA8qfwXSyJAcAFTaOjK/4fUChn6bxidElshv4DCOR7NEAUIMNkxumozZUgJDGQtOZuqGxalz
+kTImGm+M2AouxXblUcXhyjQPxWPKldzvd3JQKIdyG0UgjS+EkXQ0YbFLoDSUfI2EKXPORFSA1qX
N/hXytN4jB4fz9wKgnunUE9Z37bjOnjnTZBtr6cznGgzXVc6Apn9R9wG9U0H/nQ1M3+EwBeSNQM3
Y276TAClI8zrWsmsk50ZU7BB5gNTgtUBrNfJq5EsUcztwqnnivNIXpf0eeh1Dz3oYpxAXj8cfIxF
PFFilWgCzku8h0lPSclqmLcg1sz2u2UtVemwT1nlb9/2uJRQwHWfsuXUCEdnP3X3tpCLZhqO3TTZ
u4v+RKjaioMZ+Ti1CQ6ZN2N2FhPft8tfkayVy7NqLq0mHxAmAHm70am/z1ic2i/FevgXDRzE62OZ
SnZUpKDC0rbGYTPrBsQrmuW9Z0ckaj6rRPBjJRTjs2b2kiQSBLeeYaNd6Wa1idfmchGD+90zByXk
U3C6r4NTNmG8X5W5tt6dAefK8xaACrkJA1R8Q5z4rScqSB9uATcMO0lVd4LaTUFrZaivWCsO4hkG
L0xxmDhc+Pf+4mUhUwtZv/18SArl6G2htVaY7BOjd9zry8cWAtKmvXu0kVz3eVCqZ+aYv3gGQY01
J3VsyDc/6CNkcG5isKvMVDzz+x2EW4aZ3gAbtErAlzoT7dcafPdzXeGqo70q9I6GWCDA1qpPscRJ
1rlChoFOQhxvW2JSDjpw2tBPp5o/FvsdKQC9sx9YUhDv0SJDmpcLMsxcihqpgY3Nj6I7+fq0GYkn
aNqiUOUSUcIbrGn6aWIB1VxLm3F6ZgEOpkglsVObGDmQlb7g+P5ldKAHltsoM/3dbDceUQ6QN1QD
+o4p+Tu/m6l393etMm01N9HMeM9cRtNtL5K9JHzbq02BozmkFhenytFupLOBUqnahPKwsPTaOX+M
HinHlVR6f5IuGx4Yo7fDnIJOqR8q0uK48uzCiyNWff1nbUlMuzFF537qqKPfNQ62k29KLUUGmAxo
UsrhBuIuHMqd1Uxq6ea4+MNb5UK8DcKq784uPYK6AfTWC9N9DgLionO3qTyJeNb7sR42huUrfBtU
RZTsjXo1STdLiODwWHhPo9L55T7/IDwAlEFx5IxmP6xn+p9Qsq5guavP0eBH4P3OF5uxUWlwtWmn
pnUopjcdnFusN5eXMaupsChNi2izVzym12VcQrIT8hzVajMwuZeJmdtBFKO7ozW4YVhNUqYzLZiz
Yn8e6YMPaegQf+9y/wTYGFOM7d9RrSh09ZKAmT6NPf2fv4LZhLyzq7RNYzppZ4bPXrprro3APudj
I7Clhk5OLcgoCzt51IaHOKIHhkv0mvDCcILGOlVcxm2GYEwHBhi9/m3Y7dO93jEd8dOQHccrWvW6
Q25vCuVjAultLD5719Pw7EZ8UG8kqWcKRmwnqtzRMViQzAgdhqo+8Y8TQRYIsqCXQPBed7DqfEJ/
YOtKjEvcxexGFx6YU4kuHH3Bx2xbzJwelt0ilqPt2InRUsjcfWRWb6HfVKkFktpgT+vj5HsBqB9X
ZNM4E8kluO/lb8q3PydHa2QvW3kPSTFusz/dL94XYAwg0DFxSR6NT+E+Zf7bqBavVZzKPsKcWqfs
C+Wmh/hXEw+amFQsqUW3azlgsyYnWJaCU/vlTTlQLBKJAsRvsq46f9sXzYXBEmzicYrcKVwJiyCe
yyFr9Jmdr4dZSTlaueE7oS6U9bVsLoai5N4RRauN1jXiJhLYmh8Y5kZ4XBsCae+SiCmnc9qUO9U8
k2eIDQ01a+IuQQCZGjxqYJNjuNGoXcoZcqUJvghehPhtqQBuOBYUteDIyEiD9Au0XaWOAtIgUBH5
Zo0KMgr6VTzIzln4h5agjw5d3a5/XBkvPoV8s07dd9mwUuoq+mqbsrScqsU591udIQqS0g65DICg
MPabU4Uq7OThneV7L4mmRBluJBzU29czBtFgRf6F+X3eBXvw7XqHyYCdGor8TXY104JU37OpbqWF
RkyCwKa2UjoSnwMGMAUup40TWClcF3rtgYavAY+1zbsUi+cm+oCaB3EYiIM/dCNoUaf4u0ESub0m
CK9KdKhIKKQO5lAVpMbMKbdtEsz8K++rkY0WJxPu/V30MQ9l2rr31+2v/jSKs1EIhTXYsifdQKgy
TOqjhCOzI8BR739k00JNmnoSW7UBg3DiiiH116T1rIBGT74/WRt9VqawX1hjRLRsjsrqssF4broQ
VsdsMNDjjHP/B0ju1i3H/rkpRLQvkPalY8yfpNiSwkwRCwYOKvZSBOGDfdHMtNzOB8DAhMdMcwN5
uneweVQPFK6soLGlk9Y6Z1mRqLwcs3TRykCgXeatocSl8ZTb7uxYrKj+zXnkqNYTA5HBJPTcygrN
8iE/VT6cTOfjB4WPfz0ahYPTNF3UHISBUy6335Y3MuJPtD0alUc8P9vtMRzRlkgQCB9gGQiW1AVB
cE3TX6hCadJR6O4alAexPk8lokV+VS1cy15ZT/fmloVETBb6avymVoXB4MnV3RVYB0xx29WJc0Gh
mH9eD2gYVOQT1fS/TENgEfdbw8KqfoUME2SI7aj59buw18BotQ++OOEq2FVJqKghm68UdMhD4JP8
7ZbqAk3S5Gcr0mME3iPwJ3AS4XwijOPaQx3MpDUYsWbL60SHC9hlRR6JlamuA6gEup+cSI/GCxDy
VIMddGZOvs6mxO8yYmEjiFFgY2KJEq9SkeLAF+00+OQjI3WwLMymesjtbojEGg2qLst7dtChXv0a
J2CmFnji92X2kNBNJ/la45ervjkPWtL1Oa/Mgn8kgj/e4VSztYDBq9CDlZSyuOcG/YBMfZMKLuDW
3klxATp2m6nMYpM4pBXGQEHp/OIp33dqYQ3EQ3IgYDeZZplU51ASQXdgIrLS9F8Xke068oH3a1Yq
tQ0BvDk4cBlZIp8qMAzZS43M5TQsnmAsPNd19SIn9g8JUddwjJPXc2WDo3QhVGucYRIvtsv2hXgj
Smz14AlaGWwbK2bF/4wVdXs5hudLbwCBiLSYSNclrDywla7hFY7i/XfTosGhL+pStf78BtIZX1Y5
uXJ0hXR7Cx1TqQ9egSHsbK3AYF+GfXAR41msdjIZh3X24qM92MVptpirv4RC4IMfpLbuGm0kmcFD
9zEE2rPLhxEQoygvOXwfykO7DGH1MTwTFZ2SXYQpaEcKqK1yHhGGbFJPwDJHA1goIYcm3QmnAWpi
6ReU/3rvjgFv0bq1gi6zeiMBonXU7pq8jIytxovarUxxLQX7K7QktZx64GV5zkj2DgML+c6JsxKZ
cTg8lpBpgawOpAXNKHrX4pOSLihgpS+3eyVNeJYceAkgU1IM+SrxaJxU08cd3GErCyFLAxj1+8x9
UaW2SRzGA6TCeKprLyRr3ickCDV/c3LxZ2SkfExwFi6pmXLXiaJs1AavwzETOPE9Gq/HfibhVz35
rhOXjCJVsZPhQFm7EBDhYjG2b0rxGGIoOT5zciz+pWSBlaRC3Uu+h3PAc+kaARUYWTVWdfCIoW/J
Mh5LQRzDv2f9tUuTfWmaxqjqeuMZE68TAkwvUNixRGUMGQwB/4ylr4cg6wfDbtKCKFrgIHe0TxLU
zPYSrrapqKLzSVGLH8s3VR7u4jdyPCCOQvS7lRuNdkSmvWxfZ3/AadDJcnbQXvbYum5YTChD0Nxr
WChSAvx9EN6Wzvp8KNtrWZdsbXyNaA/ZrcTbHYdof5EHCLmhGb+Z0oXMHxK11oG24qXkjuLihxfu
tZH9b/zJOwT8lB8RFAiGRnpIqCVmnx0F8z375Ufsa8o9kgm6/h5R3y5aZfoJR+yTOxYfaCTXtdpQ
fy48XCe2HtRW8KugDNgk7zB5eS14OrT6xnHYsXojbZY3u51wl0+l8fDiVhQ61MVEoAzbEWAKE8OK
q14qpEAkvY+KXTNeyOiBg8uUdkcIisfu6CNT+d09rWCSHAofxyWSzuazVx/3OP6LdxyBTk6ME8Vl
YHmyus5ohwmDEmVgUH/2RM0s3Q7pq6YURtQ/wGo5/plakYLMUA3a6/kCgR2bAdx6lO09wueHi/+F
/plo3IPoBtUHITC2Hqb8WlV+uE8WHjmRo4jQj7cTKH2h0qimrzVjEeti9rVc4ZkiiXDPM7k5UOpa
sZXK6KOuuSqxSzHqBx6rK6NucqGYxcOEC7gBZSymiWWDvQshGIwFVTh6EKrxoKSmY+C65uAVYD+1
lwXt8qbN5QeNey+MA4i7YNAtloKvjBLe9fviRorwxwZWaUVbeHAaKOdgXAK3Ux+KCze1HSNpIcbY
FLDcFrsoy6Bp+ywcedCeg1sikLLLu61LXU2FXIA+C1vcCxsQ7s5BeuOdb1aHfB82sk47a2P7Y0rT
XuHLNwva6vdwxHkghnSRInXS30VwkOWD/Y3yLEBx+9dTVsu72DVfyDIcBGLEHtupuhDCWyyAm6Ru
axtrPDlfXScU1dOUL0D3/Vk3ajL0AlwWwzxUwRictBZW1Ro9Oew5DqVgUZ7AnV0A+Icb1D+KUs2y
HdzhL4FONj9nObd0Tkj4OgQTh+W+a/AKlPELHy92y+kDMj92s+4/2aIB20+BuvWURPXZyajb5wPT
0uoSBOW2cEeb4S45D0ySEv59eazONphUg8mmY5yJl6f39xcEvFPQNF01LaiPktajmBuFWfjHeDhH
2z7heR0aKReWpuiOqlHRcElOTf+MJBgN7+GsPvDi5LvzGHf/H3SAsXoFVLRJCmp8YbPTZaCeQQUg
NEg9HejIpd64Hj4vGhrna1yD42mQPst0xYUedmEKWUENN9M2FMCov0+7Mp9FxCf0KGEGIXv9Lviu
kQr1z6qw/lTSPEBSICpv5G/GQ/tk+cilpW45v0If0HMzOJlJi/fJC1B9cc67au9+TwWbuX15PLEn
+0gSFwnj6eAmLedOuBxHBxaGZQSOj03zQhE7qhwUjcNg/kzC44Qw3WhSXZQDPCjb+qLV/S53ipzU
rmJGtmRWsx8Q3iB9hd0ZTZrWQAkx9icRU+/n3dgeG5nlzoYpewE+UDh4PYUFh95Lr5MqE/ynYG8K
vx6fUnQ/9v3ajVa4lx7Tdzf61yl+tDMjILaXgfMImuIsWI2v3HxBx/Q0UKHfMGZF/hkd7U8Q8or8
MS8VQGZ05gatZYPvStqiflzgMOPIqsuyZl990r27HAa5l9f9drEpWGZucCn47oWqeaTMIV20cnBx
B3BMbpeYSVsbN1ve1hrfbbUg3fXfpztwWfBCnkUF0OFAvQLBypYAd7KWZUke1Dy2WTyMW221Gfze
RYWkQHZHMMnJRLiTyR0lIK83l0kjVrZyeYSt/tBdMJGdfAgW9gTMc90J/oCbWM+QI9TGhhrWCdDq
cSswwdGT6LnCE47AnSI5Dginyph5Lv5zWaHPdeVD4l4P05N5ZxTnPSpgb3Avlz3c8uH4MEqaN7an
aAG0KZLob8qi+uUHHhz3V/LFOdvVxetVz6G3xuIXscWYlW5xBwajM1WXHSsqpvNj7CmgA5sqIioD
jG9UvrLNt0/UwTbRQehfy/8ySWJ6UbRnZ54OnRD2PW+nTNV9ci6e7pBfrOBlHqv6xdbYdaj3GFGg
L+PLSDSvPfb5zGa9WseE9R+pZybQ5IYbDXWXo+wpnbh2OBehQT+TzLt/dLVArZBhWl4kCXPufq8p
jqb87YTiy52ZjYRvfc1ffZIombf+oZte21Gnml1tagkh90hxF//E2WRR37CWBmFaNYWNaMG8GrVg
PaPWof3B7GfVkS2bdzGNIg9b8z1SxBaGbAFrMrrCEAG87SOa/dTbzRnGNhHlpbMMQybi8tDhbJT6
/ovRKgG8Fk1vNnetfFdnEcq5xidHVTRhC/M5MCBf3/V1/fkIfuco/Aflcb7U5jN2g1nEgzm8PAWf
3E/3dCX55P2yPROmUb4bGs4EljPc6nleVHGRR6crwpDd+GNqg6R0OenIcsRENnwtzrVPwPetwSrQ
68vM/i+wSspLEcMbQ3JTAa9NqNsGpwb4GYj75sbP7PVqR49Muf8dEshKR5JuiBxr5rb/Vi45gI+Z
440rLv7/i1JEYla9gi+z3P8VzCdpcrXyK/DwMnrfOPsVI/WwE+Ae3QAZLJmcWded/FSRs3/M6FWt
/RukX8jOYUEQ+5xZktLQGb3VjbUzDjgtnSd5F7ZRy4MEazFo+BCQqy88CJlB2i5MMXBLuLiCLuPa
J4GWPUsoA/XK8MH5Hq7bpT5srVERrdXaxzdRrcjH2uXpKpUZ4V6dA+LkFgMNHaNDy8YS/yR3TufQ
baGN9dwDeqs1QjPlx3xocV3c10qQ0U6ARisAF9vbfYLg5FfpgqVUVDsHprH74cwgfv8RnSeNxThn
utyCJzPGt9rAEzmOwYtuqHV1IofhMCpA6G9w4M6z7X3+RNOv605AShlMWzwm+ALt06L3VPYQRSMn
WMZ0EIg9p4/ocrc4Gq/l34PU0vz3ZKOw3ZLZnfe6B3dRRlTOxzOeGCr9pNsmE4N5cLRXgelmc6qO
MP6cjQG/WlrDiKfJRwQg2DmQstD5qPCWRnuZs0nBxWGhE8SSqURbLg7BDrKsa+MBB7xTD33R8Foy
JYb5P3lfi08ma4H1QGVYKZHr3mMjSltiMxZRtyPJKFBNPDauqrEx2NK5ZGIitTEe/YfTfyw9ofsP
Dqfcp0bQ8L8aKw/FE8GcBCPZqoKhME9b43JrjGVBKYgqhnD30wJc4RO2KJOkJc4CPoT7ebLEMdYT
wbuiw8H0nC9Zwx6cOZQZvyATZsl/gyaoS57Nhj+N3iy5Idi90b6yeeZmBvXZ6VaVx0ZL1zE2ooF6
YOcyaVy6hwb2gH+ZllzwXrA/suy7zBqXPP2KYduk7F6mxHF/0ktkv7swBY3HoPE4XojKYYyTNzfR
lvDPOCI9iGU/3pO0jSgfvQ8y3SRhobbXiRtgVnNK0ecN+dW3q9LrwXSEhJaMs0iR9X3BC78NFl/W
7LT1DMdq7tAbLfEsMakzFBqI2r4n7eCz+TIMn6cLgFO+sjvAWOTj/CtBHK1RdIWDIdcclgPgzZUn
6Z3DWfdgw9SsM7RWvamV0tTCPNtm6MuGLVQwpYkUBAWOo5GP9rTQC12BrCwkzQfV8w+PyJ02LyoX
cNIV8ofcEPC7m6v6aSAxV0nbMqJsW0UW09VvNnEN2WAeHVb+OGdsXJEKU70nXOHOkM98+SkSo8JZ
dMxcsTYLdwDo7JSvoHWzbgAJYbXD3x3fY9kJFgWpMRuzYiuCnU1IFFRY4UIbBC2q6m2HEIuF46Lk
xWW6oMD3F5EoLGe6kivMtaTSzXQLsjxZFuj5Qbqw6H9CuIBre69X5GfLtNqcBkDQJZ3J6GKbFKq0
nA0DNBjH8LuMGEg3nAqrVn+KYD9omPuSkdeMF29JgxvD3mkMh4URbXgS5eIoBr52xG6MEnxP9O9a
S+eXWcQKEON8kwidZ++qn+YiATSgTNKkmlNPw5kkz+X0T5QADNbEkdNZDVOy7M01fJ63e78MFf2w
sL7/R++ZFhtvy3vCMXObjNQqI6ZTM1RuJldLPkJB2CsFaMdGDe7qEQEHHRXaKMroV1VQ4xYQgzbo
gfSpaucO1AMI7j+a2fLdkc8HkeuCS1/Bjf6wp8anHLmzWsgi73kj54/9qS0RR6DkCq1VfJXS9O6V
P4YpcASBUi+LU6eZDkfwtaPgpV0EeNDsMRnTrL1nU4wFdOr4opPPpivyXH6ohmvleGbWkIQT1cHZ
V4ZYeiXtiGC/NjST1mVaPUCCOJtlfuF6C0nsAM3UkpIBYPqntpjDDH7xKiNNppwS9xFC51VZ1e07
f4+u4BsamzjSFciF/5G2TRCNJ4tfDWJ3JICOt0KE/F9mp9EjOXcoSBSRU5RyNGi3Q6x6Ks5L/s/X
coQaBdV+N/JLhS1CLNj6KuAV58SW30u6Fzj3V94IZbx1M3jP+sQKXWW6wHvNCV1zxuHjRk2YUec9
t/RzgkuGLspXeqIfSBFN/f8xkMgsD1Bjd7AJgHAUuLrJ9t3raemta2N+VwOSPyniSlYaOr5YBqUP
b6HHWoIJkguH6DTuw2Jh35pBk3InPwUkyrM7Hdu5SGG5dlFsmXFQGEKCPsnGPmitrPHE1wh7vkSy
B9GpMF1Rhuksj3UV9Pzs9A2m2zACcr4JEVCdvXBne8Vusw9SBfGy7g8jcjqxdJnFIXuQU8x5xPak
Ebgm+bK+rP3g4B5dLygRFqnj6SsBxO7ArYP2AXvwJhGhDFR9gpEe4AW3ywwvU1oe6Wc1g5l9RXG8
5USXLHZh6q4kT6Oet/oDy287dcsdcRcDUQFVx1B1NxS9N5kJo3khgThBOaG1C1rZTpR6APXHPfLu
4mpu9PO3pOMKr1yhKD+P6BPGjAMME9v5ZgUsc0ftPxzsFvNIwgXzpoUinwlc+XmFga5vvUJsSZ9a
hIVTSxtW6sULJdbS/Yf7lgICv/my70s9vNF98nwWoS1oUH1biCWqGOb1G8rmulZBUTQgXlKk/U6p
H8lF8pbKW90n/Mx8/xaAMzIk5Ccde2o/DpXK0Fw4qvEKN5V9QOMp4RZ4glE9IxrynrXdwQeNKTt3
iSzmPaX2N5C4T2/vAcyonQkEI8+nJee1jSf8q6fGeK9Xps65HFXD5JDwxAuego6CMHmm5Ic6QXX0
hf05D2cwHmwppdGaYtUGa42Iof0829bTflYIHFWV5LcpTXw1X8cJdUepyHzVqgw6CHXMNbaU/1mr
PuBzwZgXOb/34T2NW6oMvmmTcNq3/ZOSKBM1pkDLFlhh6u4kwdhS8sgCaMWBmqNzOl6LsXXt0iOF
UbYSQaybnov9P30TY35Qx0X5uwqDLr8hBKmZKK5vwq7hRbr2yL9X6WJedaHWut0ILMcqsEVYdKbm
wGFafVxCmuoGjScvqNGqEptc92hec831xtmMVy0sZpCsrY/vul5AAw0UJW1BdSJFmJExFQLbs4Gd
HVdNrULI1iKBod7fWqf6ghSd8D7GU2GOxl3f7Usk5SrXmVAyFALwFt6cewRDYIsClhXfjGehxXG+
zyAdRLpqV2f9ZzKEyctUc/8goJ0iGo36JSUAwJxSPyQ59BSFsvclcVds0mJ31zTgGdWpaD6jfg2E
PPJ5G/gEYVhgqQ/oWoqJ7DJ8u3lJoOfdE9kAiw4vP7m9J82geS7dmljCEhyivZBGugrj+aMwcMjv
YLYmuHxfjEIg6oAmMS7fEMrl/Czd6560yuR9gBTAARmbv4hsDiHUfkfh33jj973/+lnri9K/33wb
dxmSLRGoaL5whx5X+1Yqo3iA17yF96CRfiqHD2xfhTqFv68Y5/rAwYpN3OBftoO1WjqorIAiB2tb
dGg2uKOvOh0lxUFZvuSlriLqbcWCE4OWTuMYK+2oOsg3BoSCmjKboT+QCHEP/UYgec0FFdL15Xcg
PbNU5QOKcBm0r4i6B80XWp/xIfoew/H4S4qOsreBPxMV7FJjpBTH+w+QF6FdLKTlcZyMc3BNgyt0
8CTuDR6TYmhcd0Qe/3LGKnTzSCNX5XjtE2lEBUMNr3WpyUY6Q0y/t/jUNTDjn67W5TXfGoPgKOaA
2MnRBOeiaGcOqXuEtv+Zk3oWtwGRmW3T4xCcI+qPWXWdb09H/AWkYruAq8OcHFjIOdAON8tld8s8
k8D+DYQHjvacEiO8obDTaIIE6YcLQHDUBu9aSEeRlSpoZJTTrWcRVSRSeL8FkfkzOVFZlqv6/Rir
e/uj8rS+8H85WTxTs3FYeGfyNlSB/1DLBhlvtJOGUwSdaVqXojgzZU3O/ay4NIzRyr5IMrqKG5WD
XgNXitcTNVZRgpxwHY3bHT1nNOgbxGbwnIvzYN0ECLX8OFfkA9JP/C9UUYWPU8JXA4YpjN5N0LeZ
rUA2bdXPVmII0etUg2Fc+aUmufLIiFSifLxiJG00YSGH9KDPIPxv6M6tyXNLODAJQGODg96253ph
MG3W5evSxy0cRsgl4tFsOLtzk67yqVCCaBek+jBh0JKD6oBh9pAdpwmyU1e8YuFOdntKBjLImb/l
KfSPc3YRxuIV7jqXbeL8elVl4hLZ5GzpXKeOfNC3nl22f+nb+5hDYOql23zQQXC/s63vlSx0UhNj
vcBljmOBrwCsHdNBWP1pdKSs0342c+TWVWE+1Br4/ElTLdW7i8nIbpXXgrdFDCiCrcqym7j2ZwyR
XkUXxOw61i0QHzaFs6XbGnOTFkO1MjPL3pu0QYL18n8zEZgIXFnFCZ4joznyAiuZkTsQk2HbkouI
+QY22hz197LnUx5oWQFJUfKK94kNGhxG9WRgHMLEZRDIRyXRlEr7RaxRTnJ/ZCoc5op+cYf5aMWv
uIM0rdWh+p9J2ckLGMJAprQC4cwQt+5riUD6ihh3sZEQYG6j5CiqLDHoJWfC+sXbFGs0t5ERopmc
tjdqhm9+FfTpt+85Oq4s0TQQQVvbpfFi+F8qHzYGcvoyut0UY4ZCeV9TboE7fe8h9aQWr//DBQmE
4C8sAUIPkanjhhiLYLunTsj4FZyQeSbTE/6llG06eESjvpPZ1QBcrJBH4o6VgJLjd4bHz0oZ99Yr
41zbP4ok4p6lu6WFapYbcBf13mqSDVl9h6o6sE3Eq5cdvSbkxlM0TzWVaWmBUmjGnj+VLNwy2MpX
0ZSRXA/VNsJkYeDmEyhHrNU2WQJ+sOFvU7K4sKGsL96LFNEQDIEO+coAWrlPdWo1oWXF2b4QvlFi
xeWOGbmZA8FGcctY+4F9rIg1HjpQbduYlxOtjs25uaTkTO/YfyCRAOUeQnp7GJBrqrb1VF8cG3cX
FeOK3D7Dk0jtfNW8OXw/0Fvgxw6SAegmvGcoB5tv0QnGBzQ8X4i3WtDENtZ3OycePy9YPxxVaKTT
Do5YMv+1zvOZ5YgFQ6PECnlTvrq0H2djGcOb6qGLcm3XVEx+7yxE2Fdasrr1Svd/+cyE4N6wMAhl
X0lXZtXTDdyRnZQ8YBAwCxRHKJExin2l5w1OJiGkRZAIRGyAcFuNW9QOuP4n+88LYC6NLsfeDJ4U
Gg8eyTWU+v4s5xkT65CXJSBDAE+rKsoSMqBNIjd6YvS/hh75qzXjT3B+gEaNPjsWO6/O0GE8e9yZ
NJ3a4HnpLQU6UaFD6KoYv0qEsFwd+cECTrIFlgHp5QcDEBnGC7/OIjxnbuTdn+A/mOMr5gf5oehy
ZSCQgwqFlrr49NTdHzysFP0a1TSf0zehanpEslsOnz7sVpqb1YcIxj75iwt+xxbd0UkxdmmekCom
xb/8PiZmtpAnz2Z47aS8U3eqWFn9yg4wsb2sRc+C828wbuluX/vppaR3ZXqTjMTiyYZSvwswKkmB
biH6vX1utyhZQfnpQPXxsxmQKDgbQhbNqLLz4gRdzhC5oeqYutL/510jUvHqNfJc93e3oH4bASKe
XogBckKqMySJoXIu7dabws6um4DmOXa1wh4p+jiWeGx69s/K4LNl+oJYaXmwhp/7zvsTxa3hAOq1
KO+9eU2WgHtOlSu4JjTJAPdBcsIlZrcq6w5a3XfSuZnPfr6n9uakpCUVnvAjoBfPNWHlEMUotvbT
Rr3BhI00hlstTHxRvzojMX5BvjeOX2ef5OZY2L2qaxEnwo0MdMYnwVkZN8UdLmsODiWan3S9HbEw
q5xJcPKxALcXa533ILzYnyJBICidiqUecM7V+3MEzNot3sGpq+bz+1lTHiKjLb+NBIqZlo5gHo3v
XC2zDvbxS2Y2Fv1Np97iaG8IPFnbXgCqFMY4MzJHb7mDTWUjp+gchmgTPPDmGO+l2VlMT53xR8Lk
8J+1IAB7W9m6E53Lz7d9sgcrDDo5tsY7Za2zmucnwYbbJQ49Bt6ZLKhUwAxsbGmPGQduqOWB4GPr
7LLxmR2tvagYdn3sT3VebM8nQgCItOKPAjJQjvP8yCisOEam6qbJrUT9QdtBtiUQul0gfJ+kishs
np0yxEqeFXHOYxhPEL1w31v4j/KlprymAy+gUCof2XXCgZvaoS1lvTlts3DFhqOVtOzDtDubg+5l
VVGgRK9S+4lSC/oxAqS/zLXDhVQiNUCnQMYFlgClVoSQwOtIJ8MQFrQf/iuXQqxhuOJfdEYlOIbz
dgLoZwM4HHoeieHXHGpcNn/4SMAoQjEC8cOO9db2+DxoArFjP2qEaNdtTUUIXzAHyIPOJ3IkUCWR
SDajN6Wik1/lN6i2RErm6UXzOZz4CcVbTU0FS2m3k74mA37mG6xi6vY3KKzX5bJzJCQaeu+e9mRl
JZYK53XIcPTjYFkcY/dJzQZHtZyHQ0Cj92iZBHEl2WC+DIZfLXfgZWcPfGUE1SM7pAohO+3ezDJY
n9HQwNTc+uEYTKUxZDvHuqJyTrpsvG2SYtXTjKhfcti2JrTlwr7TKepRaaBGndM6MtTgFrTQIMAr
aa5JzWpVN1v6o3AgEuKlOpilj9+U/RFiy6ze0kKAlgkc5ZBG3KIHN4yT5Sx0/Cen3f/O7a8PIbKs
mwKcjsXLNe7lHePFdkdqCzRapHcGeKQy+riqfcNX87Bp0nJJDJOSl5RBnkZQ7mDv+aTmaSDVmF/A
twdzKxa52HzE9fR2RrSGKSEXpRfg2HINYRRXnyGMC9x5HAuYCbMCLUX2zbH1VOVwmiRkFXTdzRDU
8+zjwzkK/Hf86Ghxew6IaXgQilXFtAEAKiIICh1DOe7H2eW+OmHDgcLjv4sRqzZcP78EORLKoOxU
Qiqe7ISp9SdRME/CPde7bQk+pwLSY8fTHDrlDilI0nTY8pTnlz0IUuUjiKhXlWQfvQ3pcnkWyzss
tewrdMkuJHzKyCujDJE1pLJjp4nSsuRBY1kqejsLKnRu1n6BzlLdHka1xDQp2MF9ESM6PJneQZ/D
3/GGleB48LJSdX82lu9/M65vzlMLHKOfjjWQMTt1ymgi456yRLY3ssRMwkecpJpokcUvL0DsAV/X
Xvg/q5D7MjyguI2eADStM4WA1V4lUGODM0uptKXKfQNdqWuvUjIT6CcGjNA1ZhS8fJYRwiP7QoqS
WzqU5GkcWHESEXiL5cQEIauHp5aQ8LTjnN9C2pSebWnoM7M93dBxc/YFQDeQ4wgq1AGQZdjc+aUn
7WeEC5xi5OPvKKQyP/NlWGeR/Cyu26c3jSBC48Tpqfu3KB+YGBcHZEB4X7uvm+vkBxn+o4InemDF
RX0H3a6MoQ3RY4PTildfGSibYUYRZVZwl8jFHOMYxNxsaxdO9B841Z4UQJHKUUb5LvbwTT8M3+Eb
/JBOaTE831RU3goGiFJBGKotzkIWDr0f6ISzKhHivfXRGe3BgCpi4PWgq+xYadNKBJXBxp4yBS+S
em+4EodUYqxHKKnDVvKst4efBNi6gFfRyMjnnLSuoaRlPzKI7my4sviwC6zEvNBGvvU9Z+HZIlhb
U038iHrijXiCKkJK3OfPSBW9lH9PydfVQkDofiwOjDV20GAG9k9hLnQx4oCcGQxWVGtSUFkIPEQi
ZBYFrK4+dAW2CnbeTNFBAJ9u+aCtPGZqzHoy1owggoJIFoUHisGm07ZWp5QMSiX5PoezgdgtUbcV
umLOYMeWG3zjC1uu3O6ktCTFil++2nLRUirX6diy5Yb8djDs1D7HUp9aTEZ2q03mg5oWKZIpvTB3
7LoXsLnGu5DncYTR2VYf++6Ya01xmYYv31AN6+jK+V5LqvqNMSIbqGu9MBXdlq47M4BZpraqGDVX
Nz11zrO34l3MNUa0zSjdc2DyjYc+6nfw857VWY4ZzzaTObOuLV8JbBGNxJ+5s8bveT6qfmzyiGrY
xERS2bdiEV4sngF8NOShi/N3GutXV1qDzKnZDaZyURJG38XpvLuFvV5R0o1kp0HRfCSyxuK1olfI
MKWYCSxsargsiMeCR3gd+P4S4I/aAtNwEAUhiMZXhq6O5umJsb/vFARPEY/1V+fPu2dPcncil2SH
ENgGNBPbKgTiqDxAmUHR8rFGbAV9fTkpxSBuQi7EQtKdP+sz5IkrxLA4ff+qPyadnvXa8uJIpa8l
tB86J1EbCUYxs4WZ2wUsGQDsg58Fehkc5WEkvL6W2LWUExXUm2JdfV+OWP/G6lFolbztA6huQgEr
tWpFWAseFeWOwxkjkyDnSo0u3NYaU/QdaqA7e/Cfl2Jf2/1r1wnMjA72GkcteLQiuBn+NChRJPpY
V0vmzj6QQYbum4pZL5NWgjG5/GHtlfgzY3Poi4m2g1eVMU9gRdhKQJ0JdNyfPrgOmCuRLSY+OcY/
29YpJkC/fxzWZQr3fZJ1NMAva0UfJ7YRm6QBAnS8P8AKD9GpbCKdtYluhkP1C2WmwpZCH17n9t3h
B3s53K0uPxmd1s/mzJnALPOw2jSDoo/vYCJ0BYUD4mXDdxWTzyRtXROcH99qSV4lB70bPVyfmPQu
NxAt+UPJ15xyn3mHuY/IRo0qdMMd9EQT6kpQQ4qzaPgYnA0zJ8vDv/5G8JFDuShYyBaw++GJW6gU
tIJ6GxFaG/+r+dnVh/PDZskD/k2y2VrLpHbn4I4vvmfzR8YsEG1AyNeIFmcbW5VIVw2WQzAfwGGL
1aj6ywW1MCS8++Pjq6jzu32IgyCBQr3hDuUC9+/DrGcj8160C8Qn1V7T2xQ+U0TKaY5rnXdCbi/7
ayGvyfcl5CWMtpbfyYXNERWxiE85PNKZ07YaQIcIB4qexjl1TdmO8F0DUx8qwVYXiMTagN9mIZnK
HzxqHGK582MO0DzcUO9aeXFFKFJef9ROofdWfCwL/6uaIlFJKx9EPVEFHH72NnmwjEVHncNmFaR1
4T0+ccaeF9F5g2KyFEW+/B+3cDDMUjpR+wQNc3XDl8J/A/JUtu9jMjYP4Kax+43ZqVtTeciU7EUM
27y7uVqE2CCsdGqomYWEwIJ4MY1FRdU6cbsQ/GNZOBsKq0YiVbS58hSFR6D0qtt2MCIJRF1HVhqT
R8/Gwp2Th9Pi8fe8MmmzcRGXmwsmdqs8GRTEDgZiITvbwusnOVgOR7o0psixSj9C1xLkEgMxSo7a
pq35PDabKj9mQxwo2Sd6zxPh6K0q0naJdTf68AZlDNlWUwJnf3RxV4WqFbB2Ax5Fehba3zQNauuL
TVXTCLvtzxMy9T9wLbnzkQx7UGY3rEk2Bhl1Z5W9QWC4VM1A3Cv3DmZQZu1jqWELQ/IiZJGV7Q/A
A8SX8QO7TfkPVODsaBWUzECBB3gw1yZSyHMAJvqRMbWdPE9e6WpccUXpTD3zXofnjbGiJPbOS1B+
wqbiDeERBwc74ZaNkV7+kEkAL1sEpTL9WmmrCuuLMFG5xuetm9Fbk94rCrtRjhK8wArLeKhSMhg4
pw99vRmpA0WdDlKsjRF1Nq3WUJksV6gOLmyExW+zZIGAwUhTEzmHTAGzHBd2pJSkokR02Oo7vnUf
5CmZclDMXLYVAd/x38sPsC64GIE/75G+5o3R17v8XI4NkoRE9DRcOVHWYJG48MIpFvwznnFcYXA9
WXvee/Stp6fO+MtL+e4QGF1OLqO0ZAuVLpU10m9VCFMmwKCCMH8gdQVaYpFMXg/KiK6stY0GUiRf
T94Gw//DCiffqiZJNBJLM4y78r8eoDbjHxlwl2WhPxVokSr24MEUvRBHfiOuTlG7Hnjd9uWC9UNF
DWKajEKK5lG75L8jB8/ZTMs0yxWJT4olB2CH2NjnyZBlH39eCKvZRWRAymMryNf+MjVyviBlejp/
4/4uLruC6zr/Jh2P/alwBGFPkfDsJ9yB43THW7RRG5ERQT9h6Un1rpawcH+VgPevf4laCWXOqd72
3pMz4zPYB5oEy7nM8GZfxyEGvFc5cS73svrikotnoGFNEx+drO2ysdLvENU2h6r1HND9M22qNATG
MXOu69LqgiTkoeY1wVLmUK1ji0P1rPJy+UpH9BeqKG4o0z5cKKC6jx0OGztos1soVAeUNxiPxoxv
Eo1uphVfh3ZeDnGB2UzX37P1VLlBM8Asi5/fU4nt51JwvYAZ14Ooj5RyEpr/riqJNH4uWIwnyjeU
oMK6hlQx1HAcWs/KAkZNJ6iu5l4OAgjESoLTGZyCDLXCyOtKN64A7X89O50jEfXzhfWDhEruCNaz
G8REbCh2PeEwv0c+SxPTtSTI6bCU5qNMarTZwznxTCL1w/d8TjaeeMbPss3vO6eUIO0MiWYxSLAo
60FAvuRWrAe9aocPKHc5J9y33XH/1bejsVSV5MWn3whyKaFI2ExUZ6kVvB5ow8GWMUTCV+hhWWch
AtrghI07VNCE2/vFKCeKdcN0Fz7EcWvSNdSMvXXRUD8BiAk0zd8sTw+lzLqShdfe8oy8r9Y7JiGy
u0Gx8CL7HGx79f3WhI5RN/rUSAvDQgR/BNpzS5iD++CbHQnDftuSA0Tol6EmMgG0e+utTPiuuh1z
5V7TvqNJfGgIIb7jHFK9v8wzrz0eA0mhy8BEvedtZeBxmT17Nn5mrl7T8j+eG44fZQNbBHA0YEL+
UUceWUqpWSN5xxzA31vAvdrPu97DLvs5tgkQcAP9+vk1pZ1cFKPG6MPuuvnIvT/y39j8MP60zNJd
SWcFayzRvha6m7FKob/SKJo+IOyiQ++r6w+gcflQ7dw614T9Pwq/MAN6ZW5opPsq3mg2EQkz2shL
HePaxVurHVvMgzdM4JVoCqPkGRT78xhuLYyoB+C8X4Xe6xSUflevwKKpDOb7+jfudOlMf72B9AlG
DgQUHRzucWH2Gxo5FvhSi2FYCWy8WTMS61aTR3dLKoNKREJeW3cMeYfVZg/UoMdHezW/TLU/Xt3B
xunTnnasUJv+B73uEAOC4/PjsNamcQeX5d1tANpAjkl70JBeAUZ0zE9lw9KNmClg0Of3+wLa4NBy
ym/6/eSJwQ8ElJTJmDqOf/5aKPV6chY0bz/qfnYGKtVejOfkXU0HWDzdPq0mSmZI7IFW+eo65UIj
pSL3ALVhmL6QKLyzwfaViFwGjOxJ1RjQKsTtNkEoYn1MoWz83PtqTujQrilNQizE57X3ihuMguO4
I1h7lcZC3onOrg3Iqlmc3qsj4eH2yOnTXSLGjcXgA6XMcDB34zaGB9u8D2QL8va3KzMVxBZtWCct
yfg8/ppFWj0/UYUG+ZwPtWMnvqH7hACNGuGMlESgOVVTZ/JM89tAByS4kpiLx7Rnd8ECa6ca4Ehb
cS9ICqAYFeob1v3hVkfXZxJrlGnIQTJROlV/bMuYyePdHy7WZ/NHZ1hqARIWLI81Ls6vVfQP0Bla
zpWDPaiP+a1rnhxIe3b46F80fTn/Aj7sNT+2C8ls/KYqXaLujpHTh98i2xjm+WBADvpSwGG/rWpz
A8rePCZTqvHiu/793rE7rxPn7OrgP0fVYCmn4c/453rLkw8z6LbiqpS5Iv6rvPcEJfyKgA4GAZrK
69tBeACAaCTlYF+/6sLKTMQ8gXMWU5KbBuKlAIBAIwcqga5KwEkc9gxSaN61r8pYgi9O8aZ0uAsB
SgGuAfCOvCCcypoha83sAO4RV2kjZnp45JYZaQmfgCcKdFqaXIafZ2k0kwVmhzgA7TJYW+Q/9u/o
MC7PE1WfI7oOOBvB47ti5rYG95RwyVtFYq5tUwoG8GNh28/NG9To3ibyIwx9nV+8+qd/MfyA0oJi
1eksxKvxXsq+Cni1ZoMCikqhtM66MiAJ0aDCVc2aQBg8prFGu9y+/StrS+n64eN8yBtiOhhSzrH9
qWaI535HEjV5B0s1O3IoQP1aOHsKyKhXs5Q2Ac97L3O+qd/+t4px4KkSGhuRAGj9ZPCUBwXlNn2K
DAxhuK1XytSDEJtn6HCw5psw019TnmfDRosu8xMXBp9PT29edq2IvJfP0/iHp+0Ih/955+mJ13fQ
aldByAzIsTegfsz4mG2FeTIHgg/v3dOGyvFYxD3RSa1rjuPr6Ur3CSMhF2OHtG9wU59XT8Cjms+i
ARxakzdfx6mzSIDxBsy3WWr85kkuLaw4ceni3V0AUYeK3qbfBMclfZdLFgnVVN/bpbsdVRmXuK+A
piYaX2uJ1DoAOGK5BFJHcprerLPoRYLb6RyksK3djICP1gxC5lWuxgz+M+d4cuoD3KucJtHazND2
a3USvrmcUS70dNMsQdvmRvM1IVATtObQNFgceJQCVhT/Z3SRpGUFtx+Ebg3/p5ZAuqd019GYQ8SE
BV+qrAJxWC6JJxCWaWWSLsNJoZSWarZ1IKK5hovhWocB4KNONL79KVyplKlApTJbsLglG8OMSIPZ
sSZjUGtAHVmZoK1GhiPBPIK5p4T0R6eppnIWWBWdaWMkPtQunYiF72ZL8nVTFTfT8hTwf3tOd6cs
snWkBOYSNpBMCvULAeflIN0WF8WhlOdkyj7z/noiBwaYOh6/GiXUr2hwzUtpO0nL1WKqgQHtd4uc
6LnK23KdZ+4geYslAuLPDrynacQaE3QDXPycNXJeGUXjJFB4n9U3EA9/Xt4M7XDMUYHtmQLaGZKj
HVRrLpf4z6HuKA3Q4J5FexvmS43DbIISxaL9Zg74MUNGGvNNXWYvguLdt1hj3+BwM0H+gzRmN/Cg
QdfpamrV3hCaPytt8SpDll2ob9R9fwXAD2btqCwdtwVnuWQ1YTe2B1gQ6tdwzmVUTXZmzwpM1t4X
gAOkXRE0fd1dQhV1UqHdWtTPJTYC6q8Yd7CgXXnZGI5kYqJ65ffbN2FQ++0uQObrCzeNF1i3ni4k
YUXfup05HSnKB4bUHbZ/TXVe8Tqoj1UeZ7QEVznhE+LMm51tt+y6r0Ccw1ZbOOpFZTCQ/pVJb9rI
/hmMJqLXiJnr8KeyaOy1l20gbjlwaPOVXWf9vEahqOtT98aWSzkUjQkpGkBrGtVUsOaU/eGelQph
0ledaQrXMDn0k8MkEgo2hUOg6LbFeh2c1cMRyfwPYelCKMJ/WYppuqFy6lLQGZRN0HwHXmuTYZr7
XJ8KKZfQBEjUkQoThJRTHfAZGV8eX35AzNa0Cgf/IQBJQDs3IxqKbaGpUmb2sltxnWdObTH01tUI
Rc0/iRYXrtZcskb7ScHDvKjmAf2Rd2rHPyOJUYAijSu42NcN+4z4SuTuMPiMBFLMN5yZeZuukSZa
6cmuwZqDLUUznk6DyW0yqAPibNevApsd7c7mpREBsjeGKHeJwf+L0KS4bRrYGZ+ZrAmAZzoGIUyF
nsOPWn4egmavAhUVNHAYDfCGJovDCCy3VeaET7WVhXrRlOw45gH/3MlIwiMi89TUyS/3yhy9gYXz
7K3ndn+RVl9jV5ApK9CKH+kGxFVvziAadGFZyyzmGPEOyEJ2niM0FHXZj5XMWaODF1tREV0JyNXc
eCbADlgqRg2+PtIdE18ho/4pBt89pwG7EHg0hfPIJpJwVTyfvXH5bSmQQ35IRYVs8npCK5TisMhB
VT1S4NuHl0ocFvavwXCwqVhmbPlKQLhscYiGq8nOBxPd7UL6Fog3feOpluBBPHi552vXe7fgecLA
aHZaTbnPOWUmPeoHOTS4HwSFEbQjiNZ9K3yVVkOxVckNqjuwjU583KgZ0yjBkdG4gQPmmHvl/RGf
s3I8QlE6Bjxqz+UHiu99k7M/yzONUVyaYzVVGQdbfz+2feVi3GBU25t30SVwx+Ytfi/cF03IzlJX
taeeZfokscbOwLIDkYg05DgGmkkJ0/5A1eFzXW/kTFp1JpVnXBjRrye/ra7jx79VLBX+nC9YNRyT
93dMJWqAuj8L+fu6/QGMDj5FCJNVyjXbWRdPTISTfKeyOYNsqvo3atyFsnDPbGGgXd29v88DAI9+
0fBS9MkaMwrXiyjLPr7aBw+NKNAlOSl3IPh7E+LVdmwmZmlGGiIDXW0aIZf5htVklr+fYY6y0Rvk
z9/xeJPGWcj/RDKrkDX+BSapJsHbJ53NWT9GRfJbAamCOS7staUg/31O6EA7ajQdW/VFCByFwxoU
3G0C/HvdoRSugfcpxMKoyPZ6n+H/D7kncD507WIPKeWfCHyXUYoYZk2vTVSntfwwJzfbN7Ea5uH8
2N1sCiPDqTO5rQFNEjrg7fNJ3nQzkiOCMhGqLeylFL+dzAXb0ES+A0R2cqiOuxgyN2ARu5PRNfQF
m0D6lcLMxiseZ+m0JiN6LgDj/BGJ6A7o7lKyRGxXG+IWul21AH16vWjjRrrBx0b1aooU10p8VpGy
CZq5uWEhPJ6PSmnAmOG4U+o9QOgsrfxXaiAIFgTN1+QIzsdX2h0D8ORAbGdfEsBH5vGsvYC1uTkJ
eFc1/s9C26AHRFEAFS19UXhsdtsEUCzPvzQ3NiqpLYV0x1q8U8awDvJSzm77nPxKZLpRJAxJkw+2
FkvrE+3gNKyBE8KtRKNPBK/41nFGQ822dQFa/2NcKThmPZvYNYfLpeQAI4qVySduArvUxBeudZTJ
rVR55K6fjf4KXspqLNOlROsXCAV699by5I7U+xsHaXvJhEpPftGoeXgzt4JmeXIKSpIeKu0PAQEU
VbovFK4ipLiDQiKlDTPBcZaeCVjAqD2aVpy/rw11NfT8sAsq+LWmSMDdBR54DJGWT2/vap1j0bkQ
cOeHEko74CKobIuVIKW1lvFNhBo1Wk4E8R4zhJJU8OqCoB2LxSP45rjXsRg7YcQtHEYkKs1A98tS
xbNDb1BhnDgh5bIptCyHbxB8oDVnjUQWv2YVakmqUgnuRkqupWpNAhB/ZJEB43y3y4AvkRwMIGmf
PryTRbYAhcQkVbGF738x4OVOKLpuRwr2GbF2PLK0bYon7hwYT2E2bje1hrTbNag01nyaPyxN8VGf
D+23WBIeYWpFAnDLGAnIdNkq/zQeuivb2gbJyKgw6V/D5KaISdC2dZrqx++TKwExqLHNroD8hj5e
GCQ5QRznGW709i4hKboYWgEOjcTMPM4BOSVQpiRZxVXt3pq+eDcRqMttWebeEKxwlt3hXLF+4y22
fk3+ocR355R5s+w93um0tv7NLTyoCRlXDdbSnod5XzyiS/OBT3Hv8IKp7TK9uuSvUeq2Mxm5riCA
gTeKmY69exCypMU8K9OrjqMqeiA8/rgdqjRjPP0et9Eu6M6C1gKQ88yoiRurWY6A1WJB7hdjUTz5
kdF9L7k20PBJuTW+GrayHDXHxXD6FNZrGKx7B/Ngb+Lmr0iXAAxxP7KgThc/hVVw26Ud9o7yPTDS
Qvguk/DYQiNPZuk76yRavnn2PhLze1TZQcNJLr0a4abA0X9NSDD0J/0rekrAGpr2019BPoliafnT
qw9psTjuX945mkxZcACCS1Vi54RkMevEGL4dA7MZ2ApnHOeL/ZXwMrxpLV1DlvLKd7l6WoHJOvKy
J54vVM6d/xah1Qjx8Khdrg17APJmybIwEmIAhgU46Jdt4Jj630No2AJjoOputmobmjA4I/xkc9Xh
F23L/wYsF1cawUG8A7oiVSjurWtQw2oLCkLVyey6YhdLSl4I93SREiMX/Q5eIs0asU/w/rvzxIK0
1I49tZjr9weXf7w+HE6y1BWxImOCg96ptXErbDwDWCt5XGecrkLvTkxAl6IO2TqYi0Js5x+6bW0i
Wtbcqe5UezFJ6gdq8ND9QF3IiXugwrYHWf1dN78KYgAHpD4VH8RWkeau52Cch1mmG5BIoOgGiSQU
s/oLxdPeuTXP3Se6hl5JeUq0nZ18CTU70WX/74lD/ueeXIs3kOjliK9TDabHSXNfDOkogiW4c78W
xStZA7Vy0Ys9YlQxPiAvHafByRmRxLdjBMDwysvyBtzQ/NDjueUKcq7uGz5B78Nqdd2wqvofLDbU
0bqImt+XBNg3nDNzpW87N1SiKmj+LARdamvpBNGjoj5715rpOqdk7Etmq4e8gpGEwwHY5rM0fwRm
IMhNA7LRLuAyGbrJVf/jSxasQwKIaLPf0SGpcYDWRo2q7BEK0i0COLyxTA0rRjEVRp+zFuATIFg3
kvxQ2z2POBWl+gC5iGgWmeKdtcfmUFtTRPn1XGXs3e+3aQ29F5Kjc7s3Ncj5U2IkCgd9kzuFUDJo
ZU4uFcW9O5yc4BX9I+qiS0nNWdfLHfavJknBTKNimbrVjhMTYgpNlMIYbHalVoCJxx4zRsIqb8jY
zMxR3p1gk2MKX1i6a9hBvoY7q4mxrlCw5kuuX7lih6pBt/T87y0BouUUSlx6A7prYCXnwdt5tuBd
QmROmtJ8zh2+Lajd94+DiepdAn/StzbwbHTn8a+3Vf+6Rxf9TP9nRZRj40WESuKYBeNdFQdBN6ym
HpU147KSkw+XeUhwf0jeHkpxrzGagjYxVwgHiEjapq4E5zctpD14XdJ10fOrZgkvwNHrTc03X0lH
jfQQh4GNOzsvCN3KkbMo61lsZF5AP67m+Mcmgc5jjHEIDzesRK1SS/SeUua3D0WAF8rWKR296i38
qAyKN3NeRNc0u8nrwcSXdXmpuOWGMko0vxONi35BIly34s+cwlNZ0otV6oHwFVUBWTEF/bJ0Xska
vTnQC0yEuWyg2N8LooJTDyyWjr40eIE24kx2JUcCechUBkTKRSUuqq1I0p9eM91SpKJjoAgD5HTt
rQdd+lkVDLIHctm2WEy0iXLkXPb87hHhBb90AJZ0bx9XOWY2B7MTZVB6Cw7Wn2oU82ACz1mZ3XxM
XmObtvKe2as1ttNA/oUWER3DiybWX1Gbd5Ffxf/I+XQcZjRO2fpQUY348aP7NHPN7A/lXq9jouF9
lerYO1j0P238rTNRfrmt3yg3VjSKd7oAH+3C39mWncY3Y7nsFhg8NBckT59BwIf9eRzXFVdmzkmO
zgV9xyqTo2tfUi0BzLjt84fWRy4M8IhOAlzJydenxzj13G2dHTNJxRP0uSRVc4x7OXzEMcJC7Llt
BbxPqBBRbTH7A9s+dpcN9ih+AXUxZmGS0Z+nvC+OeLzjo9/UwV3uJFgmA0jwnOFQ8rTMOe+svf6l
eiitGih+l/0JiXaL6OCNLUNmK/YekThSO/CzqB9Ab07B4idhVUdj1PpniWW6ZloQhP6WFCnwZRbw
DoVVl1n8UPqmytVBVjjLW8Ia1VmpYw4qOdGStRXXJ66Nc811LS9ePBCJ3IQFtNDtqSZgjIlBVPa9
NxOtDyb4c9NMpXpSfCpIdMF62aNtomRyXwI0XqFBoDcOybH+1GRW/BabFdXnz19UkyEAAHrGGorN
nyIDbhAoG6A3ETl0EXFyxr8n1j9C/acmRbwtjawYZQFdq3GSjsotSoJwcr95LXi5YBCdKRFppvLH
5g1Xx8OnrQUdueV9RIW55Sn1M+YvP9OvahjglQrL5TQaluEbPYKgRZu32yue9tRFeyHY7xDaPWTB
zG7rrXkq/LecB2xKYO6xMUpdPq0TV2CHzuxVI5JPdyqRYJ3qYvztedJUNu2JrXX9CF9uXkXgHPBH
YCyUtDCxnu/p4E8FGmLvuMhZMEy+qxJ/yqgSW02a+I/uHTjuqTAq8ggDteLcSeLb9sSCbc4pbdnU
VhC33Ym16b8W2rJVG2q/mV+zrOj2KwsH4Jbk/yc91DVGinjbps99zDCZymCy5eGlGyvufEMDlu8m
u+ukeXsdjOn2hSWa6WJ7q9wDLvP9XkQpAhYd6do8hjg8HDtAQLo/FXboHgv22iZs5VUEfB2MlGyg
SGbvZm4IB7Tg2+8sFs3jYT7aC5eaXqK0wqa+sf9Pzyxe9d/BRzuK9H8ysKQDqZVtjcyAKXSVXek1
zHRiTRExfuE3aYZtWZSeQo6Nzqnl2hYXEIBRZtiy38sAhYiHqEzFbo4A8Eur1pofBUYy+ZMs0HXB
P+/e/zM3eYgcSVTnQY9e4XNb0hv7nLuXQWEwdI1JQUZpzOs7gj30sN07TcuGZdg8oxe3YgM/F0iO
6QpPAI3ffWyznXHrn918vMAD2WlVNM+BEugdZIHMzkigfcrPY+BsMwRl6rgOqUGI/059R6O99tnO
0AH3SvFfLu6787AnICnJ2gjlKe36N+7N8SnL9XwFzvcsMyJ2K1d/nBw0MNhEAzANSDn2eUsjc7Lw
YMm9/Tl/grRUaXuWs20/FOsY8jp6EqYZjxwz+Bvv4TCz8/M8z1nho0g+Udl1eieE5+549agZBtx8
pN7ykkzl3cRnEvfIWH17WQkgZJHB6QbXGfiVX2h8h1v21HLQzEkAO8LsDQLb/NDGBId/oYgMDIBD
V9SUZaHimDhpSlZahMZ1WgjqmRhQS6Ko/HXCBzgh3ekTdjp9gDMT22zLarBgydmAiIPXjsqKbpQ7
pyyYKtVB/u5HTqihTSgUG2aKS0vKT8+wSlAB0gVnQQEEhu0G5We4MV53iJKLGKJ/HfjWJl+gyRPy
zXP7Tg6Jjwx5PQv5JDteyU/v+S7TnTVGm+Cenr9JUb7LJxR59TvQdIEaHFXU1MKFgM9dADiiSOiX
N2H3DCrLt/T0Wg+y4+TSEh5XvlbVOwt01Xffukjx4SwXxgO0CEIok2hUFxsTnWP1ZRimGZcElXKK
myLlEhfNy4xQw5c/K0GTm29vKXnIdzu684E1OGnjPrmLHMz80GERYXJem/4usefLaRqM9ISbVY6D
BAr1heL36xsH696yYXsEFh2dKMEAXbX1wJCSUIkhOIpNY/rdJgtrBjPPQEjRYpOJzMoWrNpyW+4U
E0/MMM5Mk7DFg2oXk0vnCzqxEFhLKIYZ7ky7SiHbANpsc5QxFptkQDu7Jjjpqe//pmc/rm19Unbb
tpWldp6GQWDYRbRSWlEX5m3OJEHOd0RU9h6OzkeU1+rCTKWBRW291cutGro10Jn3OJOl9uIhWeR+
+pBY2+qsjM7Qqf+TpniOiZuxsYnt241UierDHY9NN9cntVWzYdjZ5XXvygaB54/qLWH5RuRWCMEz
cQJBuVPJuDP1T403ra92UF3B6uqG0inic+caDScgL6plWgr7vt8S9mKKwdDsrS9zvSIUF2fT3B9m
kd3bktT2fw6stNc93QfzgrLeSSHQK/dMZyZkJJarU+GE2AC7yVYeq97dFccRZrDbABdYAKDw8Wak
P88+UQF6zGVUQvieJp58V77oS0a6z7yUFnZ0kvzfy6lvqwsz+38/zpWCCH8ZdZTAcXNVzFS2O6cX
NI/9iGeAHCH30O8dwjJgBDyvc/t79s7Rfqm3MEU+nWf6cYhq7SNQnt/0y3U08x4aU7UZv5NGmduK
RrXi5IVlDM0kV06Vrrzc6JcrAxLfWcqJ3WjNSEXVLGLZwcBCB3/Rdgdrp1C5kyGLDJS9gymFuTT8
/2Vdp+bHPkFk4BHbK3/dTb9JS90fnFmMWOrjUV8xnnqVkowWLV4fwFhF0sjNMLYnaTVNs5nrzYhr
v/q5M/j+pbI5fqu4MgTDhwNT7oL7xBlZAHKfpJIsfmdrBs/vvXGQsi5kp6SXB+6iDY2PESD5FxNt
deAXtGZPTgzcGCPxwcLqLfmHZdMp2xICJvCnbxAM3nyWlazqR7kGJjEGWUVoKyJv+eONYeO+gCnc
rM/8Jo3ISBLHNEPOxTu6rFBMJFl3R0VgE5rN71Up6EaHgzKHqEUoQenkk9YxQ80E3SRh4bT4kov1
4zNDlae5P1AHGWWTjvFh2lWqVAWV5I4A6l4pTGzBA7S/Htun2PNGSrG8gQsgBnN+fL+AqwukcGCx
4mpgmX5vXOxDfloOFWJOSI1/g/wVrX+jAQf7R/5A9NSbYLBUVTbdmI7gehOCRyFS6dPawXSxLJLu
uXGN98T+Neq60WegjVNYQuYqWnHWHPoAXUSMx5L0NvQbevjDTXvE9H15zCpBNx0mDOMVnhIbnw4F
tapfdBxl/caOQxrd9k+qj0K0xvWiSU7JjmQW93Sia+CJiETjK6MfWzcnTCb46Ha5WK1Vk66OJGMk
k9X5Q3RwoGGFqEFUIh0lHSV8axuu72k5KqqJb3PvaToXHw1BxZxIo0ISjAi77sOmPGe6txcOr4Sn
b72C6zPo5WxszR/dozSuo8wVUDBhyBleGf3CVfuB/21MnAZmVzinjDMrIT7S868heaIY7y/H7qTl
vkteGfvY3EvJpezXU6TB0g/AS7G+cV5utiCs39/V2dpQmJhPJ9PR2D/qCEl/D4Y0wl9+vWZgm/js
SEf8m0duVeQkhc/e+b8FjUn5Gt+/9cazM33qxNe0AeZ2SUvidgnOAQSddaRDTMerRLfYP+cre0Rp
8UwwNtuIehxWooB8lSRvrZavJgkSaIGvRXC4c5Ejvsi8BlAov3onB3e8CFMh0GiYyhwusVCYIAR3
DU51YS4UNm1fG9jPArX5YdTIPxYo7Oocc6/7/vfnitR3nWB5Zfkl3UCWQfvMf8gjrWzicBlceLAP
NNEjL9+BvlG/IZ6mOj8cQfK9/BjBnTvYXwrDeZj3TFnnOR5jVZbRSDGuiqeu7LdBKmXcFw4R7ZIl
XlEYaJN8SEGgZSWysmj3ApYgsVxOX8I8ir3CeeJMMqt1GmHtaSmNsmj3sWhgN+88Prwoiy/g+U7i
zd7aX4oRLO88wRRouGeowzGXnvy5iBIgfyBsEeG6IR2ce3Mle1uyoemSC/dCiWLNpuclU77NpMAA
XOeg6gkkhLNueWohchrKJPDf+cQ4nggsRm1dCrQ6qnYHc9zx3yTXw6zSw4UAbFtZybGUc3jLRm7v
o8pkWoDWIozxYO/d+jE3Vp2ufR2oHNKlD6BHtMwM9YPlypW+XCN/H9Lj8Bug5BGTQiyZYHCYTGkV
gcb33wcTqKT5aUM0cdPz/Gc93pQtQBFiRjZTvni9RRwzhRzQucY2EDvelsLIkPJlLk+LeZSvKe6I
FuIrJllCCP8Z8/pOj2xSmGz7nY1liyukupin8xhWSsm8lTbHYN03F+1jrZgLlFrcYXVNBdoKXPqB
98zQlUlzfXuRidTvy/dgV79I5FQ0DnKA+an3saNlVwKWdLXdx21w8nXfYBxPVjaUVRnPPwLxsby9
72Al9lo/s+3qOzzDjM1YGfVSBGlYx81XOe7GBVLr8gUbGs9/HeqB9H5jAw/hHHwiQhKid1uVfkt4
iAKl6Qm5hr4aOcdZTn4Nd8uEZQR7ekYmjOL4qTP//kmV6HCg5a4jHcbIGTLYsron8lGDiP6SZdSO
RXU3DFsy9xzAt7pz3THWGJ3NrWmHMViucF1P/m7Qk/51rYmDCmW/eWY92zsptGwd8IME7X3TK8vt
IgePDnuSTgS7aV99pU0axvTr93+4Oq5AKscCjvEoUg990iSOGWbJrBNEMp06/qexEGnKGm71Be9w
2PYsGE+iqTYDYZfaWfCN12baGtw0oqCmEp3UEZyipSB6Lj+DTJsue6fxXCWrPpcYMSQ3RsEHEpR7
Nh4alBu/RzEO/asSMlwgyDZ7qr/o0Vv1/M1ZGaBzpC25Vm2mZb1afyv5bbiIQLqwxZB4i8+srci0
QM/Iwc+MG7x5cXJx3coMenKd4G3UNkHWilfpaehS7Pc1WwHi2hJ2dmq1Buo6mQlXAMkrBSBwZ5g3
Cm2Ru3c3WdPbtife0TbYF7tXOsAGjUWeXMv+P3526HOwEk/3tuJFgRljBq5Zb/8/be7HF15PmIUb
AXiFQb/INDVNVG24DP1wOZ7RVyFxcZz11Q7mFwF1m9XNrX1rJRdYz2VcBVp8m3FvFjv5dUyZak8E
ppG2DwFh5Q1J2SDoDh0Z+SVpKPRywuMEDDw43yfrKK77aZPf2DIWcnsQdUZRQvjtm0D5bTGeJ823
R0a8Mvr1gnkatSxseyhXoVF3LYCWTh4xM2L1nIHvXzgumcBixotxTue6ZqyqsTFjmsip1QcZb3H9
l1jDAHxqoncXrAm+Ss0gBYOKU7Xqr8EVQmWRCDyMFeV2dCS1nDdrg/6IFuinDOk1nXKnwSntW6Di
IWXIS9hSyWV5YxKwDLfDQwnPgZIAsY30jCQsKIuJIOxRnB3Dxv36yCkVobGBbKwxEVqf0AX4Pe4Y
pd2QXfcxXuvfJKYGGyGFipyCLhqL4KJM+iJE5B6qHLpxnaW1ZKtRExmsXf0L7kmECHWbLUgYYEvG
4GMELWkHYzGTj6+w3Pts2IEob+BYV9By7W7vqhbP/G+2kAp9t634LXxugBH/SbTQgSOSvCa1JxhO
MVP9FDWV++wP87h8/jne4ZC9FcL1w9UrbT9yIVEEafC6vNUeSnXchHQDEJHHRuLH/Fp4dHJcIMEh
F1YoqRZStQPVVyA0izw5Eqrh37oZiz+T/WvP/dSwCmGVbkDif5tiviUU4d/RKPzU4I53v9h/xzX7
3np1OmRoNdfuUJ3yH9P1j+YsOXEoH5NE4eQwCQTIggy0+ixjfT+ecbx8cxyYc+z5RvmrT7rP2XNg
DLTNRqzJdpYiFHBvBnGu8oDavLi+9VdGiVw7qB5KtdLpvHuCbzRGVMYeglRnKHZcOoU6GFk+z2UD
vYh4lfEl6fCw5vYj3BEp+TCgClUJnE6caPZAQ3NwP/Q5zzjcnJaAY3xp4IuJnDAKGiQ4Usjun3v+
Dh5MR3LFtJqWgLdRi1irjwikzRXQ61zAuJrv1zOKGKL/CiHseN9g+QfkP6oGrx6hjrC99QqGjc8X
suogZ7xZQ+HA3VozS0J7w6JgZ0gavJu7mpbdMoBrm//z0QhCMUf8Dx7/aaa2thFrXP0Q7ozQA9HO
Tjsk6DhZRSPo4DvtLIWQol+fhtL/36au9uBqf15i/mTCu5xhRV3wxASSFVl0SPxS2UYIUYfh7AYp
BPlqSxRvTXQKeHe992UJbS6mvbJcY0c1QKTLyyhWIK24WnkZs/KCZVWhK+I93u/XyIgUPYK4Ht10
WT3mt/oxdkQCXDq/Yp8TWr/RrzvnTd1/SsLukPnrz2eWTp1iYWPjfS6lWma1cYG/8W0wBo2grHlo
ePtJLVulzJ+T+D4GYarz4MKtBxdIGpqZHJS1Rse/Tu4I0bbeXBlHE5WEIWNlJvjxyWYKBK9AKfUv
3KeQ34rWneG3woBScTS3b/3j5VSQUlcMabhteGFhsrCXgu5hvtNLsqZwToF/zwHB3Jyj5aRC4Vs+
/7HsVS2xYryvemPJtR281Dy+UlAfVPGwzIIyp9ucTe8VUt/JovehhtOfcFzyW0b1YKomPALGmrLF
rGPnnxE88YiRRo3Bn/2ETWKMWy6NJbweJ+e0nYhdTdPnBpJWErUZqFuk1KV6Mo2ZJj6vYpupROL0
zTSDsJez1ukEOqjzG9Lkqtb7m9dRXpwRsTznE0WcEEKF7jiMrvb7zwjIhjxMG4btZOJNZDnsiCF5
Dd00hkBGt7gNO7y5mDbDupEm9Z5e4uZ6C6AlIaIG/IwmCmv+NZEdm4RqGPNCYL1H/pSaU1OMCF37
vuybQxrLgCG1CgvtzHK2wB787p1uT0oncUJJ5jVyng+xZ83vLsNFbe93FXuFyyAGRvVST0Zenb27
Rg45SmxZ32QyM5vV5E6qqH1n9ye1Z5/Rhzx89c0CWJytAMqnCyRQwDINRFPLBa+61AWHrVwYiuNK
kBpzUMs61O3Cwpp245A3z1gcDrkF2n1rDW07JljffGAl1pj+gb0ZtXccQ03eWTLilPXZkDandQzr
zppxIXcR130BWR3sVkX+JbbmHP9k1seniqmZJWvIggThWwb/iguY/Q43oCbBWE+2gW9fVWKTVA4S
NYio7JyIW0YSLKLiWFomcMA+cLfqdjfmOuGdEZfC74CQ5TK/HrBCSgHzdTLtBrAdgc0Hywypg5p1
MrZQfJCEzCjP5Wlf/ThVTMt1TbvjDYt5cQd/dXLHve82UC2wSKbj/60Ym/YKVPaYvTTDsjHc+c/6
3nQiPPb46ZtoP8RmPQ/hm/zU9DMaoqhJP5d0aTdeH+4kw9brrOREFkxmfX8PF7QDGe6L3UJNW5ym
NSJ9vOQ8LXB9wq87mJkOZ6kO7l9qm7bQ/tlceNdWxc2UkY2jWYVDt1whyz4w4p68mnfmUXVFibJm
06NH7N440WdfPrfzdsHpYOGgemhBHAwYdinEr0P80ya3UOIYavPqlmOyqzNvfDN3bVD7PiM49nmP
HdqLDA+sK02jH1SnuNP/lgij3tm86GAJA3Gec7kqTCTiF3l1enz2gBci4ww0aL3R+yP96AzCe030
+MzFKw/Ukb/Yo6Kd91iKiyZzodG4aoeO+U5IwN4evtrzOHKWfahfZueLLYt0Z6d+S87K3H0+wZpY
HfbUWBd4203bPBAYrFja+E+cdhZEU9VxDzt4n0v1ASOHDQG5Y+BMyxC3MB9/xQvjVs7qQMjU6PnD
AF5IUaCs+z6kC31o1hhYZsiuyzNVdxW516Wkm/iC1/05MmaNPqa3pi/EID//c0aPbN7tFKa0rTTm
h19ise59qMpm+MUActSQ7d8Yw3btw4OdL+9NhQawzaaA4iLEP+Y7JMAO5cxTyi02HUB7GuiLh0Uq
FKIPFhpwhoaoA1m4pCc1ItU2is3av9/w+Lg2PIE46s0AEFsUGvrnToW1B+IPXH4L/PUFO5mRc+MM
VGiOQ6hNUBKdaPVYr5QokVvoSujd96gebqgxzPmfLM2AL8BaxDr0g3KA3yaynX5htHtF7ITC+CBu
TSeK/fM7F8oHpyTOUBqJkKAix+4c3k6IlFJWf0D8Qx9dv//Ah+JbFiDeVDgw2wpov20AUdVT8OnV
P0cWOKJXYBCz2jHJHDnTugbjJ8PGsxu5ZHJyDy/Wqxzcpw/ckfOTN4cwwQw4DKcvZfXgAFuIL+lB
8/oKZSGcrGBGOzo4vqxoEPjmSm7xc1k499avVE1gEBwC9Q4jqK1CsXN3ZwffIhkpz7AIUysmdgk/
yqND9MISy331f7/YgegeFUU3qj5e+g6o6WIcglwAmVzDC32kKK4HEdskx6rS9mCmayzs5rxFVkTj
i4bXxo+3yRmau6B+YybvD3hHoY0lC6KHplEOurLN1VoASlPG+tsPjDYUJ5ekDOWg4PS4ffbi2cL7
69grBo86PMUbjmNiaNed5tdXqeZdCQIIaY/vRwPNuYGY0VBxxLXjW6nuPVVHR899S9d/g9MuX9wl
nVC9H+nd2658XuXo5W2f3XzzWljp3t0mmriJuBYOCevDIh/n8NadmCsA+EOONwJlwGPFkJuoBzY0
4YetVKHCNWoIG+ispPjpfDxfxxyqWHzQhjTCppphcdTzkYMMH+S6ZOLysMNdLDUkEeKod+RTN73H
clNRSw9iC2Kfr4dJ2vBo4AvRp5q3aRqjutqhgm4n1MQt9EM7I1ok4MtOIdi/O4YDPnrv5KKFnCVO
rF3h4ypdpKW7k1tSo9cuTWLAvHF1hFgp8qk07C+b9jmonvf0IcenhuDflRonrdpsOzoZr25mg6U6
/jMpaHhFiHrHhFZgXQm3oRl/VwWT/bJWNEDEPTVUwpabNMJgwFolxhf1B3D6MYhlES4tXoRNTVks
lPdW2rYUnAY/Z56conzxTH9aYDAZ1W8wyAxnr5w/4RSSSsXT1WhrMmgw3suGbTfJrrO5HQGmeUJk
y0eD7UiSgnVOG/MbCwAbV9QWN6soyLRMr18oDzAiwjgbMI1bhStR4dvY57be1qGw4aQH7d42yE36
n2PiOad1pZD+h/A5H9rdlgDQQDHbHmYtm/COG5MR2xop1ySF+P9YjtDNvfX4B2c0bcze2WRS4e4z
kS4bN2LLBt/dxcXMeTHw5WHpVcO5Aj7/kRYJ1e+TANUHuddpehNn3JGS3jHD2UM7VJLtbmwGqv/Y
BHGZbx5hA2ebnD/6m0+Wta4Gt70o94EQREf5rLTnBXLrARGI2lO6069yUbgbsRNafiiyb8nT0Qoz
rh8hebaxvStnYEWMatLO/A1z8ps9CSR/HPyThmo93PwLaP/aEMz3padw5qrT2Bj070pQKm6vMvq3
bC/FW9fSdnUd/PW96yDfdbs3rku/i8T043Ix4FG0zSasUoEvCOFKaXEx3yMGaJmgV+YwX6RJsyB0
lr19JuEc4U1tac+O6INq+FUhJauxJO/5+5jV6di5iF2aDlIX19ZeNigr6jLsCAW6TcUeGlYa1rYq
5wmr0EF/QMqeNoKZmPTBXiKWCUJV6e2lXb5oPt1LEKbEhYT7onGbkOng8EP24Yhzi1FJv/lkuuVI
N2zX1wtmOK5BCgbk9LQIdYwD/5t7FzzoBqVufCQ48svTubt1Oixfh5CBjJEMil9KG4bZWed1bfE3
F6CDz9blvMaCXdH7H5h+7UqP04SLr69WBdZISNT1mltGAXTLu6rI4K1FZlR0U2TSjhczUy0HvX/c
a2xu8aNeLRLt4DaLNN8q74rtNlsm3ezdXoQFcZU63A9U1mFIurf0RIU+y0KnFrLjdBfCJ3oHCuFy
WOMldq0xbFdtpjWi0SDdUTYY+WY69A+mpSpMce4zvbonI4/IHpNeJklz054kvGTEJm+7cDhmKElh
wQoKI+RheJzyu2GKmVFdg92Yteh7YiO1JJH/NIs8BKQvkzaaK7ekgOdh0e00BpMYjjvmdURAf0w2
7tfqzT5/nC2MgX37eNtKDufLMez7NwLZwqLWTEWS7eMg9NghKFO15ZgpmYMZdrX3DT29FfflF+e2
8OsFl9c6wf2QsYueMYPLjl7tuJ3t+qGsX2JGY55Be21ipnwZaHKU+OlvDvL+U1LY/zZpcbMCUX2O
/IIpiiOJYrUqxARud6tWj12Q05Z94MRMDEbpMr9nij9vazs9s0yH6ZHRYS5BdVXzUTVAdXJHkKcI
NC2wUAGBcAjRa06yT74DACisRC/C7fUhXDhcUahjLVwuCjCcee/OnNPLZGj+uGWotXMW2sWRToMe
yEGISGQElIWnP1PkGaboA41cIiAluVVDqub4Y2wXg6cIWrLIdYy5jLLGN/6bsS0RKEKDft6bL82A
wIh8Nf1/j94fgApJr64AYRZCZbYkWvAsdpzo/mk9lcg6sFrhbrX1EhaxX5h5a/b3ArA3wlMLoGkh
VATROfGG0Jjccgt16n6a7tncs5AzGJqE8tRAXZFTzyWw2Hb9BKnEDrZzGhQS0GQImNJSk7Cxgoee
BYl5wf0WPpgLcqM5+ytdQKUYDMSBla/fCmEysWe3OHSSGsV9t13mZ8zBee9QykFhxuJh9Gj0oPQ7
3eClXHwmjL8od2Tf/VVQFECtFdcHOnWNXW0m2LeZv3fOQQAIS8ZtwjFUENWi4/CElrjIdQQU+OZ3
6fQPS0i3/XB7VYKCfaSiG7MB1zFXzSYcwSL5AhIK4l2U6AVd0NQUHJSQm6jDaQUk0oWx585Bsobg
pY9b8kfnPlsIAbTg6UwY/gS24hyNs7bncoiCEKbc2CQmvJ643xhLSEZygbxXGU3rlGbVCvW3NRyk
mdSInTNW5QVciyoRsD65KN6jQYxNccJfwe/eI7biCRPopzTmSqGNWouVZPZ4F9goX9MLDMqN2FUV
Nx3Ad3qq9aT0kRgSSaY9q1256i24+j3CvxkPCU4YZL6zaY/kO3CL/eqAouicdB95eH5iUdyzPcKg
2s6J7SvYQYsoIZakhJTomzMqd9zIRQtZQHRxgZ1k7u2tDa+pOiiQK5T5v3/Wd8sUK/6fBBem9coc
MWgkG75Tpm/f9ZVFzqrqP/ARz5Mvo8rheZviGDJa7MHZQye0CRaY1thAXf/upzr4SteTgFmOxQji
toqcnwjGy+HVq1rmE2hUdka9K/b1gMR7CbJqXZHJPRNfC94+rtDevkQ8Yuf/CUJqbsHS0znqYUeL
OYb1DTMDmm94/VdilpewNBtzeOkc6mYpDgB/sxDLbjwU3oTBbhirBACAmy2eN2PWwyX95hPv6eIb
18qokjA/xpGqWWhpjg6GLBz4TYm5+5EXdp0WZybtsCp+UbJfVdv+wYpeoks2FLm75TEBuXfk6dX/
llT6c4/etLNZxpQ/vNi+TdXXbx5nn16NcexVhMeLGAwPfsFz1e5ERBOIHp21hSsSzrNCvW6JBGRj
xSvktFmD41RYPI7D2UlpgZf+bL5yfwAP5aHh4wWh+1iap3dlvBAGUAAPmUgxYU0h1lyTBxvcz+r9
gCHiX6qlWL8fGZsdzKm7J7ZdsWU/GB0SKVta2tjMjYIZb234T1UCQYJ2GhmmUmkgdfDSJpwcPl+7
D20ggl9grOKDhSL7d4j/0/oej3BIho1DXEXvS7qrR7TV589ez7XX7bftUICkTaTTjp0GkskppB1g
xiqfKL2yHnXSwbMiJLlfPp/JZyzqsUo13fo2t2nyUnXuAt006+Ux0rOI+sICFI2rnn1Jw71m9laq
TA8nGuFHHjfI7g/KnMwnlPl5I/Ze9CwAFK2ZAQ7G/V5eMyrzCPUU4C2dwznaPfrqwUKFQSz8ysDM
zjSvugFkeM0OtsAQfjKW+bGTzaCXSK8sLWw2d0oy39d6wwtT9mGNPjcTJ6MmTccdiqyVpjOoovdd
dK+nmDDGEjHxCYrNcdYL29Pi4xSsDTxQiC2xyBb13J3IardQCa+ZXykdVmMqKlLJW6qVondYT5/p
NnetGcdH3k87bMpSl0ckl8uV/qgLOsObNNCc5lWd2K1aBRAl89fX+a+HJnvgaihZ5s8ToCgjZ9Mg
SMLOIM+j8uOsT2nW8VfF9X+HojFWWt1Jr3ADMV886mqSztWpRC2rHUTp+BIoVoXK5AtziPoKmlgx
UkudcIcYTjF/qKbaElmziRDXBwzpnnb5mFsvSZ7yNgQ1lk9MSYo620oOoiYBAbKmPdcOQM4r1geU
ke12XyqxvQy6QNKcMJv7UmOm7d605YWirSLv7Vch/dvq2AJlFp20E/Dbiw/1MydZy/ZzqV2+DrS5
dlEZopDDHptTgtjFGC3lIaRZiMt8vPbCLq7KnoxorALdEGUy1KvW1DMIR3PrJnJOuJCZfp83oIVo
MpT1QNuGcuZ5wup9JH/VH7+GgTECV42lyoRbSV7mjHrZnX4wnphIZVVvj8n/sW84ZlDMYQSWGo2P
f51H2kQwc+V1cT1QiOsckFLfwx8GXXn3hmf9oDhSJVf8dYWXmZaTTkzTcKIOV7DJl5bWGcLIAkC+
70w3fn4Aa/z+YV++39Z0byZnJzSOhiViIU/HkneccTgm7nfXYqnCYeIxAXmO/DBrNyBTvj1aGr+X
68UQCTlB75S/8TG4CBA8PeQenntlkOk1XB5VCBxa0as70HKtaFFUK5x9dBf48YMa/gSKlYUW0BWD
xZJS95wnS8kFIxPRCtTp5jziFB5V1xJ18qnSi/c04poSpaMeeKGWRE23WJTSeKhqk+CHlLCGDIbQ
l9XoWhQyIBIBFGseS9A3ESBH8t3w50i1ttkjDXq9pnad6Xnboct2I30TsRcjbZbJBP2tIM2OOr5S
byE8rTQoyiduQM3JM/91q83hIiQX8FvNuK3GiosZ3/cKFZIuAqQsiuWwGl0y9QD6lOCgbpvkfKrR
1uhvMC3QrYf15nzlN31fxWV3DsLJJXLhU0SgDZP0wfAcPNWIi09+R+gpfooeICoiSHNYsRn3nAFg
FaxzPg1sLRHTZbTPL94ywmCuaBxN8Z85ZgvoXY/49pyVQqgtHKRLDcEFCWExEDY81nDnEfM2wkJR
iCIcLfXyjM5j0zol5II9KyS/e3AwZ2IdyHQ2VSH7VlUb/E6PtLUVCBWIoF2EJe/FdEKDl+EOzbpA
1aI+/ufrU/FaI6Lv7xHbYuiDgWugK3P6xHMrzRljFLeJe9sl9kmUw/1zU9R8NJhEsChxAYifbYlh
/LdnQQaHJtGUWna52ea3o7BsY2qSTZvsicIltqOmOmcn1169KrAQrJGpwoyFrKegM9daP1YHBKM6
1cUPfcnqqh1JD52H+l1TOGiiAyfzj6CiYTucy+3EYrnH93Ty4j/7MG8Vf4x+S8rlN+k1vvkp21sI
QyTlIJCZ5GQ7x8Nz3+oPEw4lDV4YOsb805R7+Hs/KoylPZLEC8ekbujJyc9C4xJk9oO+fvQHf9D7
eSivzZAOM6AERJ79B/kBb8Pc8PkvOl2KFRfC4q0tDbBebIn1+Vv6HXcX6WC+2imPCx8nO1nw2uov
cZ81azy7uwf9l8H+YxSQ8szfjIPpL5gqg6c8EfPXfza1KnlwDIrAL9LYfHG0OTeYWmrnbdbLVu2g
7KYR24FYIIphwOp35TRFzNV4UPQ8U067dWzt9rkY1GCg/z9WSmEIBQyNnPt+nbDyXEGzvuh9qq3U
MF/YL44pNJxwnvsligum7UsRusnyStk8xJlysEuIKBurJiZinD1j3snPBMFAa9IG7etkum8tINbx
z13pblEkeylPRwaei5e3ffst5ycdCiBWnCREEs3iZ1XapvUoR1zlxl8wUcrvMT2Adr5obLkhSau0
nV/wo5gmtycCwFvQowbmy5yyZJFvtWqZ9H5Q1OXM3Nux+XB+HOSLMMffRsQSXkyeUKKo/vHLvFIp
eXTz/hj7G/ZqTBnxa47tZfWwl9iXmVWlNWchoqL5rvfcgeLk/8lYky2DkP1EUNq9cQpFVUKc2JyK
3Vw7UmlwoYEjNpKAm1rqJbkEyG7BgjBXF+3X4ezTJvMrK9Gp8xe6nuqhQy3AphISu/m3+15kdHpl
JIg8mjbQu945i66/PYyz91eVkbrTVL5reokmx8czL1EiR+qgvUrDvuTfA0t1DaKjOhZPgZvKb5Mh
stjPQ+eldDqLz9bE9dr5Dn8sYM0u1/SAXIK6qBrEKZ7zDYhtWhs3Xk8YYDAsPnk7AGcPgnIzNJss
B3vfNxzzGUnp6HF6uh6m/u0q6f0GgGpgNucpr/NfL8tXlLCEgQc5wKRhwvRCjfkRLhU2E1dfpV7z
K3gD7lgpG4LSf+D206Jwpt6nZ623QvhuqxpG3I+ZsUiP7Yzryg0nqg2l2WWuWAmeS+Xhmtdapfc2
I6tWtQ6xrpgsoba6wutFS/MSptBepDqlFfxiu0+qsaymmCUD7s5oA+7v/zWRGb4HBqdObsNgw0ZP
qid3eDbtOm5B9kjSOIT6xrcwcuWwss0athpNYlIqEnMrBEonRSb2ZuZCRDbwcU27mwh+2VlDM2z4
Z3gAFyWcWFJCW2zSNdKR6i0pkGLow32q795mmIwy6UuNaK2fD9xc0QwyOk3oiKDtYEWiKSAVpsZQ
bCghcHBPofX82NHGApPIuhx5Wi/g00RqWFxTbkQ1lUeGZPUQpo4uOYKM3GkeNXr9EOcS6rS75fN5
RenN+u3YFaQywhNj6sS52/aVrDc0lBXdD+zGoa8cz0Zor764toAyLG/LbIomW8BkePE5GGHtKFjF
5Xr2flq+F6h7SqJsA66iwsJTf6IlEu+yzIujuRN0lVFDNSyD8l84XbBSIHZJQdbklK1YnnunQUin
0lYVpcOibXMnvNlY3dsdboa83w5G/aROVc67MF0rI8ZHIPnx6zbqP16I7eWKWon9gydg8YnCQ3e0
qnt+6a/RJxpYIlPybJ4d8HVMSpwBf64QdHZUt9uM0ZEzTQl+K36tEk7bdJFM6xePWVFQ/nmNMGIS
ijs3kp0UhRbKEF8UNlhFoLyVyCvDiLruY2luw+cl4i7MJau570Nju+BS2iOWsUNFa2Onaduuvzix
Sep02MBhjWvy5d9qVB8bYupeYXDziTJVX6ROQFHmxLbDnlrps1lqBNjtMYkEF0+3BU9gpTUT9hM1
ldKF3IR+U2sscxrB+bAEzb2LeBZSP4f96QYGkNq5MFIEyHmloM8rY8jnIig0DuyJPz8YHYQU2Fmb
lvQPPRYbc6wFuoxruj3NBvvOs9Ui8g2OpA05YbWutOc8J//0IPdcCpc7LiC0+vFbWgnJiPyH7ZnS
NbpV20gZKZvy7NwPs7EJyFUTZt56F/MXzEEj1pZvJsBmBUqyt6j91/onyzVx/+vhA3j94v4dh/ak
Xo0nHn6pC+Z2LuZvjPbIzRjzATKNR+t2EqBFMll0L3YJ2lkoRWD1vNHq/v9GM78YMsYxD6yez1IU
P8KTas0dEdoukOM0RrVpjJmVLsEqQxITbE3/3zFKt+XnUhAUt7byX+9xTm9x7lkRSidMYnZDvtUT
KQmLlcmiW/jOsz1eXE6GgoWXHn3aCC60ai2TpLh1tiOVWrhn1mWnxKJe4lFZe3QfyEFhtpYnuzKo
a4YH1LJrW7TgTo7AZPeJ1VYFJojWNr54DNoSIzrN/xD2y+mKvykA/E0T5wLZ9OFp45cMBm5mGQli
SdJfUW2YtCslOYPe0HlVV5XOrcGTeSLfV+6yiw6VgbEMnKEW5pdktRgnxncAP/DL4p2Go6VPDLqE
hf97fQFsUrj0q4xoU720wI9+iz4jFqWR7hnAG6/eNvZi1Ujel33UzYue2lx0JsohjFY9nLfY97gJ
vbJY0nlCsoKwYYT0xJRJIoJZKOoOg3EGijY3da4xIwY6hwwWRa/l9X3Qg2XRpMZDRWQwBchVGg7S
qtOIJgs0irGp+91mHloBrxKgD6hBXiLoyFghg6Y/vQow8hFCzDtDJb/mh32qkttlIs2IjH8Ove76
CwMV8Pv9lR9qg4FmF9skmHQXEq3YOj8UEFF7hMTBpjimydYTXfX4NHQNDSUCznGpMoxkJqvHyRdO
PWS4SWU/wFHDtS0pCClzWF2FiqFmNA5kpwM9Em0+mz0JOp9PHhFe4j5bqDNKHHdvxcZq9jBHI12d
ia8YKINg2N4yY5W885tLAQ9ngLvlzaxHIE8n99rUl10P5kc3qfJjfz58Tl1I8Nmyev4cURJuDMWk
U5K6TuVRYPv1g5i97GC9cw8hgRSsYgZtOCY4liqz+bONPKWTJr5Jz+8DllIrx3rqueLWtmCWBwGd
ocpBj0/QTtqVI1BeX+GfbfCSrFtnsG3Xrn5fsXC87P/OBwOzFsdTSLrjakDU9Wi0uGxd4oLcVnv+
XaN0/plr558L8FoAHXIh2m1T9otZ0toMr5QaXOGBNBfzqGlYnbq0+JFjr8XHfbTMeEnEepyyvreg
af7vkwZHnHdwfCS2csyf4X+ASG/7ZscxfanWfD0k2vRpMz+Lo2Pbzoct6jobHfe67oeeUQBp6Mrf
T/yciZjqvt/5vLhVdgwpogo3Z1umvi+QeTD8VWE6sf8ilSu06SgagZMS8dkEOiXIO2idHMldgs+W
J/ZoY/9zOIT/M+R+v/iIj2SJFmGrHWniw6ZXS6009dds2sCNtSX2/wg3g0FatQfqFsNC9+9ymT39
4qURlL84BGlVI1ZSiLfKohoZvA2N3y8M6k3box+cfdH3FNubqpnY4xFNEv5PnhaOjnG/BVd4mQs1
nFA2DIwqpeIYY7t0wtxKp2ydV3MYF518EzjxV60/dXBJ/NnfjaOB9l0dcVRj392DuQZQ5KyXcy0c
JZpydi6DEST18NGOJdPNAOQxYacTcJIOosedDCWmbkuDrNg/4NLDvhwnneDRiWPvN0ZPFNCPDFAA
Mat12dRoAmsL3zv8brYeIOtdZyC69ukfer+tHODkEYdud8+l36KS49cZkLUqrs3vwc8ZPSzJTD0V
lTsqLTtl6bNO55uCy8phGnXSVzgAHZ/fEZg6pqxP1x2BJhbx3XgO14wjcLWnMVUH5E2c4yPi9a88
6PSqFN9t8w13wfENAKA4sWHZVrPXkYaQWqcGcriLn9msAYGgYiNp7f1bhHrTICn+SRxBN8zFLsqz
bLOh/bIGCbnVno7jKNuXM8ASCWfj5gpgaG02gQzhVK97/p7cqiz4Jd2PO2z0qi9eJaiIELqzuvkn
Yk2XjzdNBdFgQUb/oSZBGNdmTiN53B7iH9b8Y7an6XrVAC5yWwMRxN7H0mazZ+HmXHVUQBIm/8kq
rfMfdP66tc2eC+HeDqWYvmrcwEkI2NlM3NW6lXjWhIuhhsHZq0CF2JrWbKBR/2Q2s71NY9FJ89iL
Cd0qQy0L6DAaRkfociXjP1t00DoCL6wv+jO4RvORf3B8iHNAq5K5zjmM6Sf5ktnzN41so8jbq55G
Ze0MelDLNZjslujC7YudwB+YuuBO26/SS6dQjevDe3K2wmP/ENeu8A8JYq9iW4eJVDv0TfFZAEPv
PGcB+lhdw1IzKcs1QvTIswxRpBkaEEZ56Vtp9ronGDu8pBB/7DtY0MNeaBi/+0wR7+VkcJv2UgT4
4g3CJ4m7Dp0nxd2Qkpu9sm1Y7WM3WYX9kan7swpTtf8BSX/DTrM0f/di74PJ+AYHzuOa0YydGU5N
9Gx+v3Ihqrh5tXN74eh4cQ6ETKcO4mrtb0er3mH3IR1kh/DTylk7dgjR1n80JtLzVcsX1Vhb+hdT
8guQvcJZUh34fqLpbRjJgSPhp4ubd83l4dWg/RUo2F/O5QpkZDA1zunCHoorebF6TgzzWsqpcqvf
5WEgI/WsWhz01U8Z3hCBTx9R/jtVtJKvag32BKNi54Q39MOa9zPzh9Y8RIaKAlW7Ffj1RKw2qY02
KS5w+G+8wAJuYuAuRsUnJo2LZNiTpzQr7yBuDKCa63OvxmXNi47hrDx9Rg4euSC+RzjEzQoZMhG8
1OD/Md+0gkC1toWwFuvLeS97k+LYnO+ltK00xI+287xc31OomW1BYtQIlI5OqRT8aQJeUxBYiTtJ
5YQf6QbidO+I8ad25ciCFo7uIp79WrYX5VP//IBg2YVZLbhtzkHyn6qa708kl7++9QhfB2tcq+eu
XyHzR2LA9zP+H3jFoDfEEzNrChxjTzP7T7OAonsqbMALiCws+TU+Rae49ZLCCFg4CkRzPp2AryEj
OAdaS2lWZF5LU0+fv8YIM41AsGQHKRz3XlPMtD6a4I/FgLIFPMox9YyO1YQj4nD3RDpdg6ZuRjcw
kCONbR7u0cyfKezVLVuBHFrbGnHYFvdA35TEN96dpwU9SQmPXs1cuX8AqjqT6qFEa+XwEIg/srpw
GEhc92VPyxiMn5TPUoBJOf2rRayDGByhx9ltVEbSwKZOdp2xahsFjaBiyVZxry/FdiPkpPVImxNt
+YSEus/ioe+zF2oo5P7DB+bsLg6oo5YtkGKvX5gSqou4G5V8u4/q9AWLwUFaxIG0Pw0PRVJSHlAn
eDMOLyQB+IZvRmwI4Yb0HnA18S/VYdDpJGdS+wtAU8ACSVr4CDfzBVCyRGcavz4x098d0C6xxuP8
80vaZoGUx90LaDHNyWsLHIzsqA3RXIE68driqzFGOM4nL5M9qlboiFd8OX6d/gJMPckcVaGTgJsT
vDBEKoyZFkq1u03LnPUCYHU9jT8DtoBXRdNWF2J0h6dy54vtBq1oh0RcucJFeUcrghNxvwA6tomI
c3+vCAR3lBKGAN44VJTMbazLwVyG5VVEbWqx5MwywfMqfsfCjDjvB95mR8V3kWLKXDfoarGbtIOb
Prswljg8vM9TbO0t0d/Ya4vDRlA9rt8H/l4lNmSPTZCMg6ay9hQrzohouWHMtsU9pZFndZ+y48WH
u1vQu+Y8g8FL9Acw+4ci1b8WL5BqKF8YwEPbXuJLgHXag2DJ7STVHjUvRR+rNezF8n7H1W+i5CX4
F3aepaUsWl65uHjSFRDpRs4PDECftxr9ihm4nLSkKp1r+wlIctJ4V4FO1F/XbMY2veXbrJ9sFKGY
RpCWnxx1A+l9GJO6Un9vIgxThh29Q+y4zF8ZlryzvBNaFaLXJ7EJ2uOTtFLPsw42UB6ZmC/VF8sV
0v9UaC5zdNcaeA4xgiqfy/Tj/hMJljotQ1SUTKTG9fUZmRog0+o/YdEGZ2TH+ngwsBxBYfCRCW5n
0t5MTyQSSI2olA4aCJMsc7fAVidt3uRBpdmWr75ZJo9fyly2dB8auWT19ZpfthMAvDj4WzHZwjiH
avWmvwopoKKa0YDuLhKtoM35sRA3P8ieWEZtr19JsCawkRJqug17JwtucOqvcalGdCTuydjZ9Byv
Eu3GhEyE0wmIlirFGCUgC3cjYZ1+LJgEmSfIeuFosnHJlaN4ZObKCjRwr6qZuHSRAOkg56mP7Jb6
jqoV3xmI5Zwy34fM2R6iNbouWZmy40XKo/4Kl04zYPEpOgR5Ld8aaM7TCWelZkUKbnRgIfnLzbgu
Y4qYCtmEPHX5gNWg7cfCX6Co7Db72jorm88rVeor8VX0n3dsp6g8Z9XSQUA9/KlVvXHhylcsOTFy
sUrmj1YECQl2J7IW8SF/T76cLSJEMcmmEDJQzRQPGlvHYyiv7UsyEXZp1PHiYxNenGt3Ju5jLFF8
/MUUAHm32nW4HD7Ewpzg4MBSZLpCKSGV1B+MSHI05MhGUwLmxMuAGzhq8fnp6+bb0xq1LpAX+M3o
dI8i6uy/qKPuQEt9zJWTJ2XmK+zwsQLbZKrhv1CB/2MSvQAamW6raD6FsgMFjHvQHAkVFsWmUHRa
nNQxjDrPfmLj1t9MHI2WXrkPmmHeQVHg246/MgYYsStyqaLLnQOWp/WpqiiEY5XdrJxLL0z2kaDC
SRoudtRoy1IjNZsHZwTGbyF0Eg9xSAxc/uVMpp1FchqXb8MefoQS7fBizP8oZRU09MSoJ1R5uh6Y
Qcn1I5KqKq/I4uthc+9hd9ZNm+8FWCth2FfWQIzb3OqxgNIhvPqSeBVzOOlewtqppQhQrejiXchZ
/cyPHsbktTz+ROAN22nHSEqtZVpzHLvOwapOvlSjQqx2a1MGzbXG+EeoUn4H2oUuO9T1PeduzYDa
hCrsWbuxcyRGB/WQfPG1ec/ELIMlJlOj25L2uPXkayP4REza7pkM1uOTegu9p4sdckgkdqhd+XOT
IScOF5tz5SJ7bzJc/XACQTFLoBdsddnjBkO3i4L62LppxWQajQM/9PSXicahaHzZw/nYyOhgaZcN
zTcEARnWRAahdfN+Q1Q+Yb/N3b0tLuYcwHcGdsfQmWWqCN/QM6pxMXJ+szBP1Jr2PUyX6kPUVgvx
QrWvR8wXpaylA4bcL6Y3o8DuWufyHDnMuAq3yuIQS71SzDhyWUvBNsAIst3Y+DIh7i+MBMV74Aqs
lpLw4K5xcf5s8YVgB2BnB42WoL0KU4Tu44RF/ZxR3SLKTgP33sKWKnqaZtoSqEj8YunXqdfeDNB1
bxOTvftP44Lrop24zVJXmCCSuRAiNzBSBiFs+FhrEzUQih2g6/NLNEJib3LI8u/VzMOUXmtlRxoa
82wG+si8eFDa1RBK/1ejLAUy3+2dPNnDv0cSDTzZpW6vYqL01HqAI5TM8rbRI0/O78IF+OBUJA46
EQMC16l0M9eATkCOXhhkVi7r/NzFkDkmtAd4+eU3Z5poocYfCBT11TeUTNymv/jhQjTlTaswTjp2
YJNTNWFCtkZ8tDZ5nG0t6btY63oXEp1KrBG06a1PNQ5Yqa5LtxUnrysJEvA1b8L+FfWAdyxZK6xb
W+PAcfTCyLqqStfjzkqXZJkZUYjWOVxCEZr9ce2x9BZ3PHS37VcstZi4a8TE5XEq3BlpfurZLLpf
a/ABf1uuQpO40y+BuSHk08gZEz5v1/gnQ8hHSrIvUsf35tirNGoE/0qQrtlm/OddYJTiRfjrc568
3SwUF5AP4B0no+2ch/JHKUZmOWD2TL3lFCloMBK+BjLWtyTe0z9zhlPv9DOd8Fzn7+4tutggNprr
yKaaUSB0hafNAEF+tIPdCooF2YFLvkQb6M/aLKgEZYwvQjk1JdIdYV7jIdZIwDAwVE342si6y45n
RDBejOsKL5uJU/m1gwEcbbeI5vSbg/b3vfa0IJjg4zC1ecXuP6XzCLI9rB+FRxkPKMppiHNf2v94
0hWFb3b9qDOGQJkelfF9eBN0B/7e7f6HSDZJf8N9g2qE8Hty0OSeeIyKs7h4FKxqhHT5T8xBARTg
TtEe6v93L2R5rTqZ51HGh67awRLQK8HRFuULZm0fmzyAQghMKt1mek9nw13tZ7cwfHwEV1//XJKG
us8rX8CLJtymhOlxNz9H7guBSuEj1a2lO/fGXMp+PV3ex4uRTDTLrZ1K4OMPasT90WHcraWbv9sP
iEHaRID3rQraJ+FHQ3Bketigo+VFnOylulZIEGbaOsBOWZcl1cucnrgIWJpin6RJXZ0OxzldUJVM
18hQJqYugwypncnAhQF3NkieOCU7S8lyHezIrWyz3fW9kTIcVtNoArKkKE7P0UXSeOWXjTN8SI5h
AOLGjhIlLMo8vgsxdNE5n/U+ft4WSVKo9pG+8bOTvhzfKs+GWP9Rld3N6LeAOC/ig8lZ+4OIT6gq
qPgBxkYVKwA8nGIGuG9ytm5y/zf1+KLCwM5LIEgnwVCGpoaqtO24nANJgXyc55s2dIvNPgnPmVEC
tgaIAjwKAzl7fFjZQmmRkXlrEjX1KFwaqfj+wHqPDAZRUe4FKk5Gzzmrya8mcAEHsU1yV0OExbrX
z2zhLpTG19Z48jBmRUDsXeI4cxEPbwqKv1zbthqAX4wXCBWk1Qr0uFswlFazzVAF7IMdVwCSAIb9
N7f4wdneOV69AkndaQXhJBvOoRxfVQlyR2i8LHpoyzfp+0G84O6LBZiX4RxMK4IWp7RRB0Af4GOF
upWHI57OmJik09SQOmyMofEt9dHvcCYXSTzOi0NkxtH5QmWeRXCz9Wox/r857OD2f118Pe8+7Drd
6lJ7Pq+7sW620vlU5IndBsZhu92/1cErdBj5k2Lma8FARwIcGWluUBmK4OPUT64c7IN4eM1Utp0U
vjwznP7DhZ5c7fIdUIcKaPBNf44vyIK2Fdop/gtWY29/JLIkvGmR2Qk3aAShwtlDA2bGkQMl/sd5
pqmi3xgESdc2dCw+Dl8s03NkgXp+coQlXq7EC0z8016eLqr4itMROfqjqdn7nbejr/AiWqYt32zz
nxOUt65zX7dSuLLQmd1GggH8m998OchYiBz1kke8XtrY4vBDnpki1yLC7RlQjRzhgfcY9/aBoM81
DBGzZ6tOyVDCg+UKFN28sdVilk1b7bYf+7nYQwFkbNh+0Cm9qOgXF+QxCJXSkpd3aIvjdzKWcE1F
0OKIxE01pihkDI4gZc+5ttfp4FpDJcfvfYUq+Dyc4v0YZP00K2PiQew26E7s3HuoLTAY99aQpv3v
lpRMBFjlRPBwPXO7J0VJ4y3rXYxYmEwUiloaYi/BoE3GCWYSRP2gU/vsFBexnpHJNwOJ8tLJ8Axs
EN/GR0cS2DHubEYAPWr21hNR7u67vCU2cXwgsFZCuSiM3P/LMPCMP87sbGioSQ2qehXn2+kcMVjG
0B2EHmeZTNBsW75XrEzPSGilp0u0IXi/xKU2nBvjoM1qBlNimE0h3fb4ctOJ2I2nwfhmFO4hW+2E
dEv70yltBuHtCE2sOV/0AV48dYWwEf4ZwkFrt4dvOqilH/dauoWTHNk26HFDbZtRZLyUschImtJc
PEgeWSgaO3GJjJC2L18Aeb0w5xDmQJNe5GY15ymGSYdP5BdXc3I7BFE3zO0AYyUXRAmdUNTqcAT0
AmhxIOn5qDTCbh47WN1L8D49FyomuHfkxIZOOzzz1690/wAah7QFs+xYK7o6flU19sIfsxhOCTiF
JOV19AHuzqrN3OxEHGwm/VRi7/98NAO5yvLhhxQ1ePx2H6ORPuVmCbCfX+U/622BwZOwvSLe1m1K
eJDF+HV/5J47yY/r6xonSiAkxNyZvyvK6uBjO9eSZL4AbnEHGgu4K+//XaZGiwoqvhuaN3Z4uR63
1pSEYcJO6za1gOflxymPhZbF4TbQ1h7v/th1WplAAtoKHqva2Erf3WaZ6BZyIQVxwcHgETuySoNr
ikKiAO0fs+AUDo4Y7EQuKDsFRlsUw0T6VjRVnWDrzCCc6VYZsK34XMg2f6mzEVvgKXBDDhXpKsDb
RqmCFFzCYQWWlqzYrnZWI8GsbvMh5j9GtTo7c/MFLcoSzoYq0RSV3xPnxVQbXgzNpEnaw307OqhL
QyfU4XcPXIH+rjq9o53VA6Yh9v/hTVFcxq02sfkrRPLQ4FLUhIDS3k2vm0MokVNkHoCyLTpGhjb+
ekau/qgadwp7Q5NQPJ5m4hUPHcTp+f4Kz7YyQTxPAKDqNhsYSLw6mABAVANnuGpYiPXDVYHvJvHy
mAST46Rt7qk6opcDASHt4qu3OiPNfooVYr0DQaSl/CRv6D1hXnRRQL15yBL1UnpZmS/KviJeExMn
T6j0ZukFxTxk7rVbIisoLm4CV1JDfadLbL3kaTOC0OjME0SFOmf99NSgCNBkdEGlJwnNcsK272oO
TD8FZYOgHlNdA4DFP7/zoReY2xhfJ0XWSnN7yIAo0aBLyA9fdm8jP8avfYrJEnQlAznVPYJ5a4iA
mpCE3k35n5NYV6/qnGLvXu9k0eWInTNiOHc9hnNduyS8yzeV0Sy/A8DFYbVKMKh56bkaLoWV9MuM
KeZvt0Vs9x+mSdCJMlXkLPuhsLeGRYcjB2MTJYHnqTMFYwlkfaodTTDjhFAJSShTqJcsBuX5IPdz
G45GIVEJRon6YqW9ytyiCpCaJSUXqymqPDlBkZSoHQI9pVZ+MTzwsD2DB0Q2hPpB9opmNk+hHg7l
V+XzCEj3Y1qE4J6AdJioIOAu3ixQZYYpy6RYnLqVijJCODJFL1uIjbFhdFRjrhODvGXlNAst534l
wv0RoCquL5KrXPnF2yyDfGQdkaWbp5H4eeUu/AFtWYgyBmB8KKiqODJZGkGr66C6vPMIhUDtIPVK
2VZPWkca4OOzrkKTK5VOQJaIhRRq2FrqvF1xLLnRRIWTyDV0kQ4xbTR/Op+ubnC3knTERgbKy777
O7kZ11SJDplrZ4Soi1EGVkTmpD5GB0lY9ErP+y0uTidpCB1KIsoqKggdtwQLzVZ5+y84dSsRCmT0
VdSppGev3OPJqr4TFV92/8VVxl92TINOWFUSBn+lgSfUcZlqe6RDOvPlUpfBStqgRCzTjx5ln2uT
W/xqfKCvic+RvQIZXzp0uoun4PSAoQpcJUqeQij+cRIPNjZPzKX88FAjIeqlBtEmU+Ar5+5FkSoh
qMWmxaPeHQWR+opsQPFJLOVcq1H00RgWHibtD58E+Dv0Emjmdx1M3q4NOPxYgyhFGW49RhjzdclX
sSveUxBddxDPt8HUD1Y1Gc7xOgr7M4AXVa+fBdzf55IgUnYDeNpFnegw9RLvNCeLZbzTlYfTmN3y
jdlArOq2gEWIHSpK6jo+rR4VjQ8vW5+B9KLixklsZ9uzcu0QDRYa5jCL0SVZhdvwwnlIz8fYaUFw
JDXJ5dP4kkK4wt5/MGNIuSVCeYxDI++tfiVS5+rngrnw5jZ1c50yioKle+cwnvCvlzAf7hwDYtiz
PFnXtjq5OamwtOtlv9wl9MdcWeaCJ8HN+5U5yErpfwMLL+0OsFXATf07zpxp89L8j8CUwePFMm/8
iPcf3RfSR2+y3pKEYYeAOJjpGdT1SeiHubaNcW2LiEWt7C4WpRbBgvkMEO3jyISWGSDn97FEsbGg
HAkbDVmtJXjh2fDDNfeJQmpMFDPfY79S7X0cPE7ZxkuI4vgqmNuKKnXg0IJ/BLhuAABLruENKPbW
5ouKem4ujQIspb8grtPhRdAqtUX9ZryslJ5PPNkZD1zRLd5azFq6fgHAfJJLNlbOz0C2OvkFpm9g
cFTX25wCzi2yOQvlyR6Q+2n6OFwhYVWo85NhkZFi0GrqWizsLzKKIqxmvM32f6gcwX9Usc1nB3dP
fG70s5DFbwvdkJ6eMGhl8Asg721Cmw0NzwQBuaGd0vE1HdrEs4EZWYHze1AafJ+n1cdtAd/73tvv
fmjmf0Ls7Gi72roRdvuyuPcY3qr0gIWj2DugNNnVRubC7DJrgOPgt/ZIR2d8NgXS/ify417ugblq
sUodoh8Iaf8m2wWrQD5OMtscm1BKJdze0AJRQNZjVKPNVJimA3FrVlN8m8D/uz7YpjMSpESofQph
p7v82wGjwG4blirbSUdADoxV5lnthOfceODAgoL5NLJ0qdP9UZBJJRBEN/m4A3csk+P6KfjgPPg2
KmbmXgVcLrGfNwh/1cSCbfizJ/Zr6OS6cZnlWh4Uzllg5t1DSbuNwAR2ebx59qSrunwmYzFXHQDw
8k0CdxOQEs/PARnsdz0fogGWScJ83uBErmb5jxIpmbrUsp/BR8Qir5PDjQ6C0wOL7wCCETbBI2rA
3/s9EiRKfR65Wq9fWroJaBHJXL38xcIZbeIScEa4qLXu1R2e0pUIrkMRkDNhKZzXVwd+T8kAGmFo
zFos1sKgTuE2mlpuuoUmfBMv3iOWIu9kHxPrRi+UxtWOwoi7FdbaBwxu0lY6J/VlQXCCvWZTtBZX
EwznPquwmKT47FplgqazqSra02JlxJerANVo6w3nOIqbntiFuxvgp6fs5K8g9BFGbWO1XA1fLqj/
n1hu6xRGnN214Eb8e/1cyQHvP399LOyhM3G6EKecblplhTYkTcfVC2V9BVCTg+jaIqfGaRlYEEhm
uGsnDCQEuZTZfti/G6imoefG1Q4FnK6v00qsyTbqK5B4pCw8OdS/lD7VjaiS9Z6rCYo4i6BkPZEv
Jd1VQZ2b4fu9jCkf0xoF5VI5KKgQetpmweMI0fNM/DnPcfr6+nkERlRK/R6F3K21StB0ahHs4WUC
vtsQ0lmyAqpFh72+pwHisdK09Vht/K2nVNcXARP3kppKQvBpnOUA4VDMmDFVZQGX/qk61aIZt7Yu
v2ae1BIBeclV4C9FCHlV3uTo7DEnzUBTBfQmsgskyax8hEeWNL777IBnolQlRonSD/IaA2qHl6tm
XiSEZ5DzymexvFp3XJphVyFgnShSkMckPNomOWUAvFeJwZUWaivmAMjHoYd/aC/JVVI90eO1jSNw
h28W20Gn6EJzIuaMoQGrAZdmAdnKeqlfgBRQ5oDdjME5mBfTnw+lzhxJl6hojpaHtYTVwRQZzzYu
i1M6H5g2m0IbKOfCqVmoBfs57csifD4O45Ryyqv92eHiqYsnYi/b/rQncYQyEkHePmEecoYs/ayW
tofqwJ2aNwEh0rWoNAF6ndCXsC6PBQqOHWJINVEnAlFlSfaqiSyh5X5C1JgEbd0NCfBnUwE3uPp6
35PAbUrA7nvzBXIB6fSTPiPDdT7Xg+UW57aO5cwJ5Yh2gKImqBg/DgKQ1kezrMVcilQaAnOMNTVz
hDHMZkZHUxKltLbE+xCX2W+GuL0vn7olzd3H6de8PNNUwpDVu3Kh11KHPEU7AuASa97rluuWbzZ2
0fRCmflMwglbNklE+ba5r8UO7TdLlM/ZLW+uTbxQZjX0BFp//ZET0KP5zYMz3qgkvY9Vl6qVshFs
bh1Qw6NSQhe98lIqB7tiCATD194+Nv54o6qrONLQm1uUZnTxbT1WVrvXpQZEBAkTsVrnifdSvekq
8Lbt/JM5XCg6dclzvJt4vjodWpRK66F85j2FLK6zBvpJiDRlJi2/P0hOruu8nGQAQoojBLDpd61w
QNen4iiKXeQ/p6/x21hKRFd0FSCkgtM0bhV2A74xMA3tHTwQkpBLFwQUvwsMdKRzIjI1vMPlZ54y
Nlt+vgKSiY8JbMyjKpK66nsx9lk62MqfIdjHKx8QLSk47p1Fiv/aASzjSPEwp/xihm2DQvepXWLR
kzPFno8D0T5vdLuZ1JmlSR5XlLTQkmepeujYAlaMmvhR5r+e5Rp7JI/ccNuUK2VHiH269jqTCOjs
mx9mPDaxPWgg1iZnd7BOs0iwUcRRwNOyH70C+4oUXlkS8YZshv1WmOAU6iXQTvWOp9ZeBT1NoVoc
TqlCy7HrgU/9ZiznvXpF4FJKuqOVk77l4p6+Vwc4kHDeWth4DI8BJCHvE5f907zwtd694HjB0zR2
Sb62+XLSZs/qnBcFUsMonIPYfC87/Qr1dex/xSEgmu0hZrFHsLJ1CcfqIrmYbELvfQ9ajGp4yPgh
oT7UIv6ekxBdQ4thCuTHmee8rIGI/hbAK9+mInKrz6NCGceoJSnVFN4N44K2kwESyJVosNa8sRne
+EntM/JR5SiMwr8dAzEGjwRyxcwWfeJ5gTsUsNKPhlseusbaXWxNjSi80E2w1hxNpiWQlmKNwjIb
i0PwD3uLJhuCpg/5xQOewXdVFAwo655eOKOhveGqz30NeKFCFUwPMIoIZ0dc2fMKOUFWI5Lg6H/Y
4aRnWpefiMJvqd7re9SXafn/tH5gZV5fNvGzxZTiQbbP9VZ7Uchhjqyqh9xLEJTHItHqARMk6+ZE
ZQWPuW88K1WaosBE4/MgE6ED2L0RrVVfP5osISq/De2ia1xFj/rDZNvgl0HLSGtdPK5VzkOoEoRv
BfUWerJyYJTgWmrwpOz4ySaAnfYIrbZSQMJhz7iSkThuCMplg55MU1Ily5sEE4Jc025r7PyR5pEm
5b/7LnYX2bvXGb1ciohbXBOj0ppOzecgUDjXAZkVaquwkNRgtHXoGd2AymXZkKlHPtmcdszk3dBb
J1NS+XbgF0ykmZyTvwuzUq2GjgXn5LPTDjlb05gBcNZf3Fr2yo8OGb64EBkIeYcw/rnBpbk7FHON
gq5mynBAxTeqY2CfMW2vdiI+GbTVnbOTVrgHRosTMvwF6xpRyUV8vQFoczHJAZKjRQ4wHP9d01ir
nrpSxhlfL1us6/mpIQVyKzaDSQvnhyTvLNa5aJNun3yDesnZKhhVmEe+kB/xYsXn20G2TICA7IO+
IMsthqnOYgy4Ghtf9fHGvo5+Q/qQuofcA3OuAgogfV+1c4xc4KbvYslvw3VcQ7UPteMNjGJcJ0Eg
k60KMLo/sAkkCq/G2JSMPJqlAE3ueMvE1WfYWy1HxlSm1mPBvasEardndJv/dpYX5D0AO9NmED4Q
0Wu19g8tfbozTupQjlbAEvPf/clKMtkvZXt8ifZd7RD/qJP2ISj8JTRsjtQdyibcCSS9jWT+ZZFr
7KLlhgDpnrqhOLjFbbxtuLWzwbzh9NDBvxUwKJwAjCHgAUSp8CgUGsG5emp14uwWBdLvoM4iKmPn
vqxIUVZYAqNiAXdcZRPNFITz0CkfqjS6BxE+jrFVCN8xbpodgO8ZkwwJvgCSC0U42ngNB229wPk6
PUx54E/FK06mX8g7U7xoQHztYwMBLFt/WDh0Ic35f4Y7po4Po54M66sDs66HjCQdvWgENsx8yi2y
ciBsr6XGxyA5Dq8Kn+9Yd2Q4i+52kHbI669QfQJjERFwe7WkTl5Cf28VoNvBV62qj5CeUgEarGvP
Nb0TziJDsT+/jdUwaqaGvHLClqwHoxpyb9KIwuVX0+ncJ4OIsKhwmjG9afqsY8vc2T/tJLY+fyQy
PvL0UIV6STn1d8eYVPhOR/ieTXap+6hMQ71rZ1eaEeeeSFX0x/0iw6INp1c171iIXzO4vmL2Ao2K
DJKfMR5++93zrFZBl7NEvgqJn8BQ7QMy32z7NCGotKPtG+9tpX012qm5dOfbsU5H6Oj6/ud8jUrE
gxFKEbzZu254Glc8v6TuJc9vjhb6GHYrt0WLGYg7DeBcoMb+QNtJPVqB6rhN6C+tcHPxHGUWlJTB
uRkbAI8Eq+LjV/mV3/EN8Bqhbeb+0ZSn3ng5EMzZvM8MIBY9lDyJXZ+f/y68t86pBqJWAN09+ckU
iBL9zaHIJSQ9Z8QzA+hsTB7SGDOWpVU0C3YQvtFjYOr9qQMnhtDkCLvt6xufFy6pcZMWQVVZPYYp
iBBt525D0pTFjDhWq/0m82v4U3VJGIzJ+TMvGlnCzvgn0R2l6Gc+Dgx/MigkYYyLUaKMQ482CII1
9T3YHYhZq0ys8eQ6Q2uf+3mNAUMrO4l8zBbvMUpkLDKzBcN4NThPcQbd4MvPYquJMmk6VtOASJjy
WEvnWGNARl+V5dD2sBUDJvORvaQkCQMRIyP+9zpL6IL9Q3vJB+0Z+KJHV9yKa1b318DB/rjV+fMR
zNOG4kx/kFISFpzE0Vma0W3aQa3M5VD3EVbIBsB2AlBmUdRpyKoRXVzagEc00VkL5WSInJeN54jA
fNTs6JZ1FSgmwRIyhIbmQmP+5iIjEfdLZRRX3VOmf7Ar4JfuvU+ObmqKra5ic/2lNQbFxKzEtjdi
fgyQYNzzyd6U1PxlX95AgVk+fNaAXyW5QJ/RCqmBN31FG3zZSjH2WeVKqFaGKaP0RAxPBzL6gQvz
+bzkwTk25CFQqbVea70KM5XxsEXDMCFh7YETm06umJqcF7AmXmGu284ee6Fh/m4tdwXSTOEfEhSH
/uT8goRK/onyU80E2RE4nhwEcwvDegKBbf2Fjy98CfYb+G2RFz6Tbf6ONNoKZ9e4rnLVfUZU2IxK
gDs1JYPudKSw+bpUB4vEjYDbUulg8ZMpNIK7weAoSyU+X1MlZz0W64Q64vzgl3ULbxU0CysDEmbg
hiM99Md5zBFFMFc9IncOlr7qc8+4+efUJnyuD8rM/fC+tsKETrSeDr5DoWCeRY2JivpYmdSBW5Sp
ESH1RLUa8xQSmgVTdneWwAY0Hm3uFl1pIPyS2XE4L8ebjK71U0A9EiHScB/KS/k+h2a4z+7JHhat
XN2zbAtdxPHUgIasP1EBcEgothh4hfKbRKQWP55YsfO8Ta2/zqYvQsDCN7zFoYFlkZ1CgFMOfj0W
miRslPjTXn7qeHI7sidWv63uwGXRAChpjtdC7HxUCogRjHKr5Ckvg5xJtC2CHkaQSoDQNaS/xye6
n72TOPwfXRhh18Ic3R0pPmFTe9fy4p4QyvrvHZwImCg7tezpd/z4X9gq28g+MLCL/NG8dGldhkpw
H2QCK343KVGcri2xa3+WY9b5G9lL8M7RZNlR7s1SM6Qe/sMkfao1wGNda+o5UNcabbvMoFy7ONs0
UYW28kYLWBDxXnldb67AvNSCS7iuvlyJGzA4/wYhLj2t+k36ifTPuuu+dIpSAMNOuoBlUyTLobUc
K9XCo8T2SrkjSpd6mhKo8oBFaC857A8H2/8wSD3vBROFdxV1fjv8JkerfajUKLcB2pK0gPBKDvVu
YnD+3Jpv/709H14UTwcHxF1XzaXsBfvWV8sxaFNUHZ7Gugvmh2o1Li/uJF1W66e1lpVHOuqcwSe6
VnYuTDbfkNfT9vzHrC1cjBIivJV9RFyyBWPFcVEg8UcMaJvQZE7UIdVplvvZ4PMhBnWwIcLFIwtz
HQGKbwscOcWiSLKqq4v0yTheCI4ardRFs+Fbb7Rn1X+xXnQnKkJrBRs2oPo1uWkCjWSoz/0pOV1k
oeunpb6JHVAlRW/JScILKvyD4mz6RTW0H/YdAAXNRfJh1egdo3sHsASLK54+Z9BMYAkhF/9XhEfx
I9KGzpF4EpV0HcBVbqwdoUMVviXrZ3yiLG4YVkQVEezgtN9g/3lGUFVr/+aMyxZLfqmb1HqZQuyz
KcCIST9os9kaPP6qItfp5Us8DZP+xgPNOCPQq7lcIFBlA6AzNirUmIxWYsk7AYSU2gpta1wOGUax
cXadnYU+ySuWknT2Frg2gYFN2XSLczUj85lf9IsLlHzccNlYqFbk0uaRT9M8JXzFV94Ls642aDhK
42VUd3Pt2+4zZ3Pz8aOLPQozLswfUkMt1iOSBk/70ryZoJXDheaSxK/ezMvLUSIcyXnOla+QEeGe
u0WdBOwYoyS8x1aV5/iBhFpEOBAvxCl33HfJjq/R9UBWwPuTAIsOHnB0UQHj4HFBKuecnxOF6owA
/96UvO3O86sa9tFF9AcFaTAhd96yLfDyfIawrVWmr+eXMpTCt8vp8Egm0Dxtkgz/3VdU0A6bOkWg
LrVgM0qBtq1r93Q5pVIliA45/lShvtKAVupGh0y1dQfODQjliK30qAAbufF7yS0nyFAaH7djMS8D
3NrH0D2i35Vmf3ewe9Q/CAi4lK0AsScq1/vCVEVUWb3px/JeEO3IG+Gv0eli5NyKF2ryy01Djlst
8/jdbL4SGjAUOkUz0U3y0wEd5LA4DdQd4whbmPUX2eSqiHlXrEiDeRh99Mkn3nSwymE2gmgtCNEN
SvvMmAw0Gnk1LmrBLebOQPOCcf1Duph0uap1oAezLO68qmFVU4+QEWdmYgvuIkfSGtPAKSdq+2IN
XqWgkTWZdT1X+7IXh4HiughWgz+xKzmK1Ly5crxg7gubu8gKghZVbVhVJxAQgQwtjIhRWful51ug
IDhidqUIqI7Q4yJdG7ZfPgwGm6slFBaulGDaRPT6lCB2XsPKg8SRkHLaYdUe9F/x0P+VjGHvxAKm
wF94j1FuP3s5uVBxluqMRqSXqpqKl9B1mn2uEdO1Yg9zjgDKQ7SjhO6r8VOMr3X2LR3ooADD4Kv+
r9QOxxlYMOPbnxtNmfF+xcj4Hv3hQO0WVqgVfBOW109qmFay/Wb4VRpVikZ8kIrG9Gxi7amm/Xh/
cwzbZeP9mki4mw7EYRTHM5wzL7FfDRr+ProQ5ZsLNh80rJdEFxSSUezREPSCcRfCUdAUnUsnML2q
nyh/z0cx/Ve7N6W98kez2ozLrRgjg1exnk0o8hREv+ZSuzXsF5rCc22iiZs7GRvJ1bK12dWMciWU
iPqU21kpoHW32pzBgft26jMu3p93s2hsL+fMc/UmPyokSEssF8f9PrJoFhIF9sfCE+PkfKmtBYL9
qNuZB/MzVOGKvOj/roMe/jQaZ1L643OdyT89PL8By08rDVtH3skeEAZc/SZ8swp3PI8u131XLiSi
0TPWMt3kPbYA5oough7CK0sATPJuKLYPH65OOg5bVF+w6HwNMCQ6nCtgx4KQeFlj1W+NnfuEXEB0
0n7WAmem0cckOmmAXfdiO/qX7DE8kSzAoh9PiIwp771gcZdHHuf0mTXa7d46jhJHMXZb1RIsRjso
WMhambLoNW2tcS3hY5oFJ1MtjHiwllGZX2wG79OqKgNyUrGe145oW8KgyQuAuC3OMVfCgErZnov5
RML/nYjLJpZ343S+ChKOdbGL1BLZlG74J0PIbgZlkUw12GJSR6GlgFzPwD9jCIfS4e8L+LmHOFL8
bH4IYILPMB1KX4WOR5cFYqUGxy9mBpS94X236P+2rEJyJzkzvczW/c13GoZ7gms0BUJHUOevnrrD
64FNufKem9ncho8KckMckPINAi6zfTd9Qf+sgwj09XHB3uZ2i3vZK8N6O6Zk5Xgp6W5hvBexg8aY
6QrC/vcAW9rzES08Guf7hOfmUC6P6jYBk8unK64GmQn4+xo5X9pRNkVpX0sgCgi0YsyaS+hqYb42
d6ebEm/JSX76GT7fj8sU6MqZalllxyDOqdse5vpulUqcEeDAK1tFD/tdNfyXOSvVro+KWu9FhqJD
mQga1VRvjYtq0LHEgZ98yuYL4aJtLT5rDu97bDqXRVlytoLSHVZQBxCoa55Uc62AH4WRccrXaGea
UFbmkdGBRcV6NZxmVoc7jS2ZZWGzKzzRSL0tp0b+CuPPNFpPW1TV1bYeKYRF49FGzSdSzdF2d2Pm
UUMjqRALtvk4a0iT33OlTwgS0eaKdt3G1m1RF2DLjw81mB6RT8h2z8f20CEbkZIxYrsHW6bajLlA
cU0iT0w/9f/5vbxze+KgyMkSSJDLJqDTkIi9llgkt4eBIMiVH/REDiQcj623bcnyWHep7u3xyLNL
9876djOPKM7hRNZ79hZhnw7B78SrqpI6coN87j9Gml8M890BpVkVLnuVByvPisnsq/6xDo6W+4IU
RbiiulvE+EsgF9rxNSoVXkJSaLE50DWSSnay7U9e5Ui53oTTMRKdDnbK/avdwOKVjteAHKvV0aE1
+0mC8aOnLC9JcDTKciR7eswGVDtahRc5f/fWweoSOc1d/Xteu9kNlhoU7B2nVvkkUA8ZbvA+isgO
JlqQM5sTEyV3vtAGQveDonTM4Vy7YcFsCUtRgdD+oUyefMONqCXBI9mX0SHWYmNQ7Mm1Ws9zV0i2
fz8pRnFqhtqrIc7AvsaFAEKMWXWt9lkTZK4DHXcdWBxUVX318twpup8Jazs9sfax58RGt3qd70Q3
nZX7zP6TiLlVTLlnU+R3/AVENGnhIUTuF1myKiDrPAuwBHlTA1yHhN+imOhUI4R1DGPhC566bO1N
nx5cS/CLGr4LYeopo3komp3rTMhm8Ij1yyCD+HGhIXCT+AWFiWk6VZSrAY+4aY2rKJhNAb151V9Q
tCHBHXM1KHhujE7/EDzWq3eILbmwAf7El4h/7/e6JnoQOX+H5R4fhmFFz8ms/bKC+7unJOpwne+I
dUwzt6LgNOT2AJcV8mOfWIquwqLuf7nXXd4/IA8peGmhIBraX5i8Szis/cbN4ekOcDpbl2a1JVD/
yfWO+S5ms6w0aCAjBVauekWGl403N2krmSU14Hp+gwlD4LItPw/21l0GKGTyBHfQRcgR1AOoigF+
JwE+H+qn8rv85nU4Kc9CcuJJAF+LJ6njThVgHTslQkhinOcI6x9LQ42OMlM6aVGseXm5EvpXmb5B
zEuj8sPHziRt+v6MbE6PQieqMliUSxsAX21kEnQZQDqclJ7dJtF0IgHbdtDo1kiilgOtvjqiiJx9
W1k8GUgeBxTm22jEzhZLiTP+Pu47zu9p20qrgX2AR4zZTyLSJ/bpKanzz5/c8dzSRqgPlSAcByXq
4Q6eg+HrtkWhU6Nvm/nW21nDa+gpFewmryxDlFHJuzh+hoia5UfsxoykNKKBC0q/5UEfaxgzwe2b
/vfwtgRsPp5EyFpOrBN1yyytEa4Wc+3Oe4hZxWrC+C5kWyDmVCNIC6o2Ps0TI6EEf9JChDayZbfD
r+ogpsR2XpS4VFiKRpvnXkrJyH7Cs4AQC9zk/RENrGb/rDB+hiES0eXufMtWzqfjk9YZTLKb5D4g
NYp1tHkNnzx9+BviYpv5qS+YTK2DIcrDvxQcmdDcWNsNkxMmv181i2ptpl/tPs/XGEA36yjgOcLt
hYH1pKY+U9zKFSQtU4vlbqeQkzrYC2Qi4TTSkhFD/9S2AQAFYU//Cq+mu4iSoMRJdMNayoSY+NvB
vSgS0xzOc0eFQ4byEyO5daolQ018GyXkyQTeKRf2ioieY1gNo/EBtoqqjL6mLGF57cNSfgv6a/Ji
tPolA46QI4LqBe4LspGU7Ts0RFEei2kMpoWspoOLduYzGwmCHo1Z6CWuUGtptQj0GFPxf8oW/gsT
+Q2e1bNzUQqugyZFtWTMvnc1t18inaqjX6/wthn2n9AjPBCBCKmGpPKKugtxGuRGvQjvAI45PZot
LdMhStV3X44yvjudoe48PcC7hH1MFzrAxu2SzRJ4BhURm63nQ3wHEKs5L+OMjlvo7XtqSLk3Yn8a
KwKBkZ/ZLqfmjDBeWLEAxuVH+g5uWnQfJUermdAV6NDIjioT/mD4vPPzqbA44f3ybpbZd+v42y0e
LE1lCim7/ZMSyvcxrLvTS71k54HcfK1qzgzAT6JstYkO/2JW7c2t3fi8S6NJyxzStHd2cDi1uzY4
p3jbDqFT9Gwdrm2bHNGfCdc/rW3JiBX04k0SAhQIZpLXhaeiB2ZWW38yG6/J02DO69Xp+JNsJyNi
aSSiUMLP0+AEmAzfkNPY9ZpGrCAkp6tlYyDBIQwokVOx3NzEjAeCkx2Bm3A+uzz8jXbhqhzEYg3h
paN3z4qVk/Y3LvD/pLGeclkG3+/f4gJff0bzD/ykjdzypgX+nR/76MyDsvmh3wvpCsu1PHB3TRAQ
+AFb2Fd3gYnvXLlO53wIYyhgb1rrPYraZOy/W4T9lWfj6petaAtCxMZdrgnjUpPZCo5DorOa7c1N
IL+R4BzjBv0zHFsQ3OO0y7OS47hvVGken0FdcyjsCD3RqQquKeYA25H6bVT9KOYGe2Gwu5IgJt81
Yk+D8WtfalClaWsu+qqc0i6tlAhcMYo6mhvpmjQiO+8IGHUszlYhuz82tuIV8xVfci05fnm0XRGH
AgMrU9iYITN3cXw0VD59Wg4bdPTkv6kxXF+1aNQqp3oG/kfMtH0NcHSBKIA9CxzV9xgfZ1kVSauT
5w0LHg4VHCsIN/3THWB1f/Rn5TT2NdfmsUBiD47QL+Kej6FLrtyyW1kL2Uc+loYVMz3fusLFFJvf
Ev5F92FajVPpJDh1RyErUqEreTFrmp3HBDOXL+nBfBrRq1h/qHfD8fSEj4cZ7n4Xwpv4KNxUxZh2
RAJyyqWimst2mL8020r6Qv/6fPV1+af0kGqNt5mF0SKDyrSwDje++mY11Ulf6UvmKVMzl3rnz2+D
er2k0HXmIyLUWkwzAJiBRorjyDr3o7x9VuO97eCP+k14L6Iuf12mXs/VqnG+eod2sFsc7tAirBrK
O8FxOkG35Zt/ZRLA5liY/2Ny2iAQqTDa0FZnl2Xu7Ob3mFSbsbRnpBol3WdaE286xRA5ufEMv1/S
Abz33Zm0rSUdfIAHhkatzSPVPMTFB8mOSYLp4Tf9oxEDsPXBVk7HR49HuKl0Qd0cL3D2LUI7WdAB
33OlTJ2VrYvIjFZPQVlE34WoQeVbktvvMcgNrWmaxcGXCnog6mQNYnoxJnt0eKz4ngXLUe0A6GUx
2F3AkiFXo1Oc5Bk4sUlrt/vb2stBHZgufHud2rTFQ4fu2cMRYIAewHVpuWtVkyBvmDl2k6sbzbbb
5SxULFglG+0otkJarEvVviJQ39SahVkLCIS/jTFisjn/Xw0m104hqfnM6t2JGp76uttaBxuVOBJq
zZihxiFm7nqYYTTXnsDQfY3//SgCb9DpXR4lsG0YLu8qhRn3Df0pnLnO1UBSD8GYGl3jwyi6cuPW
i08ZCg8sv0yvDYVNq1s68lltcc4XMjbWTXCIw7iDJ3QcyFx4OVF+qwKoeLimt2Xub+yPzH+ezi1C
126qClA0VDGtfrui+UlH8U48pZ+xGUJ8nuDeVIljWdIIlTFSH83yGe791EjAMncU9/jJd9E19GF4
nWwYiSzaHpbDAP2xWyVK3HZlj8ltzudBvbX5G+pGd1ymDoZKQbVA8Cb5+3n98TWSx4ESh14NaXrN
pi5ZflVsH8wfS4ByVvy0+HF4o73fumNE+8shaY0+v+t3fv0BpPljywcslEdgipOimasw/Oc5lqm8
CRQHZqr4JkbReDlTfuYGE70lCo18n7jRULjuyyGLPhQ6Ce9tmYwl+MyLAFzOSwtvTMAnkl2E6H4O
c3VPVYia9Vgg4CexfnhacsP4OO/mMTweybMR6dIUoGbPTWNgngQFUrwFlDbjfc+ls1gIX85krlT4
WZAk1A0CWtx9Gmkoza21wMbhErkVX8G3nu6JbNVYBqreDQXzTQ69BUFods4a9Z10mV0biWERHG5n
1MfrRYHf+OFh1Urja/9n0YB2px/alZCiVMXCB7raKePMg21RwhBLHlwMECvwQQ84AFpdYRmyLde3
4HpwbCg41bQ6swhIcU2FTc3O2S0hYvfretEfOUJuNaYuzkA468rNqznQlWXDqPGWxir5Vrv0Ey3x
pE1vaTo+cZT+egViWC1v0bO4DsHx4/N1//eTR1eIkPbXLNhWKgKQM+CVuunAJ/SDziD6zSRXRd70
+AmKhUe7Ao9tpL8ryXSuNECB3+zDPq1otIYd0ZfofDWigzRseo/nY7VVFZH9i1cvIqxoT2TjixrK
L1M76Kz/CEm88ibsnTKrTti95relsRZdgRWCKXoDjW9agkwH/pDktSUP6YeevUNMXsqCAYcwmiYy
izzMTGMaBUKOODMulPhxNEEJsAI9e26JUekQkWZJCCDMdircOnOMhWsoug6sU6xk6THsMn+cqCoH
dAjnZFahtN2dtMn0LKbVktQ73t+w46o2xRo5vQ0n1ysnnjOhLfobwqHSLJrFymwU0RKuAnVhuyAb
l++2n5Hz5mbJfnELbRWw2AixLL8ZhGTHioCJVu9FS55FOhKc0FfZr+roNVODzLWAKsikn08wPKOr
DZO6pRc+DuCJYclJo1000dkd1CmXjMm/3xlqVjtZEDQR5KPio75MNOMDWiXWeVcrMWH/NlUpb1bs
taxNYkUW3S6yd5XZ1yon4EmxDCZId0M0xmOWrOnR4yDX/qjkQJileQRgis2siFIN7tS1LTVNKqy5
H3+pi5x17ynyP555Rp+ZwXdZWqnb2s60qOz83dz/jgIT17IGpoaSJ2hI8y78eGGCI3SFN0rnuqgT
1nB2wFYulpvQOwYKM2KfjxEQc9+fjVvjxI/dLa18QcV23bSc89nanhjY1rgE7ZERqo0F/GdS0EUP
ZnL7YcRcKA7uNPTYlLEUrbVugkYh0+UVJg2YPyyGFHZypVYDb1I5G6VQK/Tg1SUZBOTXZ0zJGdTz
HaHPqKnx1KmJFMDkAz6w4Mkk8Zk481m0f29srCxJZWYn1fTnR9g0sI3vmGEOe1gjOPLCr2V/J2Pu
4eWJMneanR5pDEfWUDhsz/9htrujGwgwWAp5+RNrnPtqEs4kMBjSviVeXdd/FDSEt5mxJJ65qfqo
w9vljbPz48uXqkAB07/BUughQZdS+BQe9Nvvhm6CVjJwISjNYi2yh6nO0qO7A940vUQ+L29AoyCc
uMpIlmC5Zk0O3yShXk4eBRfYPfhBZoz9rsBKf7hfktw0cPlpCCSACsEwdMta7I3NPA7LAmVemfe1
xLZGZxukWs6GK7sj4+y+IC7ishxUoFF6+6oMaTlC3WZ0E4ZrtwANNNeOBXmX724Xxe7m5bt7A2Jq
92H3QeBZ37KUHgB7FDxWO3JVZuLmyrHyKjNg7oD1dAW51ctdSyIHoizevIa/+pgik2P+SK52kmXD
H4g/Sye+XJICLupnkGgPtvnse/JHmR0NB/cKebhwCbWafTc8bsS5njQPnjOcWOoSNimhUjIxJG/s
qg2VZ0HPv2tOnqyVgrHp7i3mWHPi6z5qZUnjlgBoKQiHgxEQDZZwkW2f8NFpMghr8eSETjdyKIQ4
U5BG9/2c5A3wmFAIkBvkq5zmfcPrFtWHL+y2Q43oOlHb5H2OQSoCBpPDAQTgFuXt+6yv6EHvTut0
NKJM+IDCADBn5beSztcvuSnlD538KozuJ/MjIQGMwvnINiq5gaJ0FAmSNyZhXmHRrAztChmq77y4
pw/1WVX0CkgW4lbNHW20o+upX6VUs9qVPNQGjPAtljFA1AABPNksgNUI+Y6eF5Y6n18EGKMnEQft
SLrqY6vo/1sihA93Ti9+hBkWp0zHCFdmcnikUH00pvf7zxX9L8vxB7QzHBAUmZHQ9Gs+g4bg31cs
yuknH6lfxx80u+ZYhM4ML0KxjpFPLaZHmDi5Y69eAg/yp/8MCcJHkS7ucqaP97rKE53tQdH+s+m4
u2Ib4wj/UG9Vm1tSdNBeWZ3qwtBi7uPpPD1U3zZY8g1LmFkXFsPMNMgRbxlwQC1lXzKVswFJIOUI
8bssi+ZQG3I7RJDFRsGTqWz93ryalxV1XmlEWnHMjWFxk9mmFmjM37NzT91vaj7qhY7UMyaNiWUq
ObV3lcIZ6l91YsWSUcTd3FIRYo1/whQp8DuKFiafkwyquzbC1W3p/ifa5lASouBU6vDn2QQV6q/N
PyBR7LsP901Yz9SRGQUd5OFiMYYgkiK9amQi7B3WE/pELX0Wzijd3fvBAWHWc6jyIIxYchtFCP9h
r6CJiewRM0R3rv/beXpTuSwgtn2QO5wqaOyyRt0PuMsGDsFC2Yj3nR+nEDUFFOXiqztvjEX+vGui
DcRLo8XenqAsmOz+hqeqP1iutdpJdZJeg+5POPX6S6ggFnAG1HYk0GLx6T3xCCvRYwPf0s9UsjH/
aZu6Jv3HiRXLevkyAYPI2ynu3YD7MYWga+7z8bTdCcTqf/Qr4kVN6X+KuJrcKr6wqZGoDEz4mKCa
EnA+1zuIn3humrgxqcPOT/jwsJH/OyJaahoGINd2sD1f8AVhswPU+4hSUiP3nxRY5Kk86McqaQ7Q
XRn59LcAfWXVI5izghRgtXDbCT9mfQ8zD3RhjeYOgicAhEztzPhFrIQjMcJZ45q5LbvfJ0T9MMQO
ZlCVBwRea7MwRrSsZHmPjLVCi4YDbx1GcAom2KOQvXN3rmH1FP11LMdacDTNr4N38dvcrgsEgARm
gY349/gxTE9XZOfy+8z6fgwjgT6NqEKdd6Z5qbavoSEY3/nOnPUB3WdVzrvHgd1+S4L0EHQp43Va
6uG+VQr/Qv5jCoWlq9b6xRFPhpB5FCta3lO+XikJ4OvySVccXUfTKm9KOPAqQGY5fwlixPn/K5KN
PEpZFOLZI7nqaGLhXV2n4a4Zqr37BDfOoiksYzyrUJLX9EaPW2ok+jwMcOIPBbgJVmJgXPKZzs2s
gkPsV2jgYqfCEL8Ez1O2ETj7P1C8mGxNOaCuxi3yjFZ1faGhkENOSUJQspiH06jf/kIJKRiuaWY8
emSZm7cKFYoyh8kKNuBjfKZJnvgksO+iKe9S9/scOVuwa3VIVXKgz5KrEDo0MzZ9a9wJ+/8we8jb
WfJju6U7XxZWlCuAY3ghsGKhpeE33gPZpUJaskfaHwJxVxLFf+9vjgz1k70F1HxlPwRTY6DZLmdj
ppJJt+HK9mg38gw+LAAh2mNQ9nFscUfBUB1dbBwakq1Ch99O0ZEwTutzrqEBuYNi6beMBq7mmB6v
SCh3kpdO7IKu5bh41q1M6tF/BzB0SBvi9Ij/DWxv8Rwv5FJ6VH5vOWefiENU7a/gHJblWqt+Ydvw
65JrX7F0uSimWUHfjDhtN2Sml3BGyQuHOd3Nd0ZfWF9Px2zhglletBiYJrFzpH4hNsPTZom4DWND
7sdifXGTAcZEvoCOuYGnMXSTJH4GnhgQwkLw+9tDldA5YRFolwalU6IHIOo8+06yao+JaCrywZGR
4+Rqol6RZvEhcr6Rip4Ohg8li8aPB5pBBc5aMnnVn+3dcYfZIqqiThH6gqv7xRYx+/gP01TTolfJ
j1hBjrrtCnKHJI2/Nb/jrMPO6RDmFbhn3bRchgocOKgCg3PmzkBLJZmwxq/7JCgk0D0fnc7QFyxr
4Hqup52YH02BDmK+2GMNr+M3LBNsgAsIV2BZUlqvOTqIcZBgrJxRbrPisHwBNvJ4Zl2E+CakTSMr
TGzxiXdKIuViis6eRrbUBN8Q3FPt60mUfF8eDKX8zAsVu57SK9j8r205Ew0m9YwLYlLsyb6BDEsC
WhiDZ8cTu/K7tEIaQa21ryStI4A3/TcIUoDBFuT5VLDKzTAOHkCFkUGr/cktmL3Zgcm5fNomAzlT
usPoNgPalH9qHdwijPvRGNVwvMzyFE4V5iAYLGfxhPHs/22mEbF59v0iZ2J70vo/fdofa7hgwxHu
oVk9etIgchLtUJ0G1L7+77lf1VH+MHECSq+nJdVBJva6r0UzRiyDKSieoufrTerqj7m/UWYCjhIu
gg+Cp0Ph07hPnh1oDYiOW9euNttEZaPUVOtJD7stLsV1GGJBzT14Hldd/dEsrhuIfmURaRJiBU0D
5p8N9gvGHTSabYTjMNe6IK46v54vLoUOZh3spuOnn1/ZfZcOCi6yj6nrhbUfNyHmCuWLG9+HBQ1N
/evfp77oc+v03pe4AJgBco+d7Sfn/poNd/Qj3B/svR4EBNsP2tFwZBKA+JaXPckGxoGcr/j+ZGSS
dFw/NHrTsPRBKucaw0sQ2sknKv6SUsmPdMcynXGOS7WURwFGPTSWVxiUxtNJbpVepuXvdWmo/ZR4
yPbRdNYiBYYZX53lavhZnOoBogRgdDoA0ZIvxPYyG0YpbB1sYth0RBJRnCNu42pgK7KLuUKLDe4U
q/l7FI5vmB21GeJKZs5Akpmc8476mFcNOy8UFi6diCDXhFU64CyjkUI8euAt0Mp3mK7b88AhVP97
aatTddlM2iOgkm2D0v+WAEeGRyCR2dTAQgrHXA0xHDrrmpPdtICVRZw9PlPxmeVOuC2x6rem41HR
q1uBfx9RN8dreVqXIJOK6mzJgeAqkZXWX0KoglTkA8Lebu0b08y6d36R9AtPkPLn17fyPWcgm3tc
EnXjmneTpFYG0/RGUCyc6OgAclCksxE9BUPN7WvmYi/hhEjV81g6kA20+avoXNY9CO9MCLN+W0yg
Fc/mp+SGPQnhAkmUZO9cdQhVQGKJH6auCUW+CkYbF/EV+4COsB+/9XnBo4ggh0MG1xkboo9DYChI
u9ib9SweRWrmaw47tlf1g4xg6EJ1uDNYNOozi/D4xgoKJHNlkRi8yB989nQxwwjv9a/aeVNM9Xbi
2YdtTuv3fgMTZTgqPHZSFgQilBJ26dNEvOu3Jv5CzhuaqUwxUqsd3kuicA2fU526u+MuNNIMerBu
clPOfY+rxZbQz3UyJ3ClvBTKvO35mvKsme6GiaYKyibd9Xdcs4PPZV1G+lmAgvz8zN+IgmNE6H64
G4urc2yEzzCBgAqwkrBS4vVuYe9Y6u5wXu6cWezm6RuNS8sxVQZlCZRgIHJNLr7JCeyG5qzNDw97
yWdVrRmbg5AfcNiJMXgt7P2We14FR0sOAYLTWWMCQtj0BtWfnU5aOeSMLENhhFOFV6Gq8KbLcoH8
rXh+ATSwKTOCofJGH93J90SLdjj8OL4ZoY3M+JDF+CEKVYrhnvHKr6c3z9yBQIPPfEfEyEUA3W2s
4iZmqvlIluIW8UUaFTfe/B8fmHeyoEnBvSJ5zRgPqd670dfaZTWTF23/k8ZwiqKlOzlvQIfQsDw/
uuZgPvLFUStO0trxDhqzmMmSdrkIljWjnJSjMbHQ62FOwGHPm3zSla8Wk7TQGzW7gosiwxYmhShp
jW+5HU+plKV1gKCWuAwTkRAGx/Yxpt+xJnJtxvYHcYxcAZze55SmdmPztgGtrHaGcrlV4B3oQqZc
X1cRoxYZcRCqyZB/OVo3zGypMtGX9sXR3Dnw6ZJEgNnGQ1F6ULwUJxuuzGm1+WHu9q4E03H7/Z70
bIyHkiCCcuOVMvYZmauDK4qfhkv24NsxI2BnvKY9kknWEGzBupsd2U7qxI0g+S11rPBwxIGLvnZd
G/GZDiprKZkNHQnhMXDgVPw3zRtyTcGcO67fFd5M2MPG+Kpu2gTfRhnmjfSGmGRmgkX+WmtGshfC
K/aCLC50+V0rd4IBMplTAmw13kbqBpAOH9kNz6Z8Vz+3alKuSq8TENmRRjRJItecDmpHkf32Q5eN
DDmSZMXdnBz0j/+axzINnhmTBE2EuR1dKjQ3KEnlk3dabPkm/MfspoGDq9yIGw+QFoxFe8uNl6PW
wZMKuswKBy1iI9aAcLoEmGPpt/0Y6ccMYDbYkEJ4UC1LrxwgUrcYXd7PLZcSXcRfJD6x/5wXKnWG
Iu0ITGj3GeMfwKrWcQDOIfjmfxgj0sNqQFT4+Twvr/XawMq45NAmmRjNSVTPzhK832KEHhpwYmuJ
54nofAh/0yDJaJL9jDWszsVPnABpRf3dCIPofGHXbYQlYE/r9Zog6qNwt4ug23MpmLmr5rQZ4l15
nAjkDlKFn+vw3XooDK44ROr9n6TJaKp8EdeHB6Lwxf/s2OiyBFvN1p8VNadSG8STsZt70N+7KQnF
bkQssy4fEUTsYK9UaA7ZpUxNUTn0rwlQgZxpt66l/3lz7yXw9bmXw6cppbN3M/pWMbPTiZnKqaLb
QX4c/1LoivbxGuyiYf5rt3RcRxqxL4j94Is0XfSQNwUhJLAXRcEG84RufyxC1n+6yQrVcI2bLeZz
zxSkbP1tVJb9NdCuz8g6+7c7uK/Vq/HMvw8lKKdg2kAlgoSVvTWY23ar5eNJ1UaW05kXvL/ay89w
SW8uAKc1+nTqY90RVt8FBZUnGvuIu6hPmlHIwFom+bjezb3umUCdOvWlpvJvtUuDO4dUG03fMLOe
UMbeJP/FevXV3V+sbMPBPcYv75IpQ9v7fL+o3aVoBhtKNISzNGqiX76pxwzbvzBmHtmtnhm1AQIf
GPITwn2yIp7JhjouDKi3qnGP/ng57HZUj8k2jD2zXAhpRbDi33TfRwcxeOwDKW+7V6B3wJ+7sIiB
Sq6d6EM0UE6HhkS+hoJ8lZDHkbi1ZA9N5nmj3bbCgxVkuBpPifFzGqah2ouQcwkSsnNIW11MeilS
wDjrn12/phkZQ/FcOoQOayAZFx0h4yEF1uPpEFmUqU8E/Pt8mVH/uojAwYCUh9jkF0fdBgCH2sFI
aiIRbEqa0SnSa1nbW52iaDx324OwNIrNWwv8qs8lhyC5hwPny1KO6BlP8HZ9TuUk4KGTmaC78vn9
bmYa9NL1sJn8riYGMEtiSnGsHqk9jRqD0q01n6MOkQfJ9BiQoGmQFLx4os6i+jy2idQc6fwakVfN
TTIpaFz/0ab1HVYnfapv7VQzeb65FYEC+VookohqRW2awN3i8WBAKtaMIv6R3eU16rz/Ced9PBnf
L4whyvxHIJVAxc+ooKj8aic3HScSDci3/VZKt7aApsYk/gVvjrXJS4h9a7QzaqpZcbxnlKQtsuUo
3t265vorBjSG3ATEhkTX+1+0l3xXRD3YMPG8BeP0C2TK1qdrCJuYNPXB5KJZd6TOujzA8IzPTlYe
qtXJkwXg8zmwrIFi8awzWwsKT8LlIyuvENRF4/Dyu31antbxdtw7wDh5wJ6drVzlKsIeExqOWGHz
w+K5rT8q+VLMYMj6GllZ5z2cGKJGsxgt6Ei9IaCBCLYcxyuIWr9vVAFGpz7MN0If/NVtUgu8VD67
kH5yAF3B5R2RodDMzBZpdClH9ubftS+Bbfh9cvbUEoo8hkPZeOKn+vyrdb1fkGOlzGqt+rBH+Hl1
ecIEPvUVZxHIfzB6/pwsBeDVDZl/nF9okD26lx8f23EjuVnnobiUh13Y0TFPbXDWO/Qzvz4ZMRWG
X4d+q1IXDSrGYYL64phXkun6hTlmG/9lQjtaGRmPibEytuUdvbESuq9WNBw57XBYn04Adi1Kk7Fe
0mS8Gvy01TPnDGwqkheQxpEOX3GH0CsNWrFymk2eLdjNKTiQdch30BXags+iwbeq4QaVSUFIEhd0
+EhtwWOiXv6lhfBYXCjwMw6dBBlK5NUgSgRLSFU8q7nW5xK0RklH3pbCxZpbcTKOJ54nrDEo8VXZ
IDEamnEBeK57L5S2WKNpXAYSBxSbhVcpzv7HHOGMFxdlrQTMAA/XcZ36y2NLWnNKFCHcMS/Cfaev
RfRet+GTR+3UkttSTgPkgyq1LWyjAW9JGcND7X4tNYsYecoBR1rcVYC7/h0xzqxaW2KAtJFkdXaj
ZTXqwr0wDapncLPAAqSLxgjdBL08mxZjvp0rXeY+Sz91vcpfPifyN3gXvba+Qm5tFn/kHIMf5RE+
IYp/dpqYykJxViI+cFM9hmS7T+kPZ8tZVCKGgZVetwnb2LowGb9/BUY0yscYC5Kjb110sAcZArhA
jCshTwrr1X0QTNcjGLj9qgYqksYP0Bi4cWcx1fiFe4kuZc9YxdLNvELO1chCv2N+D1olWtqBxWrT
dzchYEgzOB4hKfw+JR5mZNuKBFUmt2PybBjQf8/AN1zHZhYqDoFrHFV8BIYkG73+hSZ650IxoGXO
TtFqRBWLrVzG0q0UAawEeldeFEHyeGUlrg2C2bLqYqCiE1WJPdmsE+mfLkDYZzGLHK6gVCdyerXf
h2RvtsFpqPMnr9n5/IpyA86BcI9pi2YXXVNGN9Pmty9qsZ5u++44kvL4+S3mmZOtZm6ElrLv4Q+U
mFwyMd95Ff6VHnDCHT94Rt8k3La0zVrvWcs0dZVX5aDjvjBh84S9xWBls/YKKtI9Bq41+5NTm1Ql
GWuPi+QupA8h0FN4N58hYr+L5F4PTuCHkyned3Y6BjW2PzwKyX4R+EfDkZq6+qUz+0uwEasfNVkD
9beu/3wa0a/oQ0vqjpHr8ZRmd+bh6xD3+Zn+JKPwsQXgiy/dqYP0RFyRolLBemHKdIp5He4aopVx
CQmK1kO/gO9zH8bq5J9uMhJZSFINHeNUX+nRwSsmcgQyywTkg+pGHRbR3ygjOfbNhrtlN+esN2oh
9PaChy+2W5IERg5tKsvVhCucUe5kTn4KHtaGBuqs4unOdCDTTttzUTle9s6+R5vuLyVferoVWhCA
TvjF5d9TZrfAh1tQ6PKhRGHgEm36ROlFRXihY8juS9s47qf4vcqPNzjzJjmQXXhv//LPmR1ZuClY
rI7BfAmxpUvSEHOu/+KSA0QUUDHBM9VOyPYKnJPo4TySVrECCc+LPgID9j3l6iuTXrvlNcAqLdtO
QBR8mSvHNJEg/zr64n+2EnpoaKeJqIk6vX5qu3+pJlloL77MPiwDfcfbzLa9iZhZS/DMl4umMxTN
AziQxwbMGyvjoI6eqsGcG+RhXCv4qK1a1/nM0E77jMa9qTQ8Iya9sQoyHWieKZwapwTCO1vKelpm
GD1xu9D8fF0HTBsNxVpv/zuqjcOI44OdstPPCm2J7HvOmMXCuOP1Fgwmz21be//OpfDdCGRkHqR1
Uu61emKLQSnNEVvAj/WmAjYCPNIYepNu8PUB06y89bdxUL/JjDNIMIiQEECfFLCvyMxfgKToFzk8
lF71S0EN4y+bir95S2Y4FMF5DoYYBNmkJVflUXf2iPQ00kAl5pivoyQ8IkzKX7remAvq7eAzxBY8
vWowvcdsAA08Xd8I9HGk2u1naloAsrnQqOjOf62fIThDfwMZ9PlF5l3Nkh9UzHXHA/0/w0AdMx6z
qjKmTnD86JYtCFallqSYh45R8B8SW9FlnZkxIbwZoxKZw2C8aRcimQb9UclDfKImnRWe0aIho4/u
EaCvfRhi0KnCYkpQBxj8ScPOporcCRw9EsB6HkFK9L7btHRSB6t92YSmD8h6Ex3zTvpYMp/n4tf+
6yz59DEgEAWtbOwNaGjG7bqAfnBEWvaNZvAFALHuWLVY71nkpHn7fIV36Ghn3ONkPhB8V75mnLaV
yeKxXOkokJ88P3Wd2nfNm4U1OfAUwfqPe+eTuBisJUvX4Hcctq1DBkxIczqZACFT3nBqqe7CcSP1
TrojkitSeWjRDfdmRDsVCt5PjCmHjyTdRP6oufUf0lVQsacF+Xjyb0V/l0hLUUIF2sHwtLZ9/YE3
FVIbcyQoGrtHbhPUeFISTMjqfTeAV0JUx8McHKCCkvyzw5ybLbgQn5xDwslG/Gu6CR8e4TLAEhGm
SJF93qk/ZcxQuLV35LeNYHibbOWgUbJfBlCaPvO/Pm2ugLw8twBvy7OkEyjSpGPfC5MegISVyC34
gNKkmlutmOcMSzd8YpKYTTP0L2dD4hk2janhbWyD43TjStcQcLW7lcTQI3WEFOPoLvVY07D521aM
xrxL8awKao2aDpR6vX/WdpKs0k+JDAOyul74SSwE9XoWwfFVXEBUyA5B6SxVrG3MZCt7RcR+JZEu
NAC0uCyqcd+9EksvA99Um37+8ct2YLhjA1dUNOashOzNagZlQRz8jmE0J1ylIlVrMFl8rYKwOBHl
I1V8bh6YIZEsQyNoxTt4zKFuDYUB6ndZGh2vZgzjotiGMld1McrbyC6lzEff+32+lGfxOnR4xgJv
dvWQU/j7LshNiSa4LgUjp0O8/oErsKeo2MF0nabMS67bf+1Umw5iQ0Evfy+IXPYSS7ml+lCNErpW
FutRyOvLcQQGrbl313ZWwbU/46FJugLt1t15AJnUuV1kIhvY7AkJ7j11y1dI14yO3M3pgjabxx1n
iVbmTImqgl9duTsVWQ7RcYQTPimPdl6sI8xuhdah0Pn030A17znh1m3eSvMfFlP7JTPyIiBJfhGF
s9q2lC5jwLO/1Q6DhQUd+BSBlRGuTDnfhSvQgcsV5uXQHZkSHOUgex8UwjDoWhoYhg+2/679gO8s
tvH7uUOHQ6WRSein8Rr1ptrfiEhHOMRKs/TjI23xM8aWIGOoPRq8x+xcWvoFVuDGxqQfw5OPd++d
1ODFPCfl5x4gay1xY7g+vv65Cnu8w9iDSiHBenOQ2gpK0QcrXxu41OXsvMFtKYIJ1qFGfTb83Hx0
/lLy1jJhLGsJ2UxZ+tUThDl2OztFWBV7xIy+skIhifdShkORbXnLFkPJepnpLQMvA90ZlpQD68PF
b1yuhE7NxKo5pf+k4vhsmqzubk76PQlPlAM223nqWAQVZO8p3O7SPA2LHLaPL3owzoHefSw3EH9G
9FawCjPRVdWyEgMxAK7uoWCCixgSRNV/pO1qn22E2yqlDwTgs2vhb/d1gpMAHG86AmuRXkJd9+SC
UDQQ2nk/NF6E0eP+PaW6x86SEkZUkXeneHKV/ULdgJFmLwPu/qNZWuGUJ3O0pwHlrcVrkOUENk2j
yaz7FdvAkCrfoiOCIK8aJRjKQtROgjyJQg3DAZrKPOSn+MfzSgATeud6pRV0hue+GnQ9whjxvkUN
sI8sxoiYiZzAupTwZz0pudrio+LuzjRX5tPAI3fmBePz6ij9YuCZzHLGxJR3dVcEvq0YVsBgsm8b
pg8W8eXOcCOUuVO3ynMX7b9i3WQgSJpBBp8tldmFoaYYtCG62TTNgPeFJoQGyVCDKPkNjOSAOij2
yWjDh+ybJNWpcPuh1qn/XMiQ8daAsiU71CTNksyBYxJRsxySdefjLKMNU4th5hk0StrokJHmrU+2
Ea/yeRM5ti5yUzWPNp0TOF+9juyXfw0QMxu/hOM5YgSviP85hOswj//kXklhYlQSsNdR16zx35SM
nXp3RVfVwZHWQc+ZW1mxdUIvrHg7Pd+3xbbSdM0nI+Ufd9ZwDNJsHs53QdH0WVfSjehCQ3o2hLqc
aTgx2xjDEQ5XWxucLeO/MldSrjJzfxmcu12TglHMAyZYUt92dpjCm58x7doiDY7XpVUcblX5odwM
U1CKgiyfZknPXX1YddRlYXxHHA5zBPADbJzL5EH0BCz4KvgGkcsMAp6xKDvXo6WMgGCOe9kLJozb
JcqeagAExfzxtVY2spNRTSD5VgRbJoYicqrKN6pDdfoPPDu8fK7FJJeBtyLGz6hU0XESOwuGU9z3
ow1dU5qz0dISUdQHBkuvemGlqF1o983vtr3wcK0ldL85pHFisKwjXL105Vw+va4cieHtdgff2fIF
nuACrPKch7sujsMXx5EFQkCOKcWEc40YUsgSOQuERAkMmJ6T1gLwLydZYdwg9WplEd2yLd9DWbQ1
lA1n2Zk5VnUycded5ZPcLzDuAXHDkfRaOhUA87WuZ+BJhrD45cqepPG2X6O80WTGSOLfbazdmKPf
7cxLgN9E/6kWn5gAT4n9xpYKwBS+i1SRfF7uisdmsvpv6s2bYYhdLAYSzjQmptlYxdHajKhciHrs
sA0uvo9X5TychL+MiVHqgjKVt8jzrN1cxii2T7s9tsBJNI93HuPnV+pokKB04DvDN8194xGtv3BL
lSEGKjS97oSp4S9Fa7BhDBLVoxugmtdxekvOv1MMbANo3TVZ32AuZEE2JUhzsRjsIASzTp38+y6Q
kToX051ouyYUEn7MVxQVkhl86Wn7QSrOdqHzIhY1QkkUQ8z/t+4G3W2oDURpzGkem2OXyzsU08Gw
V4cDPvge5M/nZNThEBaEKGj601OQ+r3lc6Imus8fVVTsCUyVrNGeWYg2+AlfYuCLVi4NSMCCRBZP
KKLLrRgSZoBHQDa/xcKHdacrvND2fHZpPKnjHWfu6pBj6OlfEnGVgZiNPLI0s+bmATuNvcKGvkem
UONjFXUWrjig064BRe1Y8rb0Es7hAJLp8K2UXbOtnxCVMroSErpcp5Tzr6LKPH4jpsrpWpe1jMnK
fPfZSUTgCsYgOtuXLTo3Cg3da3rLTQmpdE0iLH1NJ/joRYTOPLIfEzED2wqSBqsTHu6EOpHjLuPk
akzqoErTnos5hLcJWKI6xa4YafKJA0j3e54C359FKcHzx8CLSkj8kPznD7G7rpqWi0muEbckvJie
1RRFrlZSrqLYh3L+BtPPNJi8YiGCdqvHu8QnK32rY+kATOJqkfEfis790p2qygMxMC3vOAhxfUby
f/P2GMMG2u6t+a6vbtuyLrwDNfl+qauOySdU8Dy21/zcHpzK1VP9Qy/eqERAJ4jGOWBz/kEgS8zR
A7hfN0QXzCxT5iSzEtBpr9cjWpvP5V92qX1QCas1R6yda55/I1FPqjC8Rbwdpjog4sBQf6YJciAm
8xZz9r/oiEdE95s5nHHhkSEQ/5mz9ikNzbaemd7ru6LN5BxLgJOJI9gUW4BXnPB56ScCOfWvib3D
ZdPtB5vNn8daFpdgLejcG6b89vMFZ8u0JxRWDMA8/Egimz7VBopRdo6GAtHr6hbR1mn6xAJLyipZ
5a6fvB394xr+4lNhastOzHGyYle5UkJaRIHL/ho/cqg3kkLbIS6l2WQHOayetNW8bMMYAm5G0Rw9
4g8Zl9QGZLW6HatlUGrby+lln9Zem05Aa/81MGcVknec9CpKEQCKGIoEXXlhWSy5cFiFmKi0NU/6
e/Kg9xjnID3UPeAizCIL4K5NqcV6LTOQ2hk1bjJvIH82zRESDr1h1Lss+es4QJXVyqJfDhqwI8fU
c7qHbGNZrnmKWCvhoukHseN+9Ye6ouC/WSvsdwGXExB8rVAQTf38aq/S5/liIN17AjV2x2JthHNv
N9Bh3t3ngvaSD7EpMIjpN5uuoaTZGcjDkjULciyEFsvqzMfkYa3Y6FOkxlhczxPGzop2A8CdaFWc
hp7p0A3L/kN0pBhJBshrMmal8nUysK3dcrUWwSbp/srArlCqbhznf0isQqRKoG0psc/Aa6fFI5oH
v/pTQdBSnvEiXeQKx/C9l03ngrWhiFfHV800uqv1OAe+c1m8zCokUMILaYlyEf9DAt1fKGqOvZk7
3seYaWthlTDKCinofxrbOo6L/v40kcHNLo9HYOGjpVpXle3MJplkiWYGGALzRAKOK4m531JtcVJT
c5vEsXRhyRtk9Px8k9b53eCPBDZ4gP11IEIqXPJHWOzpBzf1nc0GH3tLlEOI+J0yibIWVj+oJehh
uGYKtZHSk4aXlhBoXilwzCXqRc0isJv57IQHcGDTFy+LvKsJfuWPpXbqAHCbxR44UDrc6PKUGuRy
tk/lIn4vLu/MHNj8WS6cxMa7xeLrITl7FYBIt9IvhJ0FUjhowkSOFu166QibgkMgD8GqVNznev4a
EWrlch2/qEF80GYMfZPZdSOavrs31ECEYpI9LtIjGDQVBYmc4W9HL6Vz34gcepGN1rX0oMb0l3Cm
614QXYgwR/Bt1CoUTSsiLWagsjG4SNMZPHdEyyCNpNPHBxcZfDQswO79XOmP7u5N4V0J1s/pjeeq
oydyXoTi5MzrYugHH2uu5SgNaODgr+STgN/OqKivXrP42icM1mQUtAhSQTc1gx22ri3fnPREjfuZ
Js7Qe6hpDFIloumVoUk0cm4ECwlB1ZSefHPwbv48p3tqWS44OC7/C8H45yA+UU7TCOBgIyolBW3t
hUjwehuFOpphsFWrWxAj2s1u/osTP4OZy2cHUtyiOTLQGdVUM8rkOs/QI3bGmkdcCbgnLHNZHevk
AW05ITFHRBbGYzSZEfLr5UAFJ5C/YMSuW7+YITPUvySjdvgjxNd1dDZ/D1bZMXYCoh1UQcsU40CB
H7imoiY9twWzVTKWsasgMa6Uis3C2RArd64kxVBt+RYhAVf3+y0+TgS1nsCfjdlVhmb3j47A66W4
s8iAhtULRMNXmWdVhS7r4PFWSfqDWGAz7CRXTY0ns26XgyyUCC20LZVwMsQDDARGI7+QfJp0UCOg
2yQaJV/hwLrbZVaijWG6o5lg/G4rnrlRaxX5wafuGo5wV3xymc6MLN+FV460CDIr4EVOW647otQM
IzYFR34GIrIsaXZFlrAP55Yos9fkxOFdLrJTxVWcQNGx2UTqL4xVFCU5sajj8mUM6LHO49ogpd2h
Nbq0URzZSh/rZb8llwe6b8T3KPwuj8thKnnyCydCDlWBnwGEkW6ZyhJhuGAURDkC7jlWNeKpKscz
qIAc/7zIhZJixrrEEOC+3IwhcfgUB7ygnNjSb1/1MffFWnTDOj+0MQmyQJ6EmU8P2wnPqyo1UkBc
WtPLV2SBVpJ4kA9nyL0iUa3on6PaDDTW7tN9+FF+UxuFQ1FUwboq+rNJ2z4Zg61mFRbVfDcmppe1
j0eG2sigZnGA9jt70B3CPlGXRQEpL5UTdiVzEoyvRuKip0l7XRZCJUQb1Un7tO1mlFCCLMo7oLcs
bOvvzrpmbgPJjr4aAIqJiNJEY56117VTsKaPZGBAErU5SV/txJc6VIi9v/CEf7x7BsJXgtO/B6Mz
viLEudwstRAZJ4qzXhIISjkD+E7UEZd7FB5jTaodsa6U/D/PJkl63nCCKn2CZs2AXOgO65PU80ZX
r+Hk+4SvZrU0qB/Y66LcEji77P1iuJW98msvopMeo5yx1wNkn65JWLYoSvznBiZmO3a0il8+AQ2a
L++w+/auO5qCn0sZYRPKq8B50Jglqb/CtfYORuVp5vmPTF/wInDyzKQ2z8eHnfgyKRNxXu1Clute
X5E4J1TOSrWDN9XeanIeglAw5dHxpndZ6CJzo1MB+YSHD35LGzs1x688/vhnFwOKeiKn5DDBBsVD
y7hef7Lowb2YpimXq7jNumZ7BU1TJaa7+3FH9wd8LfY38BlLIKSSAXeahMDGHGoXYawRsdrVQvmj
W3W3oKZmUTWKnpaWsB/LeELWSe/tsnnPytkWMVduZIS094Iw8LJEvhqjhQcTXl7N1y7E5fWXJuAI
sr8FtgnJW2L29rnwaDPxjBz/MHX5OHl98g6ptAhk/SM/iGrAZHEiCvGHIGcivGtCq6F6sb+ifB7G
BOBhC99GDvpQe5uqpf4qLFwJhGTx2O4H4ihJ3Y6653szFuVnWYMFV9XB36ZKdyyXxsdufRv2lz/Z
9Y9pKENTJhTjHUH3GTKaBzK7ncIbT0vSKBWizYUMGCYwjO4ExzQqyzrU7Ou2oPTkXTyL7S+HKgul
B+DUWGoKDHsSRMhdvEyNdgDbhCpvD3OIWpVUWy8WVK9DjORyyiqxkBlAgS2j5e+uVZdYrLFDoQ4G
E/sJHtYPScgl7KrLwrTWPO+U4d72Bt2nEJGLebebsYZm0+fkYxkJLUPsgp/C+TgQVi8WLWtZX0Z0
KoiyjPE8wSqly4pvx6ILxbb/5wHckQLmPytgTtNlDw2tzWxdToB56kdlZth+iMNlPO4hsNn82Mdo
NodPocawnLUjtCSLOMAqSUWDwUtU6kXWFwkvbkokSZklwm1xl68TH87MxxqulbpkG5BoI/BpEOH9
UWCQbsYlRx+Gc/axHPIez6sA695hRD+C+mEvYiFHMuFurAid94OUx3RtLm9Zn3EPPlZttIgJG7zk
N7hJVP9n01iPZzUYx8SrcIyyhUW7in8eC5pkh84Y42mF3wK4wauoKHzggkGsIv4c70DEZzXabLKq
LUhf4rfSJNy7asjqnXtsKkud3lBeL8YzH2GZ2GNZEdH0GdRD+E1nhsVOLJXRNsxxdlRdbggQIA+p
pGcJTFlAO3/yFEqKyXZEFz+sQxEJKmuy8t/QRl+Oh35wEfQG27Uuqo191u/zMKjmlk7GFJW38HGv
vCzvsKjdx/YbcCcNvoAAKm0wwRt3ktaVwxi+k4HKB73iH2zbk5LZTENM8RHqA3ZUtZaNKdUqZnTv
KPyES07toXnDb8sJPj7hcrOLMVxeg8TblZfB1QlFquoAhswh5UQjR35rrOpKZmVfL2focb8yu6aR
2Hn3cs+fwzPI45x8sSm0w7INItZd0GQJVws9mK1n/j0Fb8kq8ObeNdfPTN8uI5f6xTVgeCHIn5Hq
QetFxx10oYBhMzYsqREgvNteXzfwv2Junn51Z/mtO8fpuF7dHOIGmNSNXbXUf/Jrc9GWV4LM96QL
JoHGa7i33Ccat5fldi7X0OJ8VP9dNoy837nGoWr4ADca/Kr1CLSedVhirvie2o66N3D22RAw6Oe4
6OztgTb5iWJHfK+RMIhbavwKRimhbTfCyBNK/YBsxl0GXzWmuN22DSXiYhd+89rxce2gj9teM1nb
Qlag3I/vGGCm3G3TZT90RIW2GLD4M8XSuyeSV+mma9qXqMFxLoFv+kzvQ/t5WEfyJvOeXrQs7rgf
oyPqNvoXSFzdgw+Gx+1InA338YxOadCG/TOYn+/of3ANZtEhf6CBaKX55jPvQexv0fpv3rrbWE53
1AQetz/EWpTloIfCDZqg5afUDQY/0tX8aMPee8lJf3JLn/hksluY6UcPPg6APbOJn6H5H3DBSJBG
qtwjpHPp9zHscaYNEgUArnMOt6kxmuqJ8YYL7kP6sg91EB9zz18JNbP7pWJlmHnWjTzRaIX9tsbn
ckSyxOITeolyqjGqzr7MgME9IchfNCj320EbS08iYu7toBU288+5dxBUKfE4y426bYesAFBndaB0
2bAOdVCEKtZsrmW4EH/KStVFFlQ03d408toHGjPKldJl1sqTqnUf2HaYweyjvipnjHKeQx0uixGf
2tJUMGXvTjfrk1eW9H/ArkRCVZYWbXcUwwjn5tE58jfdSGnjlxWQPxuaCxvgZZLOG8Qx+akxukbt
b9aerwgmXbmyV9ndJKZw/gIbbIKdngO357o+pd9Ry/OD0bz4dCZEaqgbva4L6vfYAeMCQbtP5p/w
cfGjwOEXCOmeWLCzh0H9InTLggol7MOqBB66wt+J2FR4wCw4AjGlfxbx2+f9AG0unFxwEkXivFYL
PYtNNYKLz6D6mPXl994fNewuRmFg11uUGeQl8uZEYu3KjvrXCboMWQ6IHqn2at1i5P8KfjM7zc1B
pxMiZ4oUJ2K0wADMYcMcPf0r/VhNxihR2anuePH4GIVYee++0vjrnUpJXP4YPwihkZR6fW4xugX7
ai2BH9qBertb6iThzHD4Y2uyUR0JbNapqw6NmVEnT1ejKCxbi/GTSI85lIgxRUv6dJspkNcwJOQN
vaOFSzThuip2Gf8lIwcCyYhONu1DghYp5VxlO4wyZDOvWb73ueJZBH54VQ7LLfsfYY4EmBdm8/IB
EInx+geCXx6WPWxKpe8snZQGA8iVlXlL9vtM0PEhZkAMm9hbzQtM3dErKGr4VWpPAUtWezahoG0O
e4IHYDhMeeqsl+rGTDZCPSYtbz4douR6L7Kiq0RTGB7Cf9RSJW+EE6VXr/i51N/2vMw5lR8twza3
llLCaBwyvEpbm5VB2EAw3oTUqHTspXqoegU3weIjCmSk4S2qhDxYWX7hfCXHZuaubrdW1HkPXBNm
uOw+TKBRHDJolqR6V70r74JetLgV9trzpGA2aj0HgvMMFwSfYzqFjtIVG8QGeTLxSRxkMzaseEVG
XbO2ZxO82ajEKWgr4NzwbFrcEDxj2xwSZG97ZFtutCM7fSVVCAWYv9thd8+iezHKX0AWKnfY373h
fzIIDOTO7YHOm+UVRLwxYRhmcmRa0WeWqumMaT5KRGnXyWVLY+Ko45uBBYsIR3quJWXuaOHbG8x9
r0PxjYxBkCAvLl2wziriHeisv+CD29848YqEyyFAL/g+tpdv2XZh6/qIK6JiOchhcX/dS0h5K/0e
E65rx6SryD/cfScHPWPgHHhAV8wqXKl3UaUpV86sDYylQ3U8npMK/mz/0p3k3fVPjvbrXj3P7XX9
iQwlkh6k3+jA6nOzkvhCWIp5fsFh35rAI0Y1Ig0HnWq8IKqFuUm1XYVjWySwhXYyh0z/KMEFRSdM
jMblqbe577yvXqwz/zWyO8wiMqHQg0Kq1+qkWck2hKkAMy6zzU639NEqPdzJaCSJbsglJwXqToFd
Vr2J8bK/UKh4vi9fuMMdQ47P50UXGyRQVDeOS5j9EPTpI86VRdK5kY6G2rV10S77ac/9wjmbfjhn
nTTthNs18W/07M1BxGjcpBpMaYc4XgrYUmmRppy6DwbfpkCo0Xd5ny5wTJdsSBW0hd30XHn6TnkC
SF4p1pTZqEO5l88tIAHeOS0FaMdhFiy2OQY8QLfyj4OiHoSQ0BC9bpacG3U3KX9YV4Q9QZt3CYA0
N3cCLTfoe7rpEdgfXA1nTdZJuh6JSehAkt/Ca5tDoaEhcQpwue19/BEOLhRfzhF7RRq/CU/sXIof
nLUopFxsMRMZPn9DPQZYWNIFulM7U5uZbGIuXxvFiGxnkbFbFUASB/laxIKedNONfvb87MlDvQX/
uHuXpxGv30FWy81BV5t9VbC7wCouP85927Bty+bupHVPnDHMjdIE3uH75e1Dm0C0/WjjTn6jxPl0
ZnRDtFWSqAmlPVNiTcxA6ug56QAJclv4F9LKmrhDau5sWk/D0dv3BqCZyGHb2C5YPZVFHSbyxLmw
DqLRmT0ce9r9ym165jVBa3FgbBxhhM5cNG9QUwJ6IGMRonB1WkQcPZfY50JE1LcR/lNEVkzZ94u+
5RbFXXhO4T/wZGelptva6xFP+FU5VIUDfZg0ZgmwAWh4fSB1u80j4KguktV/7JRlQzYoDmFAx6oW
wuHDkei+QBR/UR3jUjdZHFEfa2byOv4iDc75bbWZ93fyV1Pb37u306l7Ez34XIhaZ86Q78Rlu/3s
jWtHW2zWpxwFLxBJPMl6KCFcgXxZeJYe70oBz1nzVeocnu7R9WmW9Qaqv0SxAT1UgeyhQc424/9L
1El44AR/bYXrqV7bcHGfO1CF3gXFmVpTXP/8hXbvYemjYQMmqAHRyDFkgKdsdg9t9D47sF67LA1C
x+R5//QjicvoYTYaPQXLSJofO0Slcu+/8RjM9+Eyml5Ej8FvXcv68pukMsXcy0L4IXbcwpGmSHwK
vR2IORBB+T0ZszzTXxlSYw0Jfc52WApQLi0kaFy2uZzgKZG+pWiEqKeLWxwnU3fyZi+hVJRm9uGl
PzkQehEWH0+9V9fr/PexLG6S91TYk6qzb4LnXtfHSmjXo6jYUg7f7tTjjEs5CHjbd9S8yRQks8lJ
BL2wuSkgDnxTcqPTY0HyHVrldGv9joymNUbMPxM2VFT3W/frslPlnCRAUVBjPv1nIKxZlTwYcame
LuRuYVEfZ3kpbrudTewySVTXSHYOXFoyL/IJ587R2kuvelJeDUjGmOs3rh8ou62+JlIhCT7sAnU4
d0e0GVreDX72w18smeWtJ2PYhw+rfzvjA67B6MKS1wWeo3+T99u9UelEM7gRkK8ybEthFlt14Wag
hO858Ek/LVsdbn4lRArzh5ZsKMKBd7Hg/TtVUvO1uAMLKHLSnSq8snCniMcGP6uKAv6ZSuZblxD4
CtDCBoSYjwqI/og15UtGieZ1ITGPkXP7zdEIIkln6xALyzJ7345uKU+i8nIdbDuHEimCGm/H5hCM
5yqu6LWWpz4gLOj87jgexfuz5IsUQtihXWpxHwIPnamznfHmHC/Orwj0gNZ32N2Yyo/K0KwFwOhx
uEortQm2+FnEkxWag+jT757DEsU0pisQ2897NjZIHHR46C9HaWDnv4Pxls0nXSoid3XMnUy8/dXx
rGX5J2/gB2S8V7sDIo+BL4xj3KtYbV7pp82/CVWL3o+yOSQ8MCVRYPQZ5f4R+fx5v2Gxu6H0+vDU
3V/nT2vNAQNNYHvWL2M3UFza61RwsS7hwyi71nUnHEdkVYfF6AVRYb+oFh51IzPiC0Onx+J3GTn4
TQuU6xBBxzkwzbr02mxbCtfX+XUkx+1YWSERCPKOd4SWJon1cRmk1Cl+V+aN520G2G8/B7tQfoEy
MaV9EO1641uuSus+1ArRE9ScY4bZ3jWdN8sjZsqBygH+IzpNJaYj+9RO4dC3rSfXiTKuxsKSnklA
CnlkcWmRF3/ehigchfMkG3Xojw43kprcY/fGTua1myAZ+ytiCg1Q56Y5l6Tfk4dXRDTqxbFPrEbS
VUWcciB9hFOr9Gfbc4MYNH1No1D4BdVeCNo/sYq6Dsh+Cr+6w7q7swAAAYWlvk++W2RvQoQXeqep
9dia7kRpnBCVDe6mjLzevM83XKMJcJUn8inaylFUWQY6lZdqebNnMBkqSk1hb//efsmxXA3dCg+M
hLjmv+m3JO5SZijRGz19zsiwTuj1dCnidoFpU8ch/wxr/eLwQeaAcN4d++zjLUPZDGiONeRfG59u
UfmyRSPgQ7dtRZk8H4D4fKPDQjmRXIhimwxg6xL2yJLITAzyrEmGluD2Q3Pe0NmakP4xvECyWdPt
w+T5KI1c4Zqm1SvLDBFHUsT8k2x2m/z5Q2xtCoRlUWgIC/DExlDwfmL261XJDsdy9LTkISUv5R3m
9hV+seqmmBCR1cpAZhbX58lAM7ohh7jO2YMu86RAxGE+Mn3pDY0bahTaceqTIQIn/InvT09+kLXf
pY/h+vEh6C4H/Xlzf+TxxzRmA8dNEY0bDIFXDGeqnIRofM7v3s2uo3Ci1XEmyRnoo+90XCN/F8hs
ET6odd3+xP+gS69GvQiVVGHG0fiBmUvQmfCcpazaXw/04mD6lC2VK57oseLcc8FBs+DYY71nZd5b
e/Q5GeKe4/2eo2UhUT+2WrvIODjZGwCAUoqZ4vUWPRaKab49zCqQZQ6092yQP3jxvTHf9B+2NTnV
yHkdUgMKDflz1WyhNjQN32OxbKIY4+rR7sIhOni5r1ZLAwds+SUb5oahBrALru0Z3qENnlO3xGex
LUXUKXRrUP+tyrzmXuydaL6pJSseakoK/1sTIGVIP9Hyug68eZF1cJZQSb1Z4nzyBJztMkQEYR+P
/uB2TM46UUHEGYQaGl/vD37s8H09+gDZW96dMGlJaP36M1kMZwvWC5Rb3Hq68Ofcie6H2F3S+MjU
LuClhyo3rMQaM9VL+mY6ffApeOtCejyHIRPD3HFSHv6ER5uNnCZ7FDGuvCy3HcNntFwR1Em940g1
o9IOxLgrbZooi9azFSLTmG2alM1qbrLsD9qaWJl33eUQpPglRmeVBkS9/FvRUrWWdsxUYf5E56dj
hM84FHOfJdyV/jOejO3j0cMUZRLMpzRIs3XwuIeGLqfO+rYrgeeW/RG4wFVlEmrAbIZTx0W6fejw
XNzXuEfr/LVC8Sv5rvV46JLYbHfXiLUafwAdcwpY+AS9vgEV3/2NuRspA05iIzsZYdiAn+sc26XM
zh1RzHmjPGV+EqQ4oZM8T/2nvsS0F+wtjfApyVlehuzgRy6J2Waz6/o7htCPy9UHhIxrvdek6nwf
hJLQmCCgw20AbYIp/L73vKyM/NndOiw9zOMB/84ZOqLlca328JF+sLJCYxZ7heGNY/MFKzpfZ7D7
QB5UJQh+FAVtufIrCctbDa7PBkvSl6Cd0BPQBL2PYzUJQPEmwESpE8I3cIh/OyZ58h6KEr/3VVdX
BSG+w2099ix4zvqTufrEWQlkU+piCSxzHVxuu7RwGb+k/HqAuBJnvogb64gY5NZpRoArLbxo2swf
9LVxmsiJePaOBIc3WSY3obdurn7rgd7htoYW/FJr5xKwiugrAEDnslX0sFyRl0qC8O3XiZd3zdiq
rJkDeZooeMR9VeQG4Xd9vuiCuaAoAGvnj0pg9zED1yT0kZHIZYBNqZhOgNxqRcn+QvRuOGzUYqfn
6WA5ZBfaZb+4rG8qplauntfoY0/lRNJX9gdAXf09Md4b2YGogbc7Rqc75pHiUP4Fci7JxTuX/swb
lcD+fZFCwV7RKiJydFzYSI0/uxunEM9Iq1rr1PYj3pYRQRKl9ubIZAxnDkHJ3LZBZIjG5b3xKB94
53oTCT5n0Rupk9Uru0C34HTRIIJieL52y2SI+jwiGo1f+5wrYyRgZwGjhrOD4LfBUt+dEdG0U1cn
DR2BYohkakzwmMZAG4XGhGNSwqApuXHhnohk75Yn3nI1pvewGIUtmvwoivYfQcr0atlxRD8xiufU
xuox4+gzrBvVQQXCBPPjpjT2ljlCK12C8bgkA47PSddp3BY8awh33od7cyw7sqjHX7XRfG16ZfFF
Q+wTGxZzTDMJHbXdU1oaI+YEdFoSpTZknza5fqacXjWhW8G4CbK96ZAety10RgHN/J7Pjv5g40PT
/MuIfPGgCCwt/u2ZuCzo3D9zD9DsITpuOQokmMouIvyEH06U2xafmOZ4wNNpPiSjDvYfRP4mJ7rz
aLujy7MuPqJszzS8Bw4CRE6pHLSpU9ZDzZbyhxrKLfllm3QqfJQc3rAMddwqaxh8HrF9fv9fj6/Y
aY56V9II72Jxs4PxIGVwVXLu67EMhtsAku0Rwbxv3sIA91UFpRSCYkPzbIp/GqutZGOigCewgwXL
b5tKERxlBICrbzqB7TL5R7QFud3emsZ2CdKM+za0cZWAda0dvn3Hs4jOtYXtX8uUM8l70FnExHhp
EK7ySIwIf7IFKAYkrHr2+SpDCduKR2aDwb87hbq1kbCC9aaeRl78N1cFnOSABrIIy+qPQplp6ETn
slu4RaxrsDrGTQ4BhcssimUu/8kkjPPW4IyjzRVkV9e5zcy/Tb+ujiRqMyBH7iiUBO33D9uIFFFC
tmb0EeTQYfVM4gq30ONCL3cp2lhPRHDHB54SKPYyOtMjnTzD2UxjIlbBPaW4k3Mml7rvaH8GFMBX
y05JGHu8niZD2IybbGvgQiHV1YkrV9oIEpCkNye0Grgq0qEIsPh5/Bjn/TZm5fVFglzOlWLdVcxc
Bx6WiSS0MYCaKzjdteiLRCqpZ7Lx4sqFuw2kGWSA6CxEYEdtnHpKo/w5MXMNmnz1S/7lfPwljtgw
Pc9zJH3Td0v6+Qr2rj9z0YDUXtw17hR2RsTg57l482ziXAMiT8phyG/7c0U4GO2DzhmhaW1MmQsH
fs3rdghP3tzJVr+q8fqY98PtUpa/ddyzfOwPLr6jjHQGoLPTIzaE/SX8C1uaWvXQRc3hV+nghca+
imYCjcC6DtkMDYVoLn6YmFOqifOsCRuvRM7J2LyLlTjXxXZcBeoHNE9aOUcpWKcNAfeo4j/v6YIy
P15iwCzEfQpqXQKQ0ZRd5tgUGq7f1uhDnm8Pc5NV/1OBrmFLmjCrhcZ8DcBRDtF2pldlJLVyViCb
s3CU3wEXi65V//JH1Se5Pb69l/3fXG3HCuCyT4hoQsn5bXKFQo4Cr/Bk7UNBaEwqpOkd/B+aFGXc
rsIkLoyXtbOdcNKFaD1STBZg1BXL+EQ8aaYvmEo9SocCK4FHaeRLbA8i41S7+fDxgstUtJbvri5b
gn5X4rxqjsH9h0sqYBP6RqwYNiq3+mfFseHbjTVx3wD/LvfXcqveOGF/egtI4joPxRIdoLQHaT4R
1aZ3gGSS6HPRwvIyuxFE4krpt4Q+fWNDaQbNmDo+LS9dj+r4mmaAX8Ky/J1/97M63zBPKDaEMGs0
UqNi3kATzlSJwykiv7drn7+ar4YeGcW6qIHyk4299Pgugsvz76H/5RNBNY36Z2MOYFvFnLCx9BRy
YFZXQuPNTCzWptlYmhSHIm+RmMDMnNQooB0HnyHIHnMA9wZfuQnU/sZj0XnQGg54ZtTNr4ua8U5C
mrM8A3H5Z3nfbplzBc7G5KVxx4XEmWabgQv0Tm7D/NNbj8sHyT75JNusZfc61i0AiRs6ZYSj7mBy
EvJ/8hcSzWihE2LEotTi/Fw73A99878PTcSjzf8ER/9O4xY1l04wSeBU7ZIPXGsXPb5X54H52oYc
4t7v6ZXPA4YBLksuNKON83RyhJMHiCHUDqZjQ2ntyTS+gzTJqMinBwU+zWOtYMgQTDhLGXajxcrR
uwI2Oytl2zMvDl1RhGcW2pYv6ReJF3lBLsOyG44ksCYZayN9QsxqqztRhz5rF1xIH1ky0pFQjlxo
FJTvPkORIJJtKg21W/YdTIcE2kp8iu7HPlVDtV/pZ1uL00Iz7PHsIFy0gTAJyLVhUm500sMjqMay
lzPx41YeuTwitoiay6ns+4EcavEKFKYIJ2cJvMnVcRJy5jPR5U/rqCXQT1SriNH3vJDP9YmJwx6I
aa1kZR8f0+AuOGc82QL+LDNH9+Itmwx+zgq4LXZVSG0dqEOJOG7m4Bx9nB0xvy54H6E0bsiw8tC1
FG919VLfQmr4+0DAG7olFn8E80UEKkDygElhxpoWGg3ZX2CIAV/UgZUvmzg+6eqHZ99VuJJ+sFv3
lnTQ9YL2aDz6gkd8Lp6GmSr1OCpr46ApzrqigY/41hj5k2SusQsWhw6LsLNLb4DmtLXLBNv6wfFO
GRiKycHWiZtR8rXF4aLqb1q1U/DSAVkynLHyuSlJZfiSz2YeVLDYGjVpLQ5f7QOsjjwXfEYPAJDo
dKoQhPtGymWk1ljL2XJhPNXcgICsKOkw480K8sssZUOpETsnzXIrn6mSY83EJby4bGe0ImxGk+NO
2J2A822UcZshBQ4xF8sbTmKEY9fijMlliXeawxlXXbGoVjICQRu/OXlI9cTzBCUylYUYQL3HykXa
c6a7bxuAAbTrVOM3BHwpEwQj96iXkYkX+OEZpxnM4cKi6uyeQ36wALQcn6WXR2Bj7P0LKckPC5bL
ulYppQPtGfAPKYXof154Xrsk6oaw3rlpVDFQ9fAQWEaJ0E1vgw/E+bdJyw45t1y+6ilOr3P2F+g0
PhuCyu+sx9qBhmUjFK9veWK64tvt03KOUGiwDG6kB/yQO38Pa3poVdrJkIzZ952cs8TohEBDF3+a
73Zzkach42rsYl3w0QRIQpu5wA8kJrR0hAZ6qNdmHvnrRmtZw9ck2fclcLJ2dDQFlcWsaHmqivzq
tzn4X3xndVt7xYhvcCpTS2ZEi/gNsMYyH9flHQIaGxILf4b56POPr6u2/FWC/Hk3bmf8WS9s+bR7
32LBc8Ij6MVd/727p/0ixkBp5ZWrL63fAbmQ5vYMuoErI/BDEW2pQQFsswxceHxOmfCRpG6S2K15
eow+kiXFaR5y8eglY84khN1obAFStqN8Rk/jANaMwN3PjPuNxAcSHebJNu/CXPvS7XR50OBeBd0X
8201ECYMgswA0qaBUOjFSz0zW3w7UOXDBySjGmFIQ7RoJUEQjjzkhtroZN5P3R98jjatx3l5oL28
W4wvsEA3Hbq93wwwR6oNHaMWMLdlsVry571+Gl7ivTpTcnB3gVS7/y5mHc3WDVT+iuhN2nuNkFQ/
QRDMwRIAJ/YM5nToijEc/6l+6qvmtSrH/AEYr7knGG9D1Oj0g1A5K4jea2BmahkkwEJD9ZJHVtje
hbua/qwp5dx+ZvRq9q/IUtZM5FIWOtSq3F3zEm3iZxWAHJ9kA8t/PuR0yv6vtc4y2aANYceOtwvp
DoZSnLqEX1oD1puh4XpGnXRiUj27GinZ5jiRZwZhGHWp4Id/Rp0a6VsMQ97ttr2Gr74unF1gm1nf
emUFIYiynXPgR1qC3SRt6LC1kBKX0j+oCWBHGJJ44c/HUxEtFMbUPRzFVz2LHjc4hQ8k91BBPZnq
j4aUgJvfoyK/6sbVh0d1qJ7QRbXhbFDK/ydQ6MOkWyWB0NVpeaE0KkX9P9zR0dBxws8xD2Idw7kC
YIHu+L/NE9bTRLANewNo+fKl08OxqE+mjHG64vqdzKY+bDay/P7eJqe88zuaZnOF6Xv22wajPgep
ExOMUKutd+g/jEoX5l3THNnXavHOLuYd/GMmY+AZktn2K/okJq/GuMKns0UAHmxHdtX333IpVCov
HyD1Rdysafx+rxxS/adqKFp5uZ1Ip//d3IgSuxZneNbjcLUNoKFNcipp3ncw3IH4hFQgaDhvlDTh
deo3ud/G+GAodML2pTFKg/PcTljbpN5b60JpItqPvyQzhGsw3VRu/o9fxP7HI4NOyetD/jGKxa2Z
pn4MCgumk2TVx3O3/xbaLHWULA6VLyGV3iff/zHXXv1nEkt4jThrValHpGKzC5DhxMlXQvqmq0zj
uUAddLvhdGeQPOZi9QeV0ic4KNTeUEioRm8OcLRf61zIkgCRO+TYlBawlR+Vks+U8/SVRlp2Yyu1
1a9Uj6xV52tb4mzjmDuGPN0eTgAP+pT4+7Gw6BHT56pEo/rQkGD9CALCl+dziVybWhqL3u4o8i3Q
v/aoZYNk7ImwYpGcupqpCgEMet71CJwCSQEkNBAu7UNYT5uh1nR7kIdMHlMh72b8qOdwEXrCsE94
o/8IMJ71Gbprbv+aVptZvIuMi4gynYsapf4qHiV0qPsitZFIxHKh+W0JpJa3kUJCe1mNhDbnzNCq
hllz375eGPOiHBMgrp4ol8WMmA84to0zTTSSj/GCS28ZkOSN5g7NteoBtcTCzhJ/lVMEtTIL0RQk
DO6Zz9CTREm17k0zGFJq0ybuXZOpmWYZbGZBtdDYmiF507mjRXwrayoIDUHPxH3BCf3J+U0mR4dN
eDG7V+5IipkEKWpsJmqFnTxngW9Q2zb0hFPsUiNXNo8ftBcF7/b7nH6V91kmGSVflDzgVhv7ZoeD
ED4rdFGGggVHZsW4hfTabYYyAtRA+X1L/z4C9XHSHIutBciXYG6QX3YyFL0zq1IJSJ+GpJNHWcEh
Kv8SP0F89q1gMSJi/Aw85JBxKp/aK6+megGn8mp5NAUgE7wm1s4/avSlELGZFWngnQM7kGRRPlC2
wUFf6aadFQJZrFselBDb6oHWTNDBlg8NF/f/jMs8Yz8lx2P0ocLPt3d8nKpisjr1ffm9UvmzkHKA
oz4FXuvirsWvZXfV2VtEgmtWdJEzI7bVe9R4/orhkg9JcA8eZ8I41av+2c12M42MuhgjSbaLLF59
Tuo65N2MixiMdJuLmpTffvcPCfYbpHwcp4XVhKl6SSaEeTdrW4mzVAQDIPso5027CKsepacMLpxV
zlR1dzku4ZRo0iYAZQJTdILEzcdwOubAJAR4TP8lDrAFH9OCtyjSw+mFNTESqhpjvSyRufOrS1zR
5rLO4cU1q9HGTEUhRfthHAPPf9gtPB7UikEBaqKJ/p7WTGqvP7b888MGX41JiKjVltGEAzywctmv
PVfHkK0bDAwWVy//y4RQSH/HBPIBGs4DF5I6HNQmKgl6goxYmYZkqVnAUUwnLwtTh6KZ8QYEy/9i
O7GRKfi90oA+LQ8fmJ87AFxoVtxKJYJBVbz38X/D+ejelcN6jat6dakcC+AdqO5PMEadXkJTumeO
R2gpTXVOkVb/23cHkqux08t9x8+VFzty06hayfz6bfrGHizhjnhuXGAJ5MFITzonoPtPT1vzwiHJ
irQ9CcMwZsE+SCQ1IejPcEuch5w/dA7DAwNEPXekw3vmr72xpTZtjPA02BarXbH4xp+VAJCIiB/u
eT1XhyVLvrzHMXj7a6ACGN+BIR7xiAtFdA0lMcC8YzYusaBzp378/jBb2dCO9kvu0iaD+rgxP4jv
CxpT+eAiQEuUxo6r5eUttgjwxHUY4j7nA2hDJcnEB9ZvGvFsdk8L9giel+CWsFO3ae/0nvscNwjr
8RvGrja/ctjNwfucTJJ7CIlJ+gASKOIzg+XZ17DGLsOCrv+UpaFspUKN6IuRcozwpBGZ6kP0f+Xt
113V6P9kKgUgH/QmuwQISh/oWx79h2E9ri3T/t9ADlrxAccjFouxCC6jB5tdzeHvQ3SoWtdsaXcp
d61oZKfACLLlNI4YT9L2S8qNtFe3wJXXcfKzFCr8h7t0Cfwj2N/5Nm1svG5ASGs59nYu4D6COi7w
ag65YjZPUwiL1b8nauYrjfptWhf+PbrxhVuTiInU9oNzFMDSUWMBQyXUTJgsHaWQKxSG5+s0QbUG
XIRJ8GlXSbM5G+hNIjcxFSdbbte+hxI/uw79myHqbjzRv1cWL8A64l+2bDeFzExpBR4/FqMx0G0y
/kY+xpwVKktuJIoiySSt48Nq/Z44dl+rMObKJt0j1HOO0s8FGbTeyt7DTgJPkB++G0GiN5a9yjI1
GIeC1WQr1kULe1588r5WXaR80rnndOkmk1hvaDTQfp2SY9+9BLVbmIIOavS1yCDQg/ZZsPQ+cqIS
NaV+j/pxgE6fEvSfQGdsYehsd0qezCJa6SZOX+9dsR9NpRw6t8vORDh7nDVf8GnugCqxAoJsLkN6
aGtkl6BJbbzX/F7xYD/HAES6ohdo2jF5e/1bK0Sv/6yuPiHiUGW2oIW/E8tgBQj+sebBDnpnNOXZ
yTAcPUE4+cFBai0rG7fKUEIzPuwSQtEWFAcsXVGuJHeMRD/dCpczdRG4sehI00iT+nZ3WifKySBF
yX+wkCyTpc6gYaTZhn0MJVYFEBa2aHvdoC2azc+Sgbo/xCa5Pgpq9iwMf17fFcUCRUKUrWeXJYfp
XE1wdPqETWZVh4jp7tEXUuwANCfJMJsBEipOXwkf/wUehXL2Wmlr0pkXfmFqQnQVb05Elmv/lBtO
P3qd8znZF/AhMk/6Dh3rO+yBny6EzldBJAZDjy6P1iXnDQkUwYfrpN5kmGvV+Yx/3Tsf3JCBdsId
cnkKPfz28Z4yqB26JjfTxfGTKsqwycQXYbv6RnrafGDoczmRljVKzLGC3l0CYIOyNPhbxPvxiYI3
yk3tpyczk6CtvZ6/GPrqyJbxZ4CIxSkHPnJeyr2Mt5a31VxPizL0qUTMd2mKDh0L62m/Q3ABRU6M
I8lp/hPo4Sy0y1TL2c18QlWtPFn1EqHAE5nnVt8YVOJRxw4gHYRUm+YCcP3yTcStp0TUHn+ksQD0
MHvllB7Nu9U9+BrseP9dZuMyGjb/q6sDAqAmqOEeSbesZFTpVhADNE7KAh4IMTjDV6Zrs+lyFhT+
QIL4jB3bN5ylNnoEA9Zr29gM0wRiwyHoIJnxcTPPAKycGQgRUq7bywyY4Vxp+CM2Tq1/VkgBFX/L
pzhYRakMz7JZP+owkyS95L4QMFexIuwCCVltOEPv6+I12C9+XeDyP6PfwcuCtdYUfC9svAmlyDkw
Cr4r3qEp4bebLDp9BBLP/GOgnLTRWEXCJCZeR7TycViMWBADYO7oZfBpgBTMkjaGS//SG9/94oFs
afFCtXwLkAAOHvwG/CntguY20KQpsOr0ujjqypehs0WFjRrp6iT8kvU9jqDE5jv4AAwXt9N2ieI5
sjjP9YLH2H8lJIxrbNhcgyfjijtF6xuueBEGTJv0K3NwQimuaA9yK70cCeHf8AzbuHwvQnCQYEGm
UGER6dAEa6Rs7ZySlyb8M1vKNbfBO++i2JuK81jeAclGjFTmgiX6ndAz38xF24kHL0H+wki1VY5M
J5dWQ28KgBiogBJbrpiYQgzJjMwkh8uaHlPn5mE+S4he9pSfgEWdVVW29IUyZ88d6F7i9hU8vrxM
lzH+ZdrcGpcOvF2Te6Vwy1FbB+BmkfubWTDZ40gj4w1bdfPpdcSG6gTxxFB/WZGKFsM/RMavT+9j
EcfG1lacH7MrIZyk/cdCp+M5ylFcBAbk5qwShSMS1PA3U+Q1HjDkwyZ49kHfmBgwC/ef4BvI4tuX
FfA/uqxzhOifR3jo8/b8KQPM8LtTmrIT44FbQh1gpSAbkWV38xKyLUuELbcfqyb/D+AUk3SDltbk
9tC6++yAc58x/v8X563tQti/dCwtUeiYgKw+gFYfzY3JwU/MJ2M97SpFNwoF/gLY/IZqHoc+hBT4
bziYvvoavaHu1ZC5cYAN41bDraY8p1b9RaOmE+YvpTyANfJ+G0Kky4W0/8XKwDOxHYSnX+TdlThm
oyEHhsuBYeZp05X4J9Vi1cJ8iSPP89qX5yV7oE3ji2h3mJoQkJGhcS4CukRUbt7+J3sdGKrxTfmZ
sDfDhQ/JULKQ5o7L4Gu1ZjFTf3iP9//0idChtxYHC/2X+zox+/g1dIWQduKl1cWXY1Jt207IRkI8
76co1OGnfavGfoxanO3/ywu56I8Hw+87+1+TbBJT7YZ/w62lcEgjVblUM3cE1CxBcxG8piyqA0Ze
PfNCLAcrBh/TUsi88f6A3Q5heDQEVZdeh2ojjfB9QeYH3OaHtq8ukNNkKnWttktBM2y1VTISB5z0
rfKAJygfN8SJZ6xwRrmGon6CIPrcxVxT1XfW/+/Os8T6EkldUhKMnvCgsbPWJbNMXJ/8buX9QaYn
Jv6hOb887b6Y36FNKe5YWGA6FnXCKk9AnI/8QPSntBUSJnwwRrvoTbn7TCqblE/IXq1ZUIfIPawm
EQ/IzImVTUn4Evbzw5yOSeT/p8/Vutj9aigMJjCz2cfXA5kAhbuqRzQBPPN6U8PXGIPSDos+YUXV
sfMsL5dkFL+3+RyxtSTu+SiNON6lMN0UctqWGMIJI1iQxX8doVxk1yxu/GxK1MsaE0vGh/TYDY8N
UXcrYAEVf23IOEtpHLGKStMjkl93y9REMPF3Qp6wUr+D+tdWm76szJTRU32QEMjibbrGKxKwkfrN
EwCQpVhBv7SldVmWR+psyMBBLhoYJEXsBNWGT5Vh7bWg5W62WtAd3sZoopBeskZtABjVE9lMBoSz
N5m1vK3YnORrDHsz/P5mgTSEUjcD93eOnIb9LgNNkfO6BKHVfN/5y5IkUO5UgktVEtKz5Rrsz81w
bhMdGz2loID6UqvhPYTE0QbVpjupQT5EjTDOtvpSLHpymuYB9SIactoyEvSI7y1PnGhIEL2sDcOo
bXj7cpS6oby303SwuEUY35p0ncLwdnGS9XW+r95hGlXpRblCyqAdK/vL6AZJTt8DB7dWQoAjbB/l
bBvvd1jd5f4Av28vbGwmmGbbMfjcRJwQ6jRtFgDbjDA53/S0ybImDzk9dlt/Xueuc3Q5d3tt3Xa5
b3HIdWFLyIzLVyofdkvrVXURPcLY+Ve0ogGX21wP9YEo56/vkE4Qhtpyo8chxQ/fk0epIwCdQ6CD
GsKBLGbx1UDs2bflzw+NZkSOUtz8ry0nSji8A668PvvQ11RA5UInD3hag17uzlasN6OSzOpLXLPA
YbuxLIxpirCNPZddR81QJ5LoCA1okzrtRLsjVbz6NO9It2ZHUHHo5ahknIzLUavf+5zZAIzr9Fl0
wKgcK+xAg9J/guMnNUPfoByptS2t7/8pSQ5PC6tPR6uT14gcrelTdv0/i1s54szv7n8EaShCALMX
IIOIMn3+Qe0eWtdMY8U00eol1bdeRN4CFxT/HgAXJALcZsRCA9gZabO/oiPDzJqICBYivbH/rZdj
N5DfdUoxUL0R6ZU89HP16orCWeJ2DHjxQnfdLt/AZqQ/dPMWiepmKSqc4CAU7x074jRqYh+PvxCV
vH6Hmb0X1GtSkIQ+D0f9HgsZ8aQ/ngvVG/YU9zNDHxepuIWAOR6iDeMCvbd1b71IL17vCIKMkwsS
e3RRuxoaEkFst10kcvQ5mN8hoPeJvN8ltMyJqRq2KoyFhQXb9qM682cLHsDTyrSFKkHxSzWY3cUj
1biVwzu7KYQHJqknq6qTveP5PAxQLHVc7Ka08hc4iAon/QWGnoe1ImjnrIGZJvkyfE4+1bkQOkMs
VwX8q/6s+X/97/mD7ueuss6qIseOeH+jaNYaixoy2K+fyW6c4UnmhcAhvldOnqMkl0MH2Lo7jhMt
C3AQ8Pj9OTeHNix+sCPVU/VJ2Kj6U7QprohLXJZDaTo2DsztWwXoCkQnaYfR9bxcNNvzuFcUPrX8
YKceXmC5Qs9NsMcLC8N7zVZevgdkHaWMeUj6xB2FvYDFN1BlDMQPBCjSIbRKR7VSppUe44P/k+Zi
f/9y6QdaGvwANybenb4HhDcR1eXwa7MajJGsYcdjxihJcpQizf91GB79v8Kudu+5FhAxNzqYIxgg
G/n2HrTI4/Zl029PUt5J0P4beOETk0m3KwzufAlk//6Pj1Hd38mkWqN2gZF8BGzHQGVCZsrDJXBl
4EaU2zF9qx1uDAWkYjeCzoyN9sS0NZAIg5OUMxq0whmTqvRWTeRuPaqkx3ec7p+/weve0TLgxXMB
SWaYCBSoZ9/9BsuAhd+9vjK++ctMk+ndPbjXy1nHMMDce5Y2nDjhIlvOJ5095KTt4pRCnV3cuzZu
DsQf+jwQ4m1/57Tp/BgHL5wlTJro4d1fWUqZQ5blpHTczIRM3TaLNYFiIQIqhr6eFdDD7wMoqi4T
B0RRfNdOqh2FUTG5esmqaEEm88WCWiHU2XC6mwwGvTjMM2ZFF1835mx0uj+6+A4409z5bNFyTZoS
lu0TYL+HNiFy0qFaBEIIbIw00YSPzgohmsBWGslu7IRw8bijtUficLkVrcB0tBW41eOEbR5vvyaV
idziJ4TGg7nYUEXg/RwL5k8UPGNVyprYQoP/mRwZUomwlHpryAo/g9NU7St/D6jxRK//EvUckuKj
dqUtUH88pbx/gLAH1AeSKx4U2xC2O67ukoC5MRBZQ7WVRug6ppZDxKhEUXKYpvLXrZN9W65K/Ynf
7QkWyVYUw9vB0x1Sx2h6jf/gIckfLiR/y+AU7M3j5kbHaV8q49M9pnLX9RutSFqWx2Bxs6J2jBxM
q9Pme2pgAGh3vMHD5Dp7svq3lbDDbdRxhsWxD+FNjNGmGErDM1aATICP+p/qdNJySIya9syM7cU+
3j5vZenX+TItuKmnuLjAljTKBkeomzGLPOAEGfRltBI2tCbGk8gCVtKqq5C1yP0sGgoXkJWBAajQ
koQrVW67s1PYQIhJIMWVgyi0RNymFdydoCpv0lQC0mqYL0memQRFUbKXlq4gW3CFk4pOYJAiq3XV
ZdEoH2xluxY77HiggpdQCNEmlncl9+Qz+oK7L0saQ9xwhDmyb/3ijZXgumdvqxF4R0vI7r4qU9GG
/k64QNy2Hd7H5oncgtikce/5YYjCXQzu7y4OzjE6qZr8J1TIVr3WUgzz2tFYtO7gNE14SDLuih/H
o6e2Sla8gE+xyGXzi9cH8wdARWp+1djpF7QvDRSS+FiRrjjoCXcQfdcVlfJevZKgvoQk9XDR+kLA
HzkcI/363a4y+f8KfppEe96i4x4Uq/S+5OA3DAweZaWT/zpG/D5278rSf8kVEbUGWEdlMnoDF2pQ
rThON/nVK+TTPCh+3gHOikoWMx2Zf1op5fIIUz0DBdFra9VAo1/sNhKABEUPQBfkHpnxgVQuGvIA
0PSDw+NCc7gjqysZcxmQsuEtxhvW3mFjSqXKMV7UuA+YWH/IcyJZCgvx+t361YWmnBCPJD+TAcDu
QwKKlHlnUaQCneOsBtQIOuT1YjMoDIGVhEMhy2j7mOtj5OEmDceQ7pZ3WS2pGjomJoosAnsoU3G2
Pm5nVYWVhp1OfaSn+BkQRBiM5AlqQmHlalJdv3W59iGz9u6NQqEDruaOuqtfZfOJbcaeMFheWCOc
UDllu6mXNJZ7bgvzvisthRaXyhwUBSe2wCUQ6nBGRhzv0N9P9ZHRWMttZfP8C4rMwBqsEOFL33YZ
Q89d3pDdz+pr7VJDPeV5tvWujNOAZFUFlLm27VSTxGwfu4rAiboRavgRhGy7HDIqilTOffuqz5gF
urXuOxe0cUlRoB9NE+g5SAkYbnjHhZdukyTj3djqBOQGzx4xWrW0ZmJWq1WJkMRsA2dF2yHJy/xt
nbvptLZUaEZ/3fRVry+3jtT4yL4WU4P5sDWQ1k39YC7LIL67o5bvvYRnykKJqpKxJGtXgRHCyhp3
g0SMblnyji3VUKXDynowNNhe97JGVQpsFCiec8KU1BllFhXTTbw2fce5/O3KJfEz8xwPRAEbyGl9
cSHXHgvWYPnsiGANzcS33swyV5WR2PLgZMszu0pKkVT2bZx6bmxoZEc8wnGL8HjU0cp5U7m8y+q8
qEZEZWhgTvH/IsGb2vTObxOPnEXOvht//YmhY70F8bhwKgvilg7cwAyMw3WhvW0NSY0gn9EMLWzt
O30M6iIP8zkxUhPua5Gj6UKSCu901u6kYR+yIf/MPZvbLGZDWhusXw73EmZa6ThAM0IuBfAYfMQl
w6Y8Kl6gyeYj+79fgT3HLlWvmL30LxIpa5rRlIVLvAlQm/pDvewvejzAoRk3sa+Yv+8oFhPxVFHN
khaH3izVAiwEmIevYo6IZ9KmaNsoDn8fg0mzpHDJB6FnU9Oiy/u8G7l+Iwa5PvFVgcxmMHtb4gJh
sIDj1DjLiLvARmhBkx7Kn4diW2PX+UOsF0+N52xedtsWV2oaZv2ehNrQzZcpzwCapplb5PjeHxYn
aXjuR3p9IjOeDdSwhm4JGvrRT11GfzMQxpblK9BBw1pbBpmJzJJzFezpdMQqUaFaN45cTGotZev2
4ovxUvftCU10NAUlJcOZpU9GzAqm59NLyDo4gpmJx6k4d6wxZWyOiqLdzEA1ds6Pe1wd8tv7QlqY
rHRyMU0L+H36rljrAJMxyKdoPYz/2OEepYHMQali7ESHX4wHaiNEpzf0hJRwRCJySgAp7V9wiyX0
TQnhLKnfySU+2+MsJQJs0SBNtgB1ixTCN/fUEHeC9HhGPJ1Jnc0LYm3CzneXMRFav4Y28WAN/Ll3
7VCVvDqbWkKBZX7z5Gh+QlS1bdkegFAqFcI1LlnOavQaPejrfWrXKUT6bIs5UsvHhI+tUHGKoxQk
of3y56Mj+J5zFgxAEYiEV3wkjHEnD2sWtbPDgxVZJUjpc5qb8Vu9tiP8er68ml44feeQsVJ7SpQU
0SD359GgUSRcr/tB7qXOx+wDshbgqdogkSPjT6ib6aXr6DH+yEnEjYLHEr4N2WLGTH0gYlBYAogJ
t3zdVh1iL6PFIxcBJv3W2AH7ocgJ4qTss1r5Ge0DSekWAjZpkQs3zxiMTODSR2enr6WviYdlqxUj
kusBAROI2Pqv97d1er49tLpOiBRRsB/wWEfeyiDNJf9DLa64bZ3xL+ZWlb03IU1ugOU1H1/HJ/Je
e5ayu69CVR2ndcsy9aTzDtTpd4z0hA8kmEQkl8GUMFjcyArS6aJPWIB7pDF5Bqn0WlZKkS/FGq2g
2eDPv3ssRIU0tA510yU2MswDQCJR2kJuHeRTQ4/iEaMQOC0WyptIdMyZ9Fio0PgPFiOfPQQESDNv
EDKI53bUt47/fpeI26+1gMM/YCPdctTPbnaUWHwtTLrwouFVyq6Yd6ULpZwzm7wkRgMVM0XGDCY2
1ByfjRzycXQFC4wTenXpRaQKHCvGqHs2odEm2vvzPGWkcpxE6X6ZxDFzYXPJQD+yHWmrtwNQpl23
YsYTz+qZXrj5f8x/k+89v8t7KzAZLIe6KuB+eFVipIRCT+KS/migdeJke92GvCK0bL+C5l5MN89O
V/CY3c70fnU+aWAdTdxqyzRkUTc3HVwxGVKsBhcFgjYdvb74z4bvgwGO3l/nhrxas1TNDjfwJfOW
dHyC753B4WDBs3CfStRXVzahtQTqZDXE6hA5kTSUYJTWP+q+1GlOFDde1rlAls8/KXmvZSkpSKez
+a552cfeQfIpD0kFDSBcoqvZztk4fIy+tICWvL8A0fgbUNBqR+pPpBnCSflkBo9USQF2AAswModC
g/ZeKImwlJ/dWRb6au8ie1+snBk6Hq6RjLiv/Ys5ixeEtzEc926rL2pwsesv9sT04Dbpez/joFwH
4Fpru3YU0UXBOEPSDNY4M0tUNoeK4s4kbIKKc/5XRpkIyhOfWDLwBNzWZJk3PyqLqUSejjK/OGXO
4Uww4GJE5IhiTAkK6ycwsFoaKJPMKA4rw+ATXLN+MCIMx/RyaOtULH/JqTKcUuNoH8KtK/cjjRbP
f3wETEtke0LeA0ILmT2uVo61201XWcOsE2WohPaArQ/q8ldU/iXD0N/4/bGTZD1r06h4dFfbuP3Y
PjZPCZHjInoPvNL2AiFtqkIwR8MQhpZcCbMNoAVMftsdxsVumUfhHU5hbvn5z3Txf388CVZj9ZsB
woDq5djklc7lBN2Pq5pAvucFld1POgsk8uCuvf5mNgFztWx5iGZBaru3FaB5P7Ri3TywKdDo69SQ
8dpaODD1lg4STR/ZT1RJZBjtcVlMPhbgtUXNgXWguRiffbjp/E+zZCdKKY6HXSywMqWYqDZLpHfd
8ukqrSTdYWFm8UHZnyTeJEEraCrhQNihPfmLcqDhFF5l8VM08SL3Wocc8GcD1RZRmRdrIreWf1rE
xlHlo1Dih5NiA7he2znxspw5PdHIlRyY/wLoFY1D6AuGa+xb6UMA3HurX0R23JuIalRLlZHulCFx
911p8k5jGy6sD0pGXCM9lfVB4snrRBntzpGlhgpdRoK/dM/WBh9xue6VWdoOiQ+M169lyyz1eMFJ
B8/Vnu/KvnRUtiRd2pr/azuEJ+zreEXub+TL+wdYES2T/n/AXsMXi9thQC8gR4F1pFOeRT16oN12
0ffbeKqOuX1QYMBGBGUOEMuvKZDrQ4dfyGhRGXxfzJCqFzr5FwPvEP0Kz3lqKOYuTiGxl6sP816V
6NxbhHwPGbNqzRq/cUNy2ZkN8A4NX83myJWQy02bn6A4DAJcrxlmY9nFT5Ujl7IBqVDS1uQdOZPd
ZzfnRAf6q6ZnWGeBgHZ4VlBhnQB+ER2+FGyjXg4zQI6Mg5T7p6FhgTzNthIedaF9x1mlecX2nmdK
IoLcNPQRpyfcf+5YKtMZP1oepBz02bw/6gEHQIOUpClZghzK2L7B3chpDqjwrU69wLAPvwizIt9O
trruHuGglRim/sUA4pFclKe1ACsQQvFwIFAs1hi2PiD2VyKAJXlRu3yNHAsAAt3+Ub0DUVtllxb9
P87k23wARXYGL1QU8dhcZbmF0xjzSzId6ZbOaXrNsCtAZNLTfmdfw/hFXUlYOP5vSTGuUoduCmGK
mn7qt7Xs/mukVMPqi2cCDEhG4w0qJ2oXnAo0AtKYuja0VB+pTtIG65Pd302+yMVUY8+sgKf77LGd
noeuoOxuuvAVFT25iccmL05mAZgKup5RyCZz0wCfL22pxEY5cCM7hRCbFjoG7MRKM48+9HnPIogh
cOZ/qNP36QpqWl8xVvf4tgRDJQ1Kxpd9eqcJS6qQXvGaS8v/eEK4OJ6Y//GdTdaKQ387ArI1fa1O
7U8Gjet/u9zBlOBfUbSzOylwj73gA2j5410Mn8p7arMlwNYVzd1yafm7Rs34YoH3JcoUMLkAydnI
bLIsSN97Pl/cdf1uyLR3H+mHldx7KYk9UfFxTY8OOxQjxk1xqFshk+9KzQLejdQn5NQkdZftZ2/8
0WUpCYCkfYzYxxXIsqyKmtlO0yjBJ4vzNUgsbtyeYSdVNgtIL6C63CkJbSb8hfnKlWcONowN32VE
htZKg4laLDy+9KtOxbcezJymQ6NMxTbJYhE95DRyYx72RfsTW5GFX06oJ996dSTZu+hLAoHjPvH/
Wg0Tvek7Pjfq0+nsjHACeA2gbry69CD7pgoxKqDmTdTqtesvMLtosSs5fOF5jQt8ues+Bw6XTOpX
ohR8XKaZJIV5aGJJTU3m1eFTr9EXDO9cY41DeMPk0T2zOqggTTh8EoBW9UziLQthdN9hy8h1FZ9e
d/CJbyu+iw97alVAkkQ3yo9D1JOEu+LGMUTLf3trRELoUkSnlIVoO+srf8z02t0wI7FYb6lGR0F7
UNRiSQVKS9M7VLOy2Dhj5SSeClfFwSoCk/2EndxdZW2Lb4S2kNNe1ljEJA5r7THyKJY4Nc8H/czt
2y5EnDXpHTMAxzTORRXGQBkwoVOt1sARacTGSxBKnFQPZ+EmjUjHC0Fnfw87DgBi2AXpqfMWkbb3
MUzw4LAEY5TCclkhcw9C8Yz6+8X+iRu92z2xuOmQ5yGvMtRCNmcRnZNqF8YBnqaLPPbPoTuT7Bf4
AoxI0uPeQgHXtlj/alTTTKpd/y2SxP4z4MkWvVvah+KCINMlN4MYH1Xp0yXozwBoRQaFh3Zmjkhe
IA8Hy/ygf29zACKYfDpQi4g/Bt69qAU9UnP1bpvfIuRF1DLY2vWKRw2Wm6Yjmzqa6MXwM6eWNtmE
sj7z1VZ2ypHIn+ZpyxRlvMOv91oFB8YpZ2ZkBaug7/8GGpWFoedOOVYCxuxBZ3YisiUr94zPfiBC
mBfflu6HSnmzIAWZSLsojI6VY/i/3+uADVGGJkWwXgGNwvnDxaIeFPArb7ft3tzFobSCifJFKwAC
re5BOkPMkX8dRpIt67DbZno5vZY8iXfezVfyVskuNSNxiPNDW+qhGn6zH/QxpIgnpzt5iXiD4s5w
lLBH3fpwxVOdlBFNwTfIgoota/HYeiYV1PSa1B0dG4/ZRHCMjI3DkDQgrv0HjVXypHKIri1gYE6U
gzr2SJfAgm1CY+tW3UkaypU7mlqnbmHBJyMrA0bpyjQsaNQtlV+jlkywwOlKDMQKOTODwVuw04yk
6NZfBzGAqKb0/XUU6HimnnCbLf6qmBpQEkdFBE2rKIoZsknbSdbI3kTZbreMFBHXeEqlEQoFYKML
RK2CLJTPKVL5VUup1HRHQVOZPqXG2uzEXeUKxUgGvmcMBfk18CcbY4PwChETN/rGpNFrIk3I1koM
HKA5R3zeQ+/cYeqC20xTEDgwZpIDPV/eDNSmVaRUmSXYVRvFXw/EeRD35clIpUGhHF+l+BGO4UrI
yCaRIX6CNtmBnJElbUpcezYDQIvkb5JGvxFWanRtigaJMars/WbRYpOOudNIdCq3PZijipTvx3PF
HjM/5FWA6CnXnviY1I1zMwLn9oSja9o/7qXVtiz3zFSjJKZCpageF+D6B1Cyksig9uXOjIhlUgbx
sZCVgiS9djfBx8LJvgHm92bTi4XnYvFFg43M4oLHfBzDePuCW74gyhgHXAWOjFntwpVz64qyFqBP
fUbFq2yBDOxl5cLvemezGCXOM+LeldE1u8J6XlpFa0gC9CU2IlKTmmio3lbueA/4k2yqS3LqMkQM
C0Liv0nZZ0ol/PUfy2TfxvF73HQvkEcSICfaePcyTF5yFcxGpXPGai+yFWN4C1G0jUp/z4afX7nO
4zuBpATxozDrOkICySAggCfBfK2uJwfpwgkRvwJlVr0o5XgMJ+Cgfod71OPQEVajsnE4NuCtTLMW
acFQ0XhybFSKh5rVMMPv767dzj/1yXNUmUG8SQHsa/bprMhzjtvNVXqtXWIPoD61EHKXBwMWhfc2
5ZSVvyDsHWwp23Z+1LVA6om9eo/oBNWXvPAAL9tt4e/2wvTlwy1PUtKPaUxUiGT0vJ6rk/uDxbPD
vyoh4SYKKaXYldh9OGsdMOMPoNPffe66lMfnmadjsvzBsax2JmMmnOSe8chQX6jL9CYGCESV+Dbe
mIVOKTdX3GXm5xzsNIyt0JfUgwUoY6oupN0YrzQjDPWpi8Vxlbj7p1rTp51A9LO2axrCGYmWlnHl
yJHHuF689njVq3rfO3ryQd006g9LeqNIPVI3qpXIjWQmK9Uy+UrbIvzcRsQSg/TxQMik/9zVWx4Y
hFOHJX+1mL1P+7YJr6AcoGtqbyuWyBNufZjTafCU0czZc0Hz16d46wUTT02vBwXy3YKvOVL44v89
7FbfIdUBGyqcYaO0m9aO7ky54z4H2jR71edXFoFgnxDmOLiaQNI97qk02LuEhGvk//mDyiyCY5Z0
3tx/dK3BHM4r1buLgKN76nvonoNiLwD9d1CWgQy5KOOgL8FzF8HjRVYSvDhqoriLsWAXYpDEab0U
U5BM3AVg2IKXjA3/c+z1YM083sD2sRCgo+CD3pcPZbi9dRSzkLucyv6ium8OT0xsex5EdNG7EkrT
v/Uc8qJNoHxLg9y/LuPYMkyEq8M4Ui/lOuLpvjU0iXa5pAyd1kOwmf4AAhlyJA351uavYzWTY9ic
7cBYpJcb3NBtQl16LdIF3IvZLBKAuK6IzZm9K5Pz7sQUqAs4cbFPBW6QENQMmBMFFTHDi/Wpv+QV
XYtre443TN6NtLbvuokkvzyzBX23HJX+6QLvd8HLeS2l7A+i/NcMvgy0G4a8LTmJRsu6yhYCjuE6
OtHoxN+9NWJCfn2B0b3rCkj+xdBYAYi8e+s0vP1tyL8mGnXe6h7EPkacPOW/s6/s1HC4ncMgzqGA
Dak2zXGuJSibgVEvf9Cy5lHmXo5Kz0ujr7PS11cOg1mb9nJxWfFjekfRu7h9WPaUvEmUBzVI3kyX
JLxk5Fuj1tyAbZ9/tD+ZNKq4Lx3sZ9SI1qGPeZoayQnNo+APQiRRrk5J5zwUu+xgfRaAk6BLrzrC
YCkgf1Xs+tJtoJXkEGYZFs6Z6VYKhbiCpbErkTT7OfRx779R0xh2N6SEUSZWZvr6Ko8c6hpVgf8y
tkOruPBmlgV1lKQ94d/IN/FWtc3Jbvkkqt7KzeKUyK7arF7vEKgEhWsmA/V9iadxFbiQBi+pvKXN
sjELnUeBhDviSfMxZzoUOLtaoVfW01RJFg3O0q2RrVOyBDWUPaJ3GeYKSvxbrxwotfQlXUXbK7UE
xKJSSnY1FsnvCvCjKz8z76LGDWZFBOV8MJszJC8L8vJ8+6AE7WCbSwe1SDNErJ27hVgOdmCwThES
RzhyWXX3LMhhWitDkQiz5KTdLhNN9232oh2oZzaalnlAUQYm+k/NNeIkoXdEX5H7AeZGsyjZwwGA
q1dUdlsjGBJX7TBBkhqd+8LMlPwesIyxGDFkXtICBaRjD6PROGc9NqAG3scBiizRoToo2xd+BXBM
r8SAUR7kbhLpZJxuWE0UBkQFmLZ8aNpvr2YcRdF6vNzBvP9K2fFnEZT9fAeiJuhQn2WYUP/O6Jbv
HUjbpj8Q5yMecZEaTEWsAmhRvIKbMaFai0g5lAiF6tLQOUgTuzrjWCR3kIYfGbS1lX1xPly8wpJ6
acyiNZ7b6A3onTsXP3emsTMIMmn1cIXtMKtU9QvDVfy6s57Ee/6rDkNW2RQ9S0nUeVOjb61aWjHS
92iZbFGZUoHjI3HzRD0BAgG69AQEzfhLHdydHdPM4MvABc2K/5+9juy4hN7Z8XCgQn4/ymWgC14E
AaIdZgYpDny+enEGGZEjSQStviyj+dF7wrIJ0a7LrGcqsNUGpCf/SLCpH/G+1ZeVA82mkMCiG6c6
SwdUOlmpjW/2B20DwdGXdYmRfshQQpBxTWOn7zNSEABOIHY6etmHkGpWH5lT2ZCJZYuMFOZglIfQ
YjITi7jYqwmRlz4jq3SfVDOPDDKmUTUGsy4X5/Yo5rOXAAv8EIANaepz2CVK+mcn8aQDbHXYlakR
qtfJLY25scZsgcDpO4rVEtzhOgm/5sP1iKk1xCI+ROFU5x2ZbH4oCElPljNz7Wc7A6gHUCoGT4+V
VEYpb3uilqS00pulxGs/Ks1HhXbdy+CRWW4SisWwVxlD7DQc/+n7tZ4OFFXhIu5nmQ4oTvAs04uY
voYaOJZVI4EpmOhCkqHNUUcxid4nJPaX9eIqPdT+Yr1mNBomZ+J2yHh1PHUZPDRrv7fPzjfxO9uQ
+zvdWAELrzjAq0AZZ16mIW8XhD9ZaWHyIf8vJnQI2NyQmq+dZqqMgxnSDu2EB/t5WaThzIDZYDNE
gwGtYHbYt1N4aGwtSneqFyv5uAF74TjH8VleHYrkYBQkCAFlmmkphB4BFCRqmo173V8H2X6TKvzs
ccx8p87poskNkCGGKM+mOThEbs0xvyrVk6lgCBs40dpkh9LrWsXeQ+eR/z4OVmxJe27h8WoHCllx
t+Yqe2m2ebH0CX7K6WiwyN3MhlbUAIFES8EXcYVR63A9e5Xu09MDXHbKIwIbEHa/Nb8TCTskb3hp
KI9PbFPiBwURw3LD2FSAPr0w5W8a+9BxTU+V5uFe+TbridVdCtWlnSjbGlr2V5Pywn3kPcOqdusr
lCMkvBI+o1kdCgZG04XMLVO8ha9jto6VSrZdbDlA9/di7Ei/XbfE0G9q1F4kHbB7SQr7ir2aVfE5
/tPTFX+h1p8ndMcfcA8UdiHUQ1ermPd8Hl7otBDbfREKmR3HnXWtjvoRNiwvguBlOe4WXsXnJ0xt
jpMxkpwUBE5KAAK2rPz1ShCuyRpG/Nm4Eo21fMFKNBQI7Hz5vexyH2B7c2htzdveL1t63kPFbCLC
3V8bSTB6N0k3Nn603qO4p2kjVr/uKJ36UwfyQP0voPhJ04WF08EKok9zH5WKrw13hVdaREpqRHoJ
gIXbUxBX8PMlLAH7vxuc/KayWzffnlYtj6KQvLfnV4RmXtMhraSLej/3YJcNl9vUQ5DlHJSzfQfj
f15EMiw4aRPg4LTB4KfKl1nm8DtQpsmR9+GRYKfTD1u4L6jpZVdCZiTpTGcPCZBIcxZoKNnV7DU1
Jg5PoAjSJoEnPs5C+k6wEZc3UHZ9dsOb1a/YvKpgqL+YRSnF94UeEld8rc/0QnyJz7PTHQkw1web
lyPOpP40NJAngeJDuGbXgRwfEXHFBlejaPCr32GSeqra8z4KFT27/1WOatYbqn9eRut1Q7mA9T+2
PO5B6lUy84aVOh8Ha4nt9PxbfcWbTUQoWqgR52uuutzzWYOOtckmBo6MhcUyVjp2/035rNVDzpy6
UDLmR2V8laO+wZ0uoRZldbY6swNMO3ZdocD9SGCf8+5nmBCqeClN+us5d1DPQKP8vULzcJdG1c1p
J9dhVM0Opr7IxTFb0kWYM8gBazHv8G7jLKUCtS+br/A4vnhoxJG3A7nLVoO0gV1uUO7xEHsEFyRb
WABNCxsbpstgAhZqRZyFfrsxr9UVTpgBFNPCgqEK92rgQGX/dPVYeneHw6+ZMHC5R5tRYDfdpT4x
r4lsJWUWHna3ibY2J3wn0ItfH9uKoT7Gq1VoRw/jTN03HuUTuntxDSr8QYDwYbgRJWIL5FusQsNc
2Alq6z3OLbZ5JYlTGaUAIMRNf2DxiefFgqK/N65yMjKg8tfEOH/knSKsdeIyAdfddH/qD2M/1pKZ
6UyPL4IOE7rhcuf0vny6+qcfjjY30b9zxlejeel4t4u6ixCIp4Lyc/e5bLmwVbDn3LDjoD+SVYWB
CcCNcuR88T0vVr8p9AuxpLcJZkGqZAj5+9lcynBNOcVTUWDtfyF1MM5rpbdVRkqvdmZn6iA8BZsd
JV5BNLmVRSaSC602HPuM9Ip0R3w2v+SkaApR6p786Zwwd7SCLm8C/PezZ3VdIdVQCgQFiYMNPRv4
GNg5zpbk/Kon+HTrmeEZ+FXV8EqrX9FSEFPgOS+/BMJTfZSKBHxITW9NTQobEZlBh7iLAav7Q4hs
pr/80gjcWMw6jOP8IOKsozoYEZf0bDDwDGmAoqyEY06vwVLappG4XJYQUlRzeYSQoFuAjPt9RirW
lLUHbTsslUjd/9y7xo3qif0d/V9B7y8ZMYOfrRCgdDHfVh7unNq8lDW/Cyg3d6nTOYFI8sdEXr/d
a9sZDbm4Dm1LBYVAPLnPnsCg3k6Dq4CzvzggkUwwm7LG4n0F5ma9vobBXz68llA4S/gL3xwLXrdm
4tTsmJVR+cr+Alp37CmqZticzHcLv6I8G1L8lQymOdb3ssntSnGMAbtNLlnbPFGXhbi1q4Xmr++M
brI0xbX1AilQHiKSrBgSDuS3cytmZgHsOFWlfIiszNlSkslCHUkzkFxiuHE1WgrZfnrssm85IsuS
kipWskE3+9LUfqrtlSoCkDFtWyMDWu6npATPY2etGgRLh32s84UiwtRI7OFEedW621TEYUjR8cid
8ORZkhWs+45MAghwR7KCpAfxdr2gKteU3zYgurOlbF8m3Dk9UZYD6UFq2F8Qz+MNFAOK9gl0JK7U
iAKCGDDE089k/7NRJatVKAE3TzC+T1ZqjlyVu59PHQeUPMvUQQHG+NQqOCp9wucEx61fz9v79Ze0
yYSjDkW9zaKiTuDtK7b3ziVOTIE5RJVcUV3SLqIpStpohtwP0LYOHkmHxDEqZS0VOWdthnM+WUEa
Th+fzHZiQMIzT18A1yQgUrq7O7aCvw4eAPsFxXJzaD/DPexY4xdWLIjYthjkL3P9V6S7MYkIuSAB
uvIBP8Thd2K7OYiB6fgOZoVmbTq/ti6BRFBVhPhdudoMWH4T1zdbvwZfbWozug6gyw9aTjHgq79T
50asicrycwvibplCrFVXV8ZveZUAx2etRGkPu73so7qwGz1LpnwsGg22z/Zw6IQ+E/fdKEkcEj7L
Fcf9ScUpW/pXtoy4pcLCEbzeRVBdXB7F6Gq5pP5mpvL4LKhZE/5NUNKv5ONGjQ1UvMOabL4wrnK7
50yHo9NWRFk4lYKGeVMP84k8jW+ozKixh5T21AaAz7C4Ea/AVj/4jLgANdA0eechvEQ5FWv0JlZq
thhOftLxjYkYq42Z9u6M4JaVzP37lAK9PjDp84hAg4k94P6D5DXyB/NLnoJOhuiOoze9P4cwU1Nt
kh0UWwL5s8Axh0EQBNv8Ib/b4HyfLdnqQYze7G97xoPjAaIZuAofYXFdLc3yNMyRju3Xgp8FFAqP
dZ35Dw9KkPYLoNoMkGkAzLxVr7mktodwnMslJ1ql0ZlDhnP3PdD7F8nxV6PuGsc4VZPhpiqDqc+b
j8XF3NLbi4pCTs/QzPQBMCwwiP5/wwWfYCH9hEzOXO04IWmagZQTeL30o+cjAQtE5C7dXjDUDGXm
77uGxTR3tmws6vx1tsPfa9zIpaUB7Db+R+Furh3kZbK/lYo9RYmt9H5iBIsDmnuBE9tKpzPWFOWm
iETfY5+WadRzLv4xbEugzRstFnG2UJ4IKZsv/0U337YYKLR2TXlgmLRoBGoAaPFba1OO+omMugfx
ENsIfUNM4WfZSYtpcHSzeIWTKLRe/CHeYuUp5mYhZYcW8pxjFsooI8HJKZ0hrKJ+ukhg6lJjriEA
Y8c2liVNGIESNDupxQKcS9zC6Ql53Cpv3h/N/NRNG/AoqnoXA/DfbuGYqqdNC0qUG4ThFPtj/Gjh
lDHEsxBc17PVqIfkpwrRk1Onqz0jh+LOr1/mOt+CpXJ3RT8Z1k/5NaaMsdID9+UPOUlglfe2Urig
FNcbxjur0AleM1BtjpjHwvMMcTkQJMHEg0qDMfgRYZJmWyl4Z+LoXhBdx/NPJLrWH9lOt+iX9Ndb
BwfKUB4Ltmsd/WNMgh0ggvewmtAFjtLQ6TCKiNDnjCzyErklssf9cuHtfQ3K4MnthbrR/lsbgSzm
cC1cet295eRLGwfZvXzA81WIqyc2JmrXtkGlblTymbXUCjlsSSd3ILw0H2bHla4IbOlTGM7ay4k4
wtkrL6/oJhV2+30Iz0o2EfxUFAHHXA4Tkr8mM2ZRPHvoja2vU9w6qFr440Go6OpuvTzPwZ6o5mf1
2JunlbfBxDgxiSgqp/rhqF287ovf9DUWPDsLYCRP2J5CiccmlGuPVxiZDcSQm7kypYGvnKUXLhIL
g5JzdA8pZxVOx68Nez92Fk+SLKbaRvNBx3zJ7sLPTE5e6WTrMupztd27r2RSuVkfG73UkDizOFqk
lf9xxe5tWByJ9Pc01awgI0IRYFYzpyd6YWyglVitQgcQEsiOzHcaf91fwsDmHeQXLQJLy7UGTIeJ
WtzqAEGpIKQ42xFJjtKjdXvZfhOdRTWPDrERghd/QESHifutnXPvBhyeXIH7iGkSPp87q+ttQPG5
YIXpBlCelWWhQNHoAhWvplyPgZzb1ssfeYW5tLe4YBUVkHQ94XScsivALQRCZd1BIYZ9kT690uOP
kgQjPidALOi244ZhwXknGtBAJX9c30d/SZiK+OoJFySumm3wS6ks988vwQX3iZ1j7I5no/4BpZ3D
36dtEgVsn2H6VQCHeV/978ZdorF7mmL+6yU/IemhifMtaQlYz7JWMkM61rtwnvJb01EtTBZWsPv1
abJsj0NFdOM6R7JDaaBKEu2aqAc28hAcsem8xWkKzaEP5hJn6DN5kvDIew0Y1UCe3UD2j+8aJC+J
A6Zox5gW2Yjmwu6Jsukv0ht7sOCjZ77ZUSbn07s12JbPCVI4fZ799qtDD6+pKTEKkcZN67iRWGc2
rOKRhiiD8XBtgZfacLDZvjmG2y5kzD6bTnWUsOxDrCeww3zX81Ki4HnuWXXkgdIfFXmemFJbuZu8
uyezrndXGWapKvgAYieJVY3oB5YtICyuVOBGw5S4+NEOpAyx2Ax1tzyBt5BOCR21RjEhsgqJLqi1
FkezuhUko7kX3pRbk4dPG/bTx7QvHW+ovyN5eV1RitMBse/NSiQKtAOsLngDKW5VPJhb/yI1Wu0V
3n9R6CxKc4IhreHgQkW6W9fAf3k2c1HVTIG1I5jGY8YSRuCmCzkSWRDxRNIJdZzmlnC5un32Qi8B
HUMARyehcgZyaxyOeftmhpqlLADNJ6W8/wKBryKYW7bLu+z9i0OFmocTX9rykyVJqiprOioVAGA4
jDQzRelTdQ4gUViaZPSrnG6FY2a6kT2Iu0VSAL0ekbjt7Z8Y846NB2T4gcTFSP1Lr8+GQAT+OcKW
emGkvLjnfFJvnizniWVoUPVX1Wms3GjUZMs1UJO3ZSYYrr6vO0IZt5Cq4SnY0QeJ7QK3rGyN3p8j
ujUAqKdSa49vWdwuIjfR/z2Kc8jsRoqbUpTqczJH37px7LsC8Ft8Ac49DmazEZEtVuNua41m7JO+
zqlmdOQUcDYYLXv6lEo8Au2d02qVw+J/FCx37oaytuFdX03Ch0Axalh+Y4gi0gjS7My8uwzhtJGK
MM5YdZY6pDu/NrVbrULlWqF2gMFFR3UO1ikjHZz5VpOgxgCTfHqIgTaKS9Onu/Mkbgpf2X7wyUP5
ZTX4YuKVFHITOkXYkvnGPh0V5QvD+XiJV/cKV1uLT/lv1EFsr7ll874oAEmdydplyRX1oMrQVmir
/+Ny7ZlfL6LfeqdWj2OEuHoILoTp3m5XmjCWbZgC07mRjmTAJrJilbaKmCMlwgNq/PNFtuQ0UKnA
NOfI1k58eu6TNlNzgFxm02LihTmKYdDRPScnWU28JaLuNxVbITDxsJEq6EiFUNOcMAax/JzTXt6Y
u9E+IJlJGJi3LLsTL6xuNdNzk652NO0JR9vbjXOMkrye67P1zNKUoNJOsFHREnx90x+3N8Uv5QJ+
jVrNHSw/sw3XrIEURS3UCxf1ycpCHVUge4/C6gVnKyAc89kaXVyDLYLEtaM9+r0McW3DG2mY/Ijg
FUhBehezzRgSfvYDzcuTn1GkfBZfUN4aC9zyVmeXhEHOf96WTad9Cd0j4g9yVOlCU4IMuJJKpHLE
objiIsQUNbwOCuVSZb+Xsz96WblFddmlC+oklSX5hKFT0BEb3TR9xMz60URQS1ogHrz5WDbXKsro
qsc36gB60IWx9exW/S9vdANGBVjzmkRpLYvmsru9pTst7R6RUgf8o80krurj36vQ6nvIsATnRr8o
nAsN46n9gHTBYTpCJO8THry4f5KvAMF8pQ63xn6eANFolb9ODNgu5ykPK6oydFrR2zU16pPJi5bJ
f9L8DWCyMn85qeEVfpiuqdt7oupQudTszalKwhmgVd9teIwss9ZmeGE3ckEFcks7/fy7ShocM38T
cICyug6AMBJ3k15Q5Johr4g8Erx8JNKLrkqQNHnLBIzgT96dTiESjFjq0VPbAZhvdH4Xz6s4JJmp
oFCf/1jNZpwgXy00hEDpBfxpRs0Y697Gg7jARXII7tXE2vwQAyD5bVJeabo1SKoeuomHvBsE3t9e
btmuzRs7o3oFHLIufK9GYNN2LrgWjBsteLmTugQLrlCC9EM1kkVi+UyrJYZBkOemGjRgCddwDlKU
M15E9hhd8S6BIUcBPFbNAqqnDYWJeyUzydXyhBd+I0SfF6IrJf8BkTfqjs/HjkrxEmrGA9BQkiHJ
7hxRkd59s5frs0/OrskBdosAxyFi/mhUeN4yFiEVEL4/BKgqKR4/9YC0AuEXPVB3t3r8dL7YdaVr
s2dhe87ELOvw2pEt9K3CpQiXMvpgYcu2PwDHl6haIF+tbdP8B9xl6JI7jzxC8OSxajOiB3mMMl3n
u67jUpeXAv/rejDWGpRwORzxP/iCTVTa9BvmCJpkAiS4Bx2xP7GwnYcm6Dj75i4XIlyNm3+RLVdP
E77/Jb/Fl7xktm2qR9lhpUQgScSp6iypxSNR9tNSk8RxgiI66qoPiVZrrxWIQJT60F2PFVeVk+My
qpvbLN6FI8hAZepUhnFvDi5F5MRHBywu0JeC0dzj6SFpzxrXM/f7fFbB/X61vO7nwg0/5qwsNVGL
RBGYH8nm8mmUFOwkbZNBHbqXW6YN3YNYYAHzu3VrRcC4/a7DrBlm5GhuEY5mGOTzY5kFhlzAH8PH
GgaS2EDRagUZxfqjvMrNO7/N05+8+EQsIdrSejdcow7yP34s3cDBngxPFT/rD78ogXCbDSmx80Ps
w4qnXlDZBip5GSPWP1/OQsjnefBcg52JsmaZDk5aVXGSSRYI74IwgwJ97zeZCMxEekPKSciTid2i
nyyc3vSEwS40qHelRYfiLzgYVUnBL0Pp4wnu2WAyHMOIKilcBPZZi4rNTSPFLIkApyhlXLXPS4n9
3bOc6D5ZISAevOEbPDXmkhzeKTtjUpDe1j3biRiZesHKHajii+SCsc16ULF3Auygx2964e2nIfL/
J33dACJwxygKkS9QeSdiALebb9JRF4swmVuj5mnaQVpDHn0W5H5qaef5P+PP/iv0KAhsYUpyLkL6
AV3TfSypHRRLaI5gBN4ET2Rf33V3RSWHw+EiKgFHgtpqJKdLxVZgqeQR7XhLJ2WrVM8xUmYz2fAN
2GEBD/NZeAdJZ4DoYJneTambbZ8shTT0rd9wgjZOvOe9yLKKfVlNq9qOXd22u9MW5ojGUpwjA5wP
r7rC21m5FDZKuYoIG25PUcDPkbUkqiGpQ3u0/1f5rh5+zZH2q7kGQ5bQi23nALtST9EjTfES/s1J
iQZ0f/7qbTYI/88m3bUb9+CLh23ndyKcQzwKRNcL/nAmnT480ATPj0zktsgw4se8bDZZMzy8Knv4
EhG2psVjyFAAKa8by+5EMa5k9HNb3P+aANF5aBJV4koyZPwNN9NVb56ai4TolSoOf2Ed5BLRdOfH
i/a7+u2Kz8eRT3J/S1yMTaCcL5qKB2dS5GocMq3ZwsLkp7tPBvMcTkYi34ur2fiDxfNUn6nkoL0f
6GwCB6iWxulQF3txD9f3vY6hKQV9A4c82u2v5CsEkAQLxcLLTJ+WaKyBxf8mzcDjBH9AAeWkEj5E
Gp/WYTWvU3JKl9KUr/86k4HPwoi2srFKktF1Hy/kZ9TDmP8fgjUptaY6A2Lb1l7VWHDO5wB4GVpJ
9CWpliExNTkxO70A6EelYZdcvCizwn9fpdITr8BULHgXm3Lmw8zfBN+abCoKQpxVbguW6ZGsR4e1
EJ3QUjCOmE54mWvUVTGqDxnw/JQfAVd4itU/48OB5aFtFuVKdwy8VcTar3xIfjg/c9hC9jUzXbAY
iI6zGKXy9gL10dVtNHll6hvio6v5TEqToKYzE80RTHhvsbyrzcP8CMV5d2ArzdGpqWXf3TjaEdO9
LAk4MTEfSefr9smL7FEBip6WF3J+vPpQTFtsyneEqna+aV/gGfOmZG69avDENVHcrICeKZ1JYkR6
lZJraRQVEEUkMd4vvBzk+vlW/wsSQsKQroOO1X2D6TEkBZdvBCW+mrmmZWfr92WLOhVgO0Slkci9
7roCiSnNdOAnux4ljJiCws1mV9dA+jGfVbRIIYSpgB1oqSpqR5wDhS/AnFgMOqyW31Jc4O1rWqfZ
sHgzcaw3+UzptbdmNsrCFTIeUX4D9Z1ixX+hhI339/Y7h7AuiRq81sITpP76t/DqxSqfwIWlAhcG
l6ztQnAPVh0kSRi45y+yodaBgOIqHcIKcqcX22KZyl7YSur/McZqux2lP/7OWC/92G4V/W5k+sAV
SoOvmAulA4ha6OVlfVx+Ku58TwdF8DOFrGNCn0nVa8Imne9WboapEuoAy9ryr3kJMLb7xOTnd/Q7
dbB9XKKDzwd+fsVUpU4BSRksdPvSDRHscoyMAuU+8m4dGkXeMwpsAOX78N+VPvgpjHvbL5C94izL
0Ffk9ePiyHgw9t+nxHoU8SbgWelcq8aZmk+OfYx6UViu5IsnVujylGkLoX2K8gxwFb0wbMtRmDTD
2zAnvNYyaFGEzzNrvI+7bECA1FagISuF+j/1XHnliglYks7uy9jeLY0XE4P0V3Zif4E+26i/iee1
zYS5L2XJcusgrB8Wt3JQQO3HBylYX871mvTB/87jYFdbvMBi3pX+7fJjJTDFr/4EotO4PCgeKnAW
2BTUUyr30A4nyFJPhC3KqnhSIiy9GCxgFX95wK9u6j0trUY2Z8tjdR/+ys5zK4tz2uWpMgoBIRz5
3+xHczf96pKpD3lr0GpNtiW4Sy4LdERCaQHd5ehVmQgMirEI031nlJusg/Gp7a/UOZLTYpBGF4fJ
YZKKE2FLN4osfstWmUPNXbczWZhUayK2ALY7k+Laj+P61KaEPHtE2bvOz9XoO88KWXBt+QLEsQrG
U1rT12wEuy5rfmv96ZaUbcZ57HzPlUwGyoIC2Rpg0G0UiZoee3NFOZofjJDdeKpckCGrKP+p1jkY
8QLGgD76fmxUk4lDmcvaGplmhjtR808ErNS7srzEG6WFyqdB40Z5cjdMhwuJG/miGNzkv6oiu5Jq
oot2ACvZ7hQXedsgEszVQ7llAq3VdILAmej+Hd2vMH3UDi2gN7QTm7XxYm57os7AqR7FlTWX1ddb
aycbpeEhWHQiBYdxdboZy57BvmXsntHnkPCc06jZ2Nd8X5ArYX61z87mJ+8E3/uAeAQfc6RmLBsk
CQ+qLm1ifGucVJnjYwwf4sXWWY5Q73mW21EQYa9SJzD7eizvmEPLNC+ZV3rM2covMdBzrZ/M7mLd
32RGpDqFyAo8630l5apKJ5y7YuuYRauXa9t3Dic/7MUv45VUPS0/TYqDMb9oWyC2/Pl+AAb9/TDC
GIPQdcdHbxrJ7GoDgeG0vDYictaIx5XEjbTPZUmu3Aptt8bycw9Su/lb9e8/2jrhJmgyt17ZYl9V
oZsDbu5GbNrekqDNaM2tjRbG+Jd9CIfxxFIJm1/kG8beDY0QP/Ns3lcssWW0x5grS3JsCmHcEpGV
DaOBAbKzGK1B88JQ+i4DUYGWtOJO4lg9pynjLDC8aNqmh3KV31zgYMPtSinnN8WBgWANYjWem4F3
jjfknpxH2NwlDthQFNv1YYMOngug0BsygJNSViXBy5WWza9M7a+4l218wXA0oKzEwuckGeGbdmSe
EBzrpXof9whty+oQac2AsRLip/OeDE6NZKTjhaEV2NRfZfnsW3MmlCdEaahlpwU/jYNB+Q/UMJ/0
ai9zG1ElUTBKaYIctYx64R1PxfrYCU2TY91tSVjfJG85zFBx9EHyKy7MJY6dKTbVkrH2o3gcKnDl
9m7D19dIgzo1Of8X4cEiyLQaE2ZpBicgwnaLczhTvJlxRI9gZupObcSRGg7EqPY3VbkF0wkd4U/8
DEitRxdFCWA4abdI/plK5Ki/TTM+GB1FKz4viYyvraG2AvidPaKhmtQyq+inNN6f/Ujs6gLxl2aK
BepfE/NqMm3kyNWunemN3kHKPmMVsfmJUQFgVFP0rmZrAv10fjg0YkJMb7rdAAexjWxFCKw6bHyF
mSGi9pI5ivGyyfodscRbc1QQIdOu8rzWSb6N4ofCcx8/m/LXrVZV4Ciwamqd1PD7zpVhcFP9PycY
j9Mzn7KYpGYejIVjGHboeSY8fGp1EjR4hLLJPQbtKhJVdmZrcTOkdfPlWv+ul/n1VMPqsem3e/da
PN3y/Ixa7pwsL87sdMuCD/YmJC7LawkxpR1wN2OJh7fECrsw/7sSYpBY6rxaAlGjygLnsfBDJSRB
FGWpTuJkiyHMI2/tLc4nqIbwLs9Y1G9aNxqegIIpTcM7yuYGnI6knxmKb56t59vY60H6OYDh6e/1
O4MEtoBR1k+YVyL+otuJxYfDt+8MBWRUeu76E2+Ct7iJjXPooA+FHvx018q0hpcVZF4fgokTdT/I
l9lxRS4i+ZDfutBPR54PEatATUM2wfHak0Nf9nzcOUXVmjrB8G7yh2EzjR7y5J3+7tenVKL/6I6T
rrv3sBRgBsO8qfJSR9WSJqg8zgF8YkGtK4EfbW+6HfLT5z0yGQYECOzTyLAMdcUIqgrWccPFkt/j
Io/18vIhOEor0CLA0ujcLChCeblrqNzP895gjMztdKNdGu3TG5rVj8XcSQcBqyb65j5zDW6WaNqR
3hoZYwxtrOT+e3TgAkwJ05v62xGwrTov+GaiPJZ9gI4X7qgKmNwgA0mVamJMEzndXD2o3+ZslJpP
UpkfpLKp/awgzQZk0IO9Z3zGEQkXgKDVFn+C6gTBmHeFKEqZnA2AyHfq6M5QzE0dmWcgBo7NrV/r
rWc0NtpXsUVsng2AyY6yBLAud25r9VOTqiwSZTt/sNjCzItGdGriKxwjjB1XyS5OGEwRyPl9hBZy
INNJHjLMdW3GWO5ZpgkJ2nL4k72R5tWJXZF5dP28fkNv2NZIcfQwUyAXWKSr8Je8E1ogTKdnOoVe
0IruERjVjes3YpWJHNUfNiPMTPOq6Xlmzc5QIl+pOe71/oOxZJM/G3IzjUCkYRVJdst00GnXj2to
fk46w7XcndNne9C4bLKA5Dtn4y5Je96hPcHfMWhJGOlWCZJXspzS1E0hmf/Qq45wcv/76t4aXUbd
vBmhD7x4zNai6lByW4cXcUFipO4iDdzRCRyxtdTn+tqMsxoBdJa5j7ZqsQlIupG294ZJxE+tFKxa
+xRLmbCY9Yix60UuW0IdSEZlPW9wQ1WsDY1alX/sJvUMjTd2Bhloa9vp9tbgLlOI3YzZBsdKmIek
GPLQ+FsFoXn1r8Om1xW+6l1OnQAuC+LFBFEGc+yzcz3so+6JPHLCDdiBYNYDMMne28cj7QB4Iaxy
/9ISHhNfA3RX9eTjuUgH24X8sVOceKzGT4znxxg0SJVKhhjbqETKj5Tq7kfRcIJrQOw9CGah9710
hHffK38q9ty9MEyIvwXsDXLObWishZZLZffjKo6taTaBTjjVIqg2nASE4miM8I0jwpiA4alxSYwV
qSF4JJnjB7vlEvMYjVbLZAnfgXqSlmL/HQnpYTYefpdkof0ggGj67Ayg4gBGgDYtmie5FJenmJvD
LKevg44LtFSc82h7+qxV5UnWCTG38BXZ3pLMXb4WmgiEEknAa06yTrd5Y8vrvDoi/skBQsuzbkcw
q4Xj6tN+2ek087a15gZeGdtko8KnLdx5fyxwx7hbvHil6Uq7DmPkMlwpA/RDDwcPqLyCWbGKNbuz
W8Rr42rjxUKfCOo+MeYicNicz26cIAUzl3SB0wgMZBKFnF1aeY5Dtg8EMvwjxTMAUmNmUoSHiGSh
2IbdVGxPkGuWO4Pp42fRmHTPqRP/uJCCPfLHcz5dVdkPmKR13YIhl9gcMTs3IeWtuQWmbfSevnBm
QkD/oON9o7OWtLWNESsoRLjH/SlXZoXlLRQUJjYxiTYJUm2Nx9DHM/P4V+iwDROAZc17zL2l+nII
tX5gyHH1h1v3uD1F3W8QCFw8eAaO49eI5XsCiW4ZLszy2e0ADwWFWGEy64VjprYEhE0ya6/pZFCJ
4lJsUhs8OAZGpSS4y+7KfBX6ImqioctwfulXTx63TVDUFOA7ig2i0qi8FrKdzbUDohDDc5gZoKHi
V2BsET+Bj5UbRY8/uXgRcgTEWiNx2uJqUECnjXu2uNJxyKkZgXTZcaTSRE/PvpM+rGDTYNLLyrA/
7+V2yTD3NvZlywDgNO7TqSAPf3pwaxy/KqevJu2jlyQ38P63utTILaxz9jgOqBaKKeAkR8xQMkqQ
3LMoj/y6H9sUr7bObUwmrtMYGP+r+Y16v4Q+5OyTCTR+kVavg/BcvB5IQqc0nfb1exwD0S5t9jCN
IAH9RrQ0RCeOpeECpWcHMH1DeIMgwmJKZuG8afHnkPpvRAE0cAYGFEkz175B1ZIKWw3KulGMqRZK
keE2DKQDPDfrfOWitCT6OZkixVLMNxIdomnvV0CDzqZ+u64pRyY6tOZbSUE3m4J67EV/nWvCxW8x
KwL9YyUnPpVhNyPLPrsouE6baWb6bw8rIViEzOLsYdu31H/Q3WoZ0UxmXwmqLgmuBx0kb+c5CaEQ
V24UvE+2tLVje5R6GerszdKGvl+BxfPy/0PzislhTWIY5RUywdOi5p9qKWfuDWZ1brZPEfDlA8S0
XkSsW0XN6Xb4dtz2KJkcinVRX+DG0IR05Jho9c2v4BuIhD4ktnhU00+/tu0yhfH9w0+nuJQXrbvN
hBASsEVIrAaKSUfjKJDcilEdqh9aVsTFtDicgqlYY+t9+z1dXm7Xk4bip3tKNEBkE48AnxYC8Jgj
E9HJ4dTlFUXK7IgiConkD6wnnMw6o62LW1GXn5cDgQm4jv3sEd+OqimB7ZdCsUi02mSGPLo/d+Fy
8wePjEYld2+iEbrNoWtcAReQz5Ef05/Ih3jScdKgcideS9/ypl2GfSASSHiUmarY1f5DkS5oohjx
UWOxtM4yxH4GKhWLvL+2+Me5knSu0S1IMq3yVRKWZ7TK4EnJ1rdwGlYoNqKtkc6i+HBzgbxbJPq8
atHLNEOIDIgjAtGYj3iCJeZusAm4Lr4b78g63uye0w5aLqY0KSH65UfyHNtmQx5dEcKDKxehl+7h
UkbnHY7syLyL7l0gTJv6XZTWTJnVhcxc9hi53/Zo4/LiJ1yercJUCF6rZZf52XLuet27NhrvfMxo
xi4uFC/BktjDt3QpCD/yTuvAYQu/Fpr0rQE71YldsRqGUc91twx3voWvISber1mgV9Q6VxFzVSFm
NFaIffjoW9DyOENrUfahfM/oE3hYIht7yaXyn2/HSDODvqDTt4XIG3k9kkki5meuC7sAi1syP+Z1
x7zLclq/GPnWSOiDf5x0LipjYrvt+ijZF0lvkWbznqCp967rwlF0VoegZGF+HdOIt+s5ArFuUZOr
jszk/uALd7lVI/PtfDub+Z6zHp6vKQXf4ivfYNR7bt+f+8isQO7r5+Xcw+Y1gLmvLqkArCcf6urH
BhOQ89kGU/0kR7Ed4jrwTpwXi0EfGL5Q98GhmnSocYj3/CbhV0j65i9Q/PvyEdFitl68aSozB552
TJjtVeMo1V8QEGrC8LCEw24004NwQl9zvccLBLM061l+HUMigGxoWAkXbjY7oPftrpVLZ5YdANvq
IM/OboqNw7J+sps1jaJlRNP6PV5IGBQrEqOLbtrkDw9U3DRs9HgxYZG1NtQzj0YpeoAKJq5yXaMT
qEb7QBFyt2EDPXEIiLpuxxIiNB+/cvSZr2U1qWNs8e/yx2y7fV4mesh03AxwTQErZGETFTvmV3vc
Qd+qPWWW1liK6NivjtpnX57z+m12dVmelN+pimnF4p0oC9YabMQ75NnhiX1bJ8m2doyYm1rutrB7
QSNV3lXxX1v0pH3dkrZ1HDN6risvnwpYqoq3S8l6ewcYPg1xFPQt/cWhrDv/EqUnrDxHioyUBzLM
j0Pku2qUT/eGppD+NYZt0NLMXPA2d/pfPnbDeA2EQ8GCBfZxBLOQuyJKypX8mkJtNV70xT9HJVYh
dGgP5u3oMF9PspYUrRZsxHO9tLI/lP9S5mJLHkqJf2BpuHzwOwO3g8kXIioMDygYJKr8PCOhOPbM
zynzEZSyuSlJGoMo+5GdfYR9WkAJbnYQjHaaWza69nEe0wOJE7H2IsqIV7bad9ORFhyGtfrHebnW
e2oxa3pch6rfSm6KZzum7m8YsgV+JFLto5X52pZdQvvojekq7fUf7KWehJQc69+qDS3yYG8e7bhj
AXKEra2TAM5VCil572H7qO3Irqw73dSWAg8XAGk8CG1Kv9IOIqYTlnpXU+b3CGhdsg4jtqnnaGIU
FMSkuCZr55VwiK3iTNC+OxQ7wh+9KLwBHAqiRLKez1WKygZvtdw+MFktObwBOJCLmHL90ayo8u08
eoWA8uRWSxOSgDWI5navJgud1vKo7eU18PEIfokC/56ofTIbYICV8bC7JP+65tfksaIwLNVRqppX
Ci1PFEg40BtSSfYGtndKv/cZfks20bGILlKddvXvCCYTYyr+36AfcOfh7hFecCNGBAXjiYFAvpIf
yXMbk1L+akcWMFzlRBo+gciyZuQR6j3E56Ea6MzEqIIWivYoWeE62Z87TqAVHYboli6DjbezXTLz
hHb4HHJjGtE0EjrR7uIYWF7DGDwvknVfJZOetoNkXtF2XjEVhZxNEvB9Q0Gha/j4M77d9lTMtd8Q
rCPHy2X5/w5e0TfPPnE5pmRVZEc80ztMW0/Zz9rqKW7cfdBAzg7E3Fiw8YS6RftqavceThyvE1rW
8u/bgq9hUxMjSrIKuc6BmghAZhjUxv5ueociHuNUTd0VKzIQHegd6sL2PrRBmjdRcwSyVRgQ5LxC
T4WI6hnRQ7R3NB+k4vS8+M3HQfIq4vsWgqX9kWY/Y2vppGqe4K0z9p7ibed1c2x6dcWj7GvWZTl9
8mw0paZUantO3KnCd/ymiuJMTKooXSVq3KoSL9DDuyzBETKdqU4YhN9B4vdpNfwZuR5c9OvjcF0U
OxDHRasBxNESftEJjjE5Vnjcfn6dg7qNj2MMN1mb04z4JSbSxgwAQu41lXYREVZ1AGZfLKRtJY6R
LkbVs3UrDQ0dblj9kuYE8zm1QD03z/RXwSsuoLZ0OQUfyszawt5a9hV0SsjbPoNbY2IK7eVjNXqW
cSoqKNjpNC+UAt7FV8YrTAcO64Bklwq3WEC6i1Ihd/sc1d5FHYXNA3Qc2k6NXA/1gFy9jnUJ+ram
JAn2tQdu27GS+T0jPYcS33vm41G+vUbc+uGO/sgY/vZ8YhuEX7RgoVwVgVRBertIorfmH9sYYGOI
XoZw2wrVQ+eAXfh5tfllC3JgVpmY0bNBVVv3ATQAEcrvaueo1CUhkYTQfJq5EcLUVYCW/OyRukxa
6e4LzS7jgOzMc63ncuuyP1Uh5sGAfc7t7eH+BLAF1bJKAd+u/JZigsMa0rhJC6NNjdPq+zacPlSq
ElcHD1aEcXNR/N7YaF2SKVP+ZMEPqXwAiq+MeFHiRPS7mAXyxjLhPKv7d8c6ZEUmO7N80g4U1WIn
QAU+qfwgI5c4+h3hXQ2wjB7eQf10k7COgH1CX2DUvpLyJvAi8jfPgcRbadaUQeofa2AOFrinlwHZ
mgYiGusQg/z3OilfmG+8lGdMJHWconNi/s/yRS+jqDkLxOOH8UNRwQWhGyLNiSI7j2OVev153KLn
frU6q/MgzFJl6kESLkW/SGGztcsHTrnC+KxpCmFE1d1xwg8xqo36LqEAhlZ1LsasFjJDx8LnH8dB
rJ+hXBiAhxVmKoWSYb3JwzqQP+PUqCerTqzuVz/O0O7hs45Rwv9qgjZG+z9bGQSR1TwQXdWQDcTd
ESvWeWndtjI6sOFIdl8K1G0FntbqrOYsaNj06sTZL3EuWh/xfm+uyl33ezf3CEJq0N32jL5u+hpg
UlT+O4gHzT94SjIBj+xqKTDSPMzeO0MUaFI7WW3zw8RP+9MXqoCSRGTfSlXZu/fOXaFKpMNXb6Z0
SfGgEVow/+lJE6DT6crkmZIuKlSGpDqsrW2Mb8mVs54bF3uy9h1kA54/yLAgsLD4IXmj/BO9uob0
/6k1xXEABFqua6tMaN7KZs/vc/bZfdqsbidGofuMxhDRdPM3MwU/EXo7SKqG+ME0jcmkBypFqP7y
5KDX0erxBQovSUxiuUzTTbvzW2xVaoYQxlSS/UKObDparZjeGN2QtXRHxxVtyzi5J3XLUEnilwWE
+w0t0yx9C/MJsoOQ9qPX0PsFbZykWhAJnigMi/IaPB7Bi+JVvEYGECshuxGUBcGpPwhVyYYhkH2j
vb7DEvyeW2icxX0J++kA2xCdv0OqHrbXi74u5o/d106Dq2jY68oMazebd42tLrmJEVHPABxPBz0o
9a+LwfdnLpsG8clF+1hjAoXkX8ih1W3E1OufYrHk9AZs0VcMQsfrDzo7hiXRsLid0+1PTfdM+Ph/
yznWHZw4rNX9CrV/slatAThnQng3j4qV+gbIFni+qfvzHXeav6tl+Becy66O5BANgLLgW25hoOQL
qA+OVJzEmE3Wk6MadJ836Csm1hfhuK7j80VwTCqPH6jTaEcmbfYBL95DjMaCM5RhkAfeLvyysqH9
Aw8y4/SEZ0qZi5dgnSapCvQ4+3Nsi0jr2/1ma71ed/BHpN4DkmCdhkve2E6xZYhvKwR32VlDr1uo
QYYv/XwZOL3YRdNRa8C9NyWQsSxTbGCVNl3L6Tm2PaPhMNN7AsZcWHVPrGtT47wpJCg47Pih7IqP
DO7oL/OljP0YBpR0SqCJnrcVoWexCTbiljmx68CVJlSDhq2esJH6+ZhGDT3oByyfR4rnzrcn9h7a
6vbQrvFtHmUH6sSSgsWtRabhY9X0YCZDKNmwAikmD/6x6Eju9zZKqTn39naBnNdfQLWTqMmnDXRq
63cb1vs+fUs5rz6aBECrVmp3N6HBxWtI4sIkeog7YIegj361PNywkPGJQIKKoHbWjGMgRZvavJHf
nxF0MGr6Y9lTCjsrdGGqcSlkRyCxXuUtf8E53Wbn3TaM68fKt3wvpqyAdA33qQuKEgMO31s9cTDR
Q3Cg9mR6fURj2TxO7XBQhw4UXz7U/MYP8z9HKxtj1tKJqMh/GD9ko4oagr1wDuf/4jM5qZtByb49
SOAibm0cueqAKEujAdtkniDxxQBjTVDuB0wAwO7yk/1JRBMeqpbRueeWfvYkgUpyr7xqmEj66FEH
7jPOglsmKdAyc0gkDqNRupf4vhptchH+DdxzlOPrhIk4nrAi6q7vwjiE/3ORxESfVIEPTN60XLp9
SHlB1MnvAgga1R7jmyI1FAnis3ffQeJDpShnhF5znWGJSXUCbmhs0atLQn1DLjR6xufigWDt3J7/
O17D2zbDZ3HbR3+7GD89YzGqu3sxR5/v3w7FkqaqtICPZaqscEQYDfLtnQSfirbJE0mmBGbYvNjs
0vMSO0Dv+O64ebjPE/K1ROYxinsU0cY83+HoJmAvUfxGhZMzKhhvV2pkJXpQ20HDX/yyCc7PEPKu
ZEDq7wABwZJ9VOP8xmOErtFNfpp+llC3J8Fruanq+o+MBL9gPUM7aDyjMLJVWQH3K2Kbas6ULFwD
df0R8iW2uxvqqWFVjIpz2rQ89ucyinl/eS5YOPt39vXa6s1Gq8GZwrEDkPgocq5YhjZZk0qhbxMu
iGsz7nUWXoZ7Gag9NuWOx5F0EFiIWcRaMQ/7ztSeun+yXWh/Mspd+ryn+cPTEAZu9yYHlfd8tq13
RGBSYR5PTHTxl/090sV8gM4aNpodo/0KwplbNlc4kbCG/NV531/gAqgw6R61QGgA7tsXiMvqXsPp
TVpwSECbV7UFdCyXy46/sXsCtzdeZF/ZFVIHAOlVbHuT/P2wUr+225uJwUcRVsSRzHzZTQzFR+qE
HiL/3lhEadiIIS2egaZJNFkQyWz/BPIUAWPLVenhlVmAB3czBItvtDfiaJCesZB8eAf/Zf8KhxZD
wq0jzqEVuNoivEIE1+o5MRY4c0/swWeNw++5MbS7y9hnEi3FHgWhHuIImuqFY51tT9D00Mw1WzL6
QQvMFmxCYx/RSGOtIckmQWVmMMh5QXnOOvwXgyr3G8RqeiH4AZHXU4jF2vT76qGsLLZI7buOllHJ
BUsxPPhxeFtfBJhuqEz4JIUzgtqwDBuvSQN1BSclpdgiKAH7hNYz1QD5WOWWbW4p3hegMTDweROB
LUpZ2wlKpY0BuMtV8FXXLYCl7NcmJ+a5zCftnxX0foaBNlJ76M3LNjg7oFQ+OSxyIJneppedcktY
AgfsAV8KNeN2NsgQm62h6TYoOMmeNBeaDr3T9QJZpEa00aaI2KslbunU1yMX6B9ovFPLxCnKhgQM
YV1DW+c7J1aLzGMO0iHOsIn895r//ApdWeHWuLGZ8Xws5NlluY/ZwAXSW+pxwdIf6MwVuPeGqD8A
TgJ8xLAxslTdCCjm+oHNpEeQ/X5+BAvG2RsAETcI23FX2bnvOlCQRf+DQaqdXBDtbsy1Ts2Lokf/
+2QVNivVDw42lpNh8GXA6/JXafpaITjfdzhqNxHcCIRffIhRglFq5jt5NlcIx9uuTnh67H0isDkZ
T1zUHinvnk/cs8rEyTgQz/ujWXcNVSL0vMRIOp+949WtxnIf907MUmd/URh7449zktMLIbmN8cQk
kTOYUOMkyqrVXkFFVGUI1Pq+1opqDOWgtPlybfTxrCJ5JctSi0L5TmSo7XkJig8PpWBgFSLmEYJe
zTf4AmI+C7vR11jjzcW5onx/SFFaRJ1edyYCOVOGSZGEC18nPy7Vnb/PGi5cFNEmYpxgnQ/TEPyb
BNVL1L1d7QcAunyaH0ZCARzdgLb9s1IhAQfyfIJpgbPklICv9MAGAFSXX9c+0maOESGkL1eXhKdq
tQQ642h6DSnA9eNfKUsA/tB4Qt1QjVALlaiJR+6hvh5btHgh2qGk9kj4WZlT9LbicAA4+3YdcT7q
HztakSrVvzdu4mbMc3QcdwgifM2C+OGe9CBWb+oNnaq2faz46HzK4AHlGWCfdg3jgWrocOG1yn1M
nsxWul1kaoDsBe/ZsgKVe4HTBro5IGDO1L9cwdKeTvdJVsnDPc+j4I9WSJRvixZuX5O5IMylw2QI
OFBdZczexPBsOM+ECrMiapxGtFCPetIc2vo4OE8Tcg5vom/ylDLidhXqsFa+yaXUJJZO8fLJd3UD
XosPn4wxbSrsWhnVLccQ9VrK7R6UuveEfVeeTAWWzOcTnIeHjMfiX7Rxfzf6nxKlt3zu/XeKxLmm
i5QOZulcrkOCbSl/cxxUUw/ywztSGmI8jB3gj0rQY0HIR5uMfvgyDY/7XPCT8tjNBpOv+5zI4+OQ
rjWNVjMFwSt/XSh4TjtonxJsGtWNxRnavmQ9lzTB6vTjneiLhxz943yN/8aIK7boR4dzR7AM1iho
/E52ZPrdHsoE9gXRZR3hLhSxyyhNePRqNM12sAWta+cP1V5b5ZDv8eF3zthNT6r0NxB6T66Ob1Us
N5x0RwQrp1gNJJlC0Uy1ZyVpuf0ryXy3lyH01icGjAZ3Px3SWfjBKBoMZdm5Ge+8IJJOkf81zmzZ
tJ1c0xhr7QVVoKawsn6GJSc0kPlN2QYX0PU66I9QhAxvyWkp4mW7z0OsbfK/qIr0AOkgScW66v40
NYg/aTbxMQQzBtkBp5PUIZEVhgIAkL53O71qMaTvKqSIn8K0ZbGZYTWJlH91kQksruaNLCqo6Kng
lPGM3ayLhuFKQDqMbD2nmK0hpQu81O/p/aZasN5gJt3maz9Sb2cczXVKL+oTCWaJd7KbnensWZL4
rM07ohn6hej0RwybwEA7Y9aC368YP3VtnqSYFpJFkUaz3J1mLvS7/7GmiD3yzwIwm0j3uNZoihH+
qe78/9T1tvbiGHckeHuYNq1qYh/D2KH3Vh8zCayo9LkYKm871pGKITzzZ0vRmwb3QuWEwIlkqF2c
MsehM+DCvmnR066JjTUiZ/Ht2bnXtzquXv9UO9r55xfnZhMiGA0Xe4Ti8lahdiHZ7wb878l0ie2k
5gHIuroMVbYaTT/0/bvZ1Tvm46DXUjP/faoFcOJczvNvdhzx+Zmh73VZa7HvY/fwBXGgQP9N9n/9
D4ONGnCjeEsjEPttBVrmGzhB7btc9D6LL8Er26tUu+eCcs7ymkRvRmv7tCm3iBPOfYWHANYWIt+f
ANXbf2Jjd6U8yQkwHypzoPdJxIf0dizfYdEDRjhd43Evb6uB8BZR8PlqCyA3QxmnQDawwZBnGy1P
cx9bivsrl/stealCCOpZF8CzdbnotFnTvyPdbNq1mRgwY2JMUdWM4nedPdsuM9sAOzWw8wrbQC/z
ClCGIs8I/suBc3dLzpNDO2mu/4wKdw/nJtHoftEphgjGMrePIoFgvEwxfWm8yQQqeQM+sTNrb5FJ
vRWtItrWMG5gsBl+Dw3k69dr7Q/tkvZOz2lpIVnVfuIkB0yJvJBAVuGe98b/UC9WCovZH97MBk7B
IKAd/Fg622Xjk8RBXk+Tj8mw1vZcvI6DwpR5vPWAvWzf+0lI8UFmHLHJSqEBLFfaEeVyUUcdErIn
5XB//vXmjjf4tbRmMFsRhVv9/6z5lUkYV7pAvmtGLvsEuUlZYjaZnptnPYzQV/OyO1HMhjJwA3Yb
owWUJyRd6BTgS9Klkid7dL87ZgcD/wyZPwlRP1MkJ8PMrM29hRnhHWBRCZK/j9/bYyg68baRFcPC
lZ4qkJNkz+PUC9BhKoAfcQ3baYtrxS+MWAjhoobHHbDY3VQcMKr+2U5CL1GMBHkcPkmyFzlz6dhQ
xcqesLfYfWjvuQ2ES4RAGNLwPMcFzknbHB1FfSj3Nk0ce8ImDoEG1QZ7D+CNHydv1pXCxLmz88Y3
x0ljv/1+JHK9T932Xzmd1YFWTHl86tM259T51WTTy6pDQMqfj59XMkA3Ah+M7HNyJiT6Fmhxk/gi
7z0M7yGA4dOiQ81HzJNn4gg+zGrWXCSQg85Xg3YeQnLQ4RUKDf63abPolnrbfVLS6+SXdbbWAli6
06ANjwa7f9bAfFD5NijUkm4z5xrgQCf1QczRx0z4KaulmK29wpuaHLHaWSTpM9+byI3s0u/+VWum
igeKe8+dcOH+LfIPGIJirOQS9zzTG1nkMFBU1Vd1rQPK48FH0pBwbjGvbJoQjQTw5iifm70yw1MB
qcQoSqm7ERMW08VY2bvRHvvtw3WmkE6p/h4bBFsiEkrGxmAnlEfvhsYRfREFX33ncZaP8j7Dj8Ks
6izrUYxgK1tZuoFhxjv666g4+YlIlTAdWwi9tmvniR7KR8rS/kMpm7ScNPO2Q3CH2MPFXInHo7T1
SdLBqEcn3zFsuL68KNEHZKuqQZ/PYWi+283mYr/6agIqs+inJaxacvPpSKmA9Gr5mw/tRkW5Ed4v
NFCSmcCjraktB/AyeOEFNVWeGGREW0Ykgc3HJfIvwr/7i21PZ/UKtNafJohVxjO7o4rqB/qc94o9
068Pf7Mjlpk5DeGD4R7eGigXBy6z08jtK0xcDI/ovbTc2EF6ldDlUptSgeo3VK15nys53CUHGdtz
tnTRRhEqSx/EliKJhlnWHVG50eAyJLUuLdm1P06QzN09n2xE8ra/Kp8CaNEc3efvuHDNs0gOqkZd
9H6iRiuU3Ly8QTbehEkPucnZwOSlrfLyYoWCksbHP0f6j9dCO1I6NjcyPPfgyJklttKNB4DeQx8g
PMINBsAneX//qlCfPJ5xTYLg21RB5TtFus4vy1H55+Uzyp/67MRd7ZYSvj49B+tYQXTrCrIsb86a
Ghi0C/rjlrjZyB5T7cKkIwnL/sHIowNmiaULPTWJdJnl/exhfz3a3SoTO5cCwon4variGjbIa9nD
7YKpD+Pq/LO/3N6qe2nct/ALAxw62ZJvNu1dkpBLyRNsMB8NND7LjtRSj9OLZ0x48HsF6vXmBr+J
fsu3RVc5CZDTOtEKfYSjuvORHzPF6chuTqAB9WjHOoB1vx6hazl61l/lmvcOqS6n68PBJgvhsyhR
5aFkiYiddRhDFVPi3FBLyw8q08rBrjIp7QOS7QsjanqlqRo+8AfFrNoyuTKwr2eA5s2hrfKjpv0G
H/rK1yHOMKzqFqz94Jol6ceOGbat91/thm7GwP2U5FJkUeHLZO0v+Y+PDfTk/V+C19r1kq5NMcwr
TQol+zwLLV2ZNFrckmta+J125z4z/K6uwn5zDC9eG2t3Zm57YOxuCBIHeRGzheY9jE1yMFxEqHIs
59/ubvZLtR1W5j4RgAU397xST+ZdsIvC9Ib27n/FDjOuUYqIRYdnQbLnaVAODtxr32AoVOT49gGb
vx3bzPchRFH92ijCWvopzOpj7aCUmhFqEU5JSJ2cJRC1woLNOl/DmmR/bjDAsKMiXyFrhlnY7jiF
8ZThG2iupe+gRNy3b2VGCfyPYHZwnP2SxDiG3IVPuHpDGqJ2KCW3zTIxwaNahVgrN43TLqDPTaOn
kusvANJ4LFqvX/RgCGEWHU49AhT10teMhaY89v81hQvU+zVlnK/Qg2JwJQo1jPtQ4cg4V34FDSPw
/HMtvyMEJR3RWp0TFGD82vvuENg87KcaoCMYU8BPk+0VGlt3n99Rh/NSp0UhZgtbafSF33rjdmF1
KMvw2GLEIi7BqTDwZOORK+3EQJIfHwl/aYEL+SROpplTkLzdr5Mag6SK8Q+bg9mXL6akOpf6nnNI
K8Nve5lNy5v+9qDz55ex/QW5fad+GV+V3iPiNihVqV+//IHEegZM3WzK/mCBEXFQz2XkTDUKV8gB
XEIGZ1LxFNxftwZtrVyf8DQLT20b++6wEW+rU2V0kqvJeqwdYFwdqtB/gVyhyEqW2m2Jvsq25m5R
bBBzVbjlM6U+gOx4Dd8gOVtcPOZJAjuN82uevw2a9TnS7wD+dnO9exdrRD8k/0Qpk7AR0E/khZaa
lkZsECAORNLwHulmROMQArBWiX6HDycq1l8mPGT08vpo6Udaw9qYXmNHYa7Wpf45ioD22+INp1Ux
OWsBgG6zME++triQ753VuC3olXlJvbWXcuK0q2EU/PELTPuutfG7ghYJzwa5x47KLSfJL+Zzfgxe
CJcSWiS7/dHWR0HmnqSepu+iDXIT8M1x4vOUyE4PSOEZ7wxnr0zksfmLbFkROexW7wRXOQFg37cp
4GpKN0b0YC4OIZTNKsKwLIVlGve7wqrh0V5M/O5Hkx0CstDG3w59I6dPUoarUjMDVjLSXbaAadla
4pQa1FlTaoetWGvX4exTFRxMog7k0Mt6j2X5ryZ1Xh9Nqcadt77PD4zfHNJfejPtM8ofd8BgU9so
H6MBrVPnIwt2bU5M46qOS9fNd80oP6JlonZAMtUdv0IAX5DTqHFJI8YGbFy2xi7WWFdhF0c5y4dM
qnrVvVdKeDjHA0m5h46vxRUG3bKFItZZtyI9Gja94P3TeG+V5tXj0YoN2lZeZU6ca9x2TC0zfh+6
6tOAW3TEzozSq/NrnYsZQE5wwTPcwRcSZr0iv+0QGvB6ovrBN6a3y+tY4W5yuNGLYOaalmc6crOH
8N4UCO3PHd1k9hzcLRoxj+rqFvy47xwQSnOQU7eJD6c0F2bvO3bOOM4xp2wXJpQNA0Ey6VCbTdfj
x0B8pi4Fb0cjkRNJsv70WhKnyqHZKmFcB3JRtk6hHDVhKVncNlXvThdJg02iHhJcjhfjpCQkSNPm
y5Ac650TZJHHsgkS6NutnNK5zykZpFoFu4NLSfmgxzjKrqiAGfNodW+J/LyWZesZW6k6ma/7f1wn
SMadHHN5+QnZfD0LFBRsY7q/0FY0Qg0Hjdiau46+qUo+PPT3SOKabJpbKcFL/AuAsYAlfITszdaY
sPSCOUGx0It9TQfzc4elpP15M8nGkypHI2NeWK4h24YnJDs3tKzC3U23pa+z4X0d1f9zk9CBxBZo
HDQW4LcNr4LpqGYFmfYc+/pCmYMGQuK/10P4qRo91yDN46qQA+dBskmwy7x6/WX84wYpkTwMv5hD
NSR6eWg+8dT7ZJyBIeB1xQaQEItp2O2XAF/FoeEE3l5cpHHiDUav47ARBlYAFCc9Zlfysrbl/dS+
1GH2+7+H8+m0NsbVsICdh6S6uJHYmZdNJu/I5eeQSpjkknav2w+ikIJSJTHl6C1FcIGUeb61ADPO
VXC0h60d38Sa5qKT3BL4zkXENqJGxU3f/OoMLSk9r3JBmtt+icSWo64o0xnlGTe2+suXiNA24Igk
v8rjduHqDoreOslcMyYqjQEei/8jLGT6Jr6ct/dmbUkng2lO7brZvn2A9qr9DcVNiVI43WA6U0t9
S1BNQuMsDwKqChVuFmO8dd0B/XRIXU5aQWVRRtARo8AiOavPU/xOH2NxGM/RUNraJ2HgGt0xIiaH
vCOOo0kfLkYZrejpt+wow2GJ3bLjCxlO/eCePMRDARWJjJibywiZWH2CZ5pGgv0s9nx6EdvsNhaX
NzfGLM3S8CdEu/6J6oSU4JCLZvZ/2Z+YgrZFfRDGAknLWM5tKjWavO2K/njjUwe8R1NJRfX+6Mn4
aNsmRRULz1mMRmWDcpkyHTQoMALhY57yOpmliisk9MQSsmo8nvXay+3aPz4qxgfEC5R9Z862jcvO
UiQHwFa/5JmLGvy/+0EY5djsjB9dVFf29A4BJYnFyFYr8U0AkGLzZWQi0a2efsaipcXOltJn52VM
eKQo9GmD2Y9rHbXDre0pbY6UXH1hikeEBJ9l2866WRuvAs9lgSjd8/zhETrNY1xKFMBLRr7lYb5b
C3wQcWgSvDgqdrx2Dj8SWm2FwkZgcY/Z4XJc60Pg8GOZTP3+yFHVuBg1E5D4agGMeRjBwp9rdoXf
tdOjvYTaEn+xM6q+hXjiT1jMGq1m6eRhdlk/+HjTXc6847a87SpDRFVP7+OjQosUkvSgRXJmX+39
kBrmdIUsGDZgHCe/OKsVamHMUKAHs0jhcs9b55ANqL6iRNDVPbc1fzJWG46mDtR4YFqIW1YCw+qV
TQH+NHhruxc2nnuFyDx/IomFqtqj9C1bZt74seKbwYPR+0cWysnbAntKU2L6xgcwuWbQq4o19FnD
W92oOmtnZFgpgrKvpHsCkeH0UO7oyzw88Gpfg7Ul1P8cIi1paZ+YpVuoZBKIJ548p+Hos7ApEevj
XWMBo+fdDrc6ONyoi64lYYJ9yIa2DCUT5LXBlVwSgl/JD7CPQL3vgMm0rhKyM2ApezKeDYYbQ+cP
faRaYnpKxoGpVIUB1qXUtMbaxgWF2FYMdbdFH2BOKLrpOTlBpIQsKipG8uycn3dWki5sZzcTYGmh
x37aNd+nr4EwgN8A1i/qsy3zdNzL00bbMYPsDXOh4FBcvzOeB3j7L+L39aNxIp092ESQLRzh2frE
klIyDiXpZ+57JDGBPseGTGcB+fCmGdYVlgGtRSlebl+cTzwZlhjjJwx59Q2LSF+Ewt7PlvP5TYJv
AAAiR6poHS6utLoWZlnvmDpbFVLxmuER0AXbdWrY0OLDk4v7A7x5inGn9PUf28gymM/fG1/BciQy
GKmlPjoRi3sT0eWWRZrXU1uW++ORtFDGeEQVm38BmU2IGvXjPMACjfB9WD32BCxv/6FdvCaPMB7l
q0vF1XOZPFwBFGUOG1U+gKmseVhlaYkr9yQeYCE1+IFs1+s8u7CSNSov8PMHp8P7hzusyq3raTMQ
9VUxN3cVNhN+8/Zm7Ng8mfwO1xmvIjCQqTOsDwwMGXVBk/Coe4c6Gebz7rIzVqTzBaZiu5BV2YwC
qJc2PLY1m3vPdLmx67tE8x0+E9y3lYPF0VmU3cigrtb8/dZ3zucefbPgDsyslhYO1Rwr5+x5pMKy
4TM0pmMt6Utq2xR9BZ8aqTXl9GFVhKkxlLKwKPhPke71MDCUr771TNuNU2bvGEaPjCcz1MF4anvu
z/AJwgIP9Cq3ghnfdnUwN+a9poG1RZV5xzIqw32tHSuLhkLmc5E+I/xnTRbd9h+mMP/OPDNHNXI8
cX1GMIDf1RxgN6f5AA8NZcdZ+88rYtmm6PskNn2HS8ts+5T3IiKCszqTETKgJQG5Ju/KarVDBLS/
3PyRrpkLYx2SMuPOjflMZ/jENNOJKTpe8w3k3vdQQpHV3HRAYZ9qL49jXKzrMNsV/h+0l2ilsHBn
UuxCOhGp1Us0TIT+W1r72sB9HxSOo0/T80hGN7578fEVIHCJ043SMDYe03nespc/1vuAiVqMiKot
VflvixjieMtgfFBXz/6uHH0nKW8Hx42yJKUBft/ksrlbB5JfS8ZtF1D/gAz6VpWk/su3JPalthsc
xk+mjytSU5yUJbn1XCB+yqVCPXdZJaQ/sW8iAZ66wC3x9eohBBSoH4XvIOmnIM3SL55Vy/ijaW+G
rYqHLt5iWI9QN2e7RGJVKWNh/G8TwCwux7n8ff+q6NIbfypuTKyThLH3Fd5zoizagKlCeW2nZGNM
CAnaZiTyrajy2JnPYbGY5hoSO4HYVWnTZgIbBhfz4q/Fkn6zDB7fMsI517PRUPnqFq5aJcU7BunC
TBnR7Bd7x2Dyoeu1wNj5I6UDuIO1jmlQcKzRT8M/ghB5/hwJb4zRGQQoWjnV4scDHGz8OaActaXy
g4gnht6iVVUsVQidgYHc1lJtaLnvL/ilPXp44bi3vBEp5a+w/HKntXqzmYCPoJIltZxrQ5q3aq++
fhidtF9jnXOZ9YH2TTltrynAVBAH7/Eh7r670D3kselv1SbcNMXxV4bM+0W0jOJkZzYf+eWhcRJg
YK/sqZ/ts9x4ZOxzGIt/kg92pihfgeBLVxDYOn2lxZZfny8/ZW+X+XKKhaqvlVQ0xAi7J5Zawzai
19nBcofFiMNKTZtBWvozDG06v05GNHKjq8r/wu+mVWJMgiAKQO/y79OV2GirTWRD62CLCWdx4XW8
Yw4xqetPiApSQ3kVpN5UQczkE/8fU/FFFZbG93zNkZxNWp2GG2P9LsJQmMLbzTb79vyB4ztXuMyS
F2t1fi8396kxDL2eeAmuwud+kadw6KR/cpK3kUVVDbDlZhuPRi4f8sL2rASkv9Cw3o7jKn+5GYMU
3umJsH4GnFWisBePsHwxrKlhrOZ1A/on+HFYe4WqPvC8KeIbf/+Kg8bJbrZ03zl+Kd1JNiD+3C9A
3/EB41/AZxkFPndNsjyFLJWY6deVwyEK+ukYNJKreYmg+bo4Nx8GwdRudX14fvWGv3TuxcPAS8NU
hxWlmXCiTjVcj8mrJrlI5ygwJuSzk6oJ+T7x+0gmriWy6jsX1+1oj2J3JO38MbPIruNjuHCl3eSZ
axZAcZcQSSvP+1qdoxdE7c9MrE5ndnivKTytXxIHiQ//jyaeHx1mvGimmOnIFOTZCjim/nV6nEQp
iegbcEcUDTfYjM3x8kOWAEmVLvdljDjQq1Bm5dhIGRLd1ANOuEypfQyLyd144awxlSoxjlZHfXC4
mzPVsIKZLwqKkWBH3hE+En0Bwi3v8u+K+VWsNK6FW/tBm1q6xNh5CImBmXAW4FQ2J/kH07nAU2KY
PH2+Tx0lA8Zv+LnAarK5CKRDVOkI00d6pGpycCv67obarB9nkkSv4ProHhhi4zLOxp+coLlXvnWh
wOaux1VHGI4qEv4ux8O9OpYU52jSGatPnl3BSSVT/KBtDCrtqhQgpReGRBs1l/51nG71n5WpfRYA
084i+QqjUwk2xTxHfZIc4BLkxO8MkSDQenrm4/duyyFnIedt13bHURcQE2tvmsHSw5/kgNAw/0+Q
E2iUpS60QL1lUS025dr2BJYdre3/XB6QibxtSnnjovdEbHfzFmQP1aw7G/6No3Yhb6M35zfVazsL
SKgiDSLzOxrBsp/jSV5lQyFnLyGsLu/8zU8I4IwHfsPEQW4X5hYM7Xmi3EloDNp9XBBhpOOdtqyF
xi7KC46dqeHW14u5+GEJyXJWEe3ErXC+YMX5HsYOLJhdAmAw7BR9b5iiv8Zj0N9e/F5VXO4q4LBQ
CeM0b1QFXpjT/PQeKNIIaeNwcZ8A1NVJPV8Ps0kBh7qgzCTq0oXy+Ad5C7E3LKPBuziBmTTvo/C6
sxUxZGYI9r5q4+sbiKZd7kQbKhd1Yed2JRUe241nMO+/p9MEeg1nYFbRZ17cxZD0+yxrW3MKXU6R
aa2H5Dt9cVi2TtAgzKoYXkt1EpqNAvVmGBIBZCf3EQJ2r1xkfoJVDpBRrCqef3QLSuLIDZm6DIYf
KiNj03AJpICg6WFIxlc4hrivTt9X2a3c1ZliJ2gT1AzvNI3YVVYBDw5uGhn0abC6JNIKb2T6LQ4D
0KAsqX9E4G1ufjKjSPbneC0nrSXSKjU+pNovpg6JnGBF/Zv40dFMBpf7n3m9HwvDanDFjnqrTSGQ
QLTtDgrSYOKsunh2/udP/f+5xbv0E1iUeopVwzduSJ0Td4MrUboxFTyD+3GxnIGO+VbkL9HW8M5R
BoMxC2vJdcU0jU5d7BKo4sKpPXCmFvHagvNvAA5VclOf8Y737zTWaYn975dAxWHVVgrJcnXLWdNy
nvRGeQG3FKquwEWHhWLH7LouLiBvkwfcxx8sa+uFwEc7oiYujDiyQ8iUOPjFinaxMGRP5vUZKNJx
Vh49qtC+RPRU2Rp3spRqRDoYF+NTvw/bKOVsW9ji6Yyjaw0Hb33FzsDaAct4y0cb5NJQUxJIHaRF
peuylvvjOkwltVFKQU1oOnyYB5W1YcBEO72slSOUtIQRhK7DpqhtJVcNKAsTJxBWD4S4ba9OwTDd
70QywRXCkTrukp8yI1s7FSIAw6O9E8kxTpvZqtEwo64MYU49YjB8cbRLGqwiwPZaTQcK+gQCMJtN
MKTR5F9w4aM6fR5RtNX/qDWg7mgtApw+kP7CP3VsVO1DZb+ETKu2vJ1m1WGF8ymzrMZosc2ymSB7
SbTnYXa443zjx4asw+Jd/cLKcPgDkZoRnmVTzqWZ2uaamjNNZ/1pti81DrnZ/ciQGvMHSngox5Bm
/Cfrdr394vEyv7Tq6rfO34XgRQjQG5HSnV3HUCpm09fQEUGQ052dACyPGnA+DDD/aU39O7F3o2tH
8qV2L4nuaqjuyA4kB381mpHqZ3lMeZUx4pbOX6PowQTgfBeHZx5T1EdyIhhKyniqP4K3y/9fNaFo
hkyrzKyCPLs2xp6waHzlWdoiN9j2McFnSEkO/dRmHcc0yO2sdHRp545LfOXmDOvD//fx3/Xi1wOn
gMslexsJDdxSgOWBUZPzxdWtWhi5cGnw8m1361MWbEBJTqRS1X07P1mi3eGIHqPnXQE80q/WQMc2
WEKqoD4DS1BT68thd0oAYasjIE1auSXuRBd/+ZNQUfANLfmF6fGYABw8mKjPtN6emWvTOG5nYhD+
+9AHxfdpywKtcvG8zCIz05l/06eZLJsh0jmYXFUsGfjfJIdubgHbHirMRdICmmGQFFyoQq7J/fhN
eXZ7U3F/oJ3H9yX2kQghvn99C4AKLa9T3qGvGMdyvtWUKmBpuqNOsgzpO7Wqea5pBHRTB0JEox8+
9qqlg1U7pCbIwui55JSmBWD4GZqJqUS1XesHyoWRfnzhiP6aLXk+tMzRT9YbTLG8v/OkgGFUn+n1
RmI5OABpFL4YFHQ3ESxYZFHVnUDmbTG/RdHNgjD85P7sSLnnqZICyd2FlbmwYwM6Q1+8k5pV+JYS
pg5G54JI9QIRPTJSiLJpwq/achReF9jaC6ZRvjcxUoyLAMVdKMEBHG/FvZWsEPHR5V8QPFdIzPwS
4jIj8s15HgBUWg8XEFtYKzptE5OO2kPXiI0qUvfQ3X8GHCTG71T0sVt/hBIoWlnFTHxRSP7dxdr3
7rlUeEVYJXO6W7aobw7emwDScTiQ1QkCG+Z70uYaR1YXnv8n/MRjW6DZFPyl8ZAT7zhQoh2jNhcw
iGiX7cu3EGnegdOdQUxRCjUkFqA1qbLqmW1BDm4qnY8XJOysSNurDqUAHUZ5+9nxy9Le0+8aREVS
cWkfGin1a87A64XOV/iGafugo42vhn7OwngEGbAA8BTYgc+n4m7Ol7vdZFtR7F7zDUVApF7xvZZ3
e4TB3Z9cy5P45k2nKr7kLCUtlxdtAaKeglfxGRpGr8YKFiRBuItZTJTSPtpGvmucSkbwnecb3PsP
0k+hTh6Yiq2JntPiZGw4vSo0iU0pteAA30hgfwqPVPipXBYHfk7XwsND3v2l9ZYsdG/18f0fyoP9
7PmBRjL3qsELTVIA9x4LggxoltXo/kvgp5nJdjg49h59KAmNspFuS++CGZgmTbsO3yvGkmYRZvod
AKc4Y6SbWg5N4pSt9WkgdAmMZHh/UyLRK37RNqBc8W7/DrAJ4T6tlqVUPZNxUYcCh6K46GobUisI
Eqq/nn9SfQmBAmzPjEmuSDX8PAVW6Zm6MH02/SStjwT1gSYn/KLKJ12ff2H7wUKUkhI+rg7f4YoK
InvBOSTz8Qdyuz6a03ZdYBY9hlg3yM72i5pP5R9eJIvAed9Tn9W5buAVMCaKzpBUv3Nn5PoLfzfK
21AA9i3YlaPNSu0sVQFOj/xDRVCST/z4ikOWh79cb6l3yr06eNrIwlwlmDZCDPyX7+43Y4vOp7/z
kAir7KAnUgIyhYdqX/Npd1GakcKJVU3+FQnQhnd4Kv+E2N9DZu8+/KpZ7JG5Jao9x5FTknyS5zNQ
H6a6GGznEzIXc6c3yZ422GabABf8taclCgkB3lvSoEEI1SuTr9LEl7KTQCbEi2T+0NpbZWTkPEmX
8Bqp0tZe/e4YOMmm8NBOyABxXDLRNvY2wBJ5VHgFYijuTIZ6I/bb1f8mAOJVwpXQ//oBhrOv0ODi
PvEJRV5nCWy2fSvhTADFS3UeePMIlPnnGR9KcLnTddV0vtKJMIutYuo/5AQLsda28N9UDBSOJ/L6
Z31NQwOJrzY2mGAnfqkHB6MaVOOaJuvgXnqgGmo9C+HIkCdStikwVMkKa2P5dZReWnVWL9EMOE/q
2lF9ghm0+pS0n9ovz3aIp/GPCECTRxUggLiA3+/W5aetmYBi3ADB/jMUfHwPFgtVH0o6No9OqwRM
1RArI2FrQWTWPACqzkU2xnUXk7++sFjQB1cvurn5xG7ML/25heJ50rHcEo+JiUVNEseDaHGqjF4K
5LkICnH7xBcmKdnERmOZf9aYimbr4y2Ee0O1UjFQcrzE70W86h/xpq35iJCHPi0Tr4ZW649dcaOF
a+6v6AOfB/V5jEiloy5GCLblWWcnbaz0t3YQ0j44uxkqV7iSVeRwAXxdP6dltCf9V4cp9gzKRxq1
H8caSUpanpIffG2iOl5kmaJZFb30zDp0q86hFx/U4kTIdqoKB9I+vUDCL+RHJRDFG0m/RqH5SgxT
LqevhzTr+YdyoYX9+A/pWBldaDdbQYRouGADf6FCvCjo1+HARPmg5YJyl0hNd0S0fxH++RMb4wA0
LYyOkC2iojuOxasUxnt3VXApujrdXbATgem96w3RfBGDEs686OqLcLuLdr6DPeUdvcZP3HMCWB5h
sJk9iTiRgNXU3NkGYFzMgy8AHArqXFmTbzO3F1rSUNqtYhc4bpVWXxwb9oNtRclwXs702Ab36cWl
WdIKRFyOJQN/jdX4CTWy+HU2OCaeCwuNdP9gdSYqIIvMuT7v9gOewlPfcwoq2V47HdJ9vnr9Tr+u
XgbkOhWvn4lm8u/m4fNyU+np6i9Kg+/s6rexEqf2Y29k373Jlcq4W8+Te6ksKksiCW0HtCqbhqTd
pd1vRJiwd6sMaLAJfsQ17hM6jrPw2bIaYKLM6/hKIvumnlpnfkzVAJU9SGaO9WbRPUZjORMGJNuC
7K2KJPZGtBD3Sco5y7ZILkub8BzStLfbJyC6e4inTUeCXiP4HRhBMt1eSkSQ7mZD0M97WGYXF6pW
5tvKyVyi3S6AJUXOzwNK7Ds2SihLOI8sl00yUAKCxBlduF5fsHXhzYaTGOnNZLie04AVOjXWTanY
4VsSVbF+fdacTKq7rwcatAdvLnS4AcC3gpW1xNZrvX3abL1+X6H/zAQe4GkqS3pD8qunC8wR+V7s
xrApGp8ToJOfcSIquc+0/ea2mkqs1E5Xf9r6u/+DkCyfOLudUm7siZfOrwqq92hcHTz681x13duW
qyiQ1xZHrC8DDVu1Ky5ayq6JcaHBJNVmMeKNhbQDtqgmjkRStCwDnRvLW0Di4HqAGfJiDnS42xQQ
p/EipG2w05Y5eNL/EQfPOs2rCtrB45cQni90GyTNTjp60QbC7wmbYxU47dK+orlP6MhZI12r/jm/
w3WznXyI14e48FtMZeO+LNl9po2RN3H63AlFOxpDKfA1a5Cko0h/HTjEAACV9sMvoSB0oAnGEpd7
SiYl33Nh9A5xgl/Jwd1Hn/i/ovM/28Lh0i9E7oh+iXVMkytFNBIGduxPW8i8G2as4tzdrM9WSPlT
wNRUZFURfn9g+ZcoRl09X9AVtGmtCFqh2WZcfanJOVQxkOwjAfiTWrEMaFKGRlTc8ThtSQraEhRM
+bO/kDYoJivSJ3vC+vk25a4MsAIde6w7HK+cXVrUh/B+h5mf8u34O5AJ03yCsuP9yuzdR/6cN72k
9L0fB73tc6OUmtkKol8i7VFKVI7WmUKXbMkccbRxtgBUPhVH3g+qKNcPhuzfkdJ0QvvQ7AHkxQyK
+nupZl9uD1cwf6qr+WBYAF/eo1deT+KaITW1268Dr3v6FHV0+j0iVBEq1KPgdSsu3jYYHdvoYFNS
arrA3K+T4lR2+znINeS7j9CN7kqknotQTJcuBYTKgDb5ghh2BpBFpcDAb5NB8S+pBFuBn6s3KVjo
1IEEdKsAkP6DycANz558fhbAM57Pt87h5y9wpx9PAxjfGUq+KLdwPxPuSmZ+5VRHVkt13urNlT6P
oEWifkdiQAp50nCo1MOluazz3oCVLpXJPDxMm4JhTDGJdK+Fp5HLsoVY3NfF1Cwro8QQa4BEgMHR
O8JEiG92cZiAxkpQHHhZ7NkTWEZdkdDxANUwPqGhR8SrC93bfIbXT+UDNgetwJOGqnK/l6c7Nsei
uVqiJTvCM2HivfwuPYZzhBjelXzNlCVOpo6owBvCYHf67f3e4Z1y+MdyGr7do4VdEBmfMWLyBxXz
zHl8EMOVPal3PBArWpxOTiClcL0CPHQhKNQZjn+JebKSXr4JzcUyPg9z93sKjQBu0KgztN/YhNWQ
U0tZB3pP65yTBszsaFSjy5UevjUvGqD3Fz1jdvf/CUG9+dJvxNiCod5MG1860HkNIU6M1gEYbdmC
1K1FCRzS4xIA4AT7CokokqCc6N5f4HSaDgs17CirypEBJJnEejLgOvkroffoGzBiMvBH12ULeRYu
0GM1cIv6KUDlS7+EuMDL/1MonmLcpWj+txJaWtjbdW0FrXJy6UEIcir3I/uvR9t4+VqNcpyAbIBL
DmOe1cs1zJbaP47QOzWd01+fQ2p+xXFaK9plnOZtn1s7olTZTLYlc5TEDNYy8RPHeBnoGvhqHcav
cC0RAmcrWmkm0UspG4aI+ZwJiwSep6BTLhwARc4NiaKRm8r+CngG+BR9XY5YLbYTrs2/crbxN/sl
G28uu8euBWzGdkPsCUiYVD2Q6MusXu1lLTqsXLtVEDZ34nxGEvyoFL7tjeVQH8HwtXLvRliHRIoT
i6cLv29r+gmtlWGfzvCNa2fMvBvAew57e1Yj5n6xx4jfoNqdidXVbjdld4wXoZS0vycLne02cdXF
NhiRRF3vOlJYl47z1oFqaSs0InmM8SlQ251EbEzEqAsi6e/t3Nn9gL0Y/FkwcpHu+ZAE4gwyBml/
8i8tRcU6iXmqQIfubABmC+WKrndmSuPqiZ5uWOR/0ACFN2Xmc1/CGBdHvdH16tJRubS8+8vpfTyQ
yHkTIU0vy0YrC0XJAD8Hfa5B42x0+0XCmGPUfqGpcN1KIMGMRjKZyTf/mar8DngYj1iEDKFqrEOX
R9ycdWrZ8RAOMSGXolIoA8X0bHc9ENGQSTLKuJcHnzc50nEBAMHAgBBec/dOXR9Xro6pYCzUorlX
URHHfXYqVq0sHSNx/j4vLPYauJuk0BL8ZGYarEsfVCAQjXpYAvg9/20DphM2Uh3y9aRa5lh+22MM
KQcPPx2lmC9PNg+G7kQJF1ocmzIrR8IP6pn99v8Me3Z/DuUyN1Nsj/pDKp4vcOl/RVB0l98l+YGW
HDmcPOEnLLZBK49vw6K52OTKXMWHVG6RNtGF37qxP1BLJQthrkcTh6872Os2HeY51dIN34ePn06B
drGc0mOiIStKgzy/tRL5gvTW5r1CjNXZszGLcEtW/yYWDTvwE4urjTLnwUxNKhOYV7TOOeu62wNt
79PCl22LHkkiwIoRUG3l7uV2++YADhveTFt4Ift5CONlkTUp0c0Nu+ddX1UpiYwsZ4jfrpCrD5bm
jn9o0LtuFQIb8afpv8W9BXBpJsHSWJYxVgJZHaGZRFkSpulFApRcm0Xu0BnBtrS/0uI45MddsqRp
5snu1X7VWyX6log3ZfVxbYo3Hdt4v7VGspDzl3qf60hP+7GIRHb5FxT37FTOE/DZSE18EL4RRdx7
4xYwDLiKz+1fVt6PrmOsFjOPzXPn1KLsp3iebixQBJoV9vElOeTmqztriWxnr2uRNnv0FEwc+K+0
KQo4c+ZSkweHj+xWLT5t2UCfkcPlDjspRCsC4rBUxrW6ecwl1sQyAZUmbQGEPtKmPfyA4tKtwAlu
ygvrvYmyzRNrrgM8PyH9urXgdg87BMR+BiuEjeJojg9GZWMECxdtk2BnDh8h6b5JyMFwWPylC5vt
Qn2lNrb49wOJJMjODqeLV5vAROV2Pe8T4EfX0U2U0nSZOIu5iqBn4ALGeT3gjH7C+wmh0LyLFT+6
nzMVKJmiuuKrB5zWlWFq3/JNzroa8M+kTOq8wen1zARizhow0CgxG4j0Qkt+fbD+x31lkWkRo6MS
38lrUQhGrlbMT5v4XH4ORT44oZMC3+1KBdKAlYEpAyKl3QICn2adAYpv5uatmq2bXwGEa2hgRk1v
le+2gKOZMsI4gibuBCQ7waQQFc4+fgqQrTB90CvtlisPoxDLapItweNmAedVlFkOkyRwAJml42/e
dAVRV/z5oBQusA1sktDNHyXFGUU4wTft/U8+C6+JF/8usWi1SfqDIG9A3ywwzsth5d2K8PY2S5pe
7GUVLFVNvI1nbXLq5HApAZ8CPTm/JI115j1Mwc+qCg4sKun2S/1ZzYV+87b54aUqK/rMnDh9oiX3
gjcqwJTgIPUE3XAAMDdaE4EZ4Vkp8302mBO/I/bYR/++JJyw4rqzB7s5f50BVHygSMDISzSQYmIi
8z7MtP3m/Jg+mw0OVqDw8jl8saZeqNMPfqPhFfZ8Vm9LJuCFmufCjXjXeFG1gQG6fXSTt7Sd9g0e
q7RYbJ/ODOfllb4n93acJRCEn+cwSrEUImwoKHMs11NExjIbpIm6qEq+hgHf5VQ7QUGt6v7tWkVd
bvaZB+LASaxRfvCzALtvRrJyMqpn+ksaTG8QfjFMAkcasCLOgo++39xFCaPrhVMGWEe3yN7PZ5I4
1IRvSwEvBBWGw7oppJwdjqb/REMz3iVWPcckFRYhGPK/JumzrXMrr7X4OZNFkwjl+KCxkwJRDYrZ
F2ETJTE/GX/I+lbNsdgTTVd1tz0UDt3TDFsdE/t3YvwCRSO+mltt5vvo6CrggfaaAlYarEru2Qsx
/JLtZrf3ho/74S7jey0uUuQNwRXoW631ZYJ69MTmRSLur2xMi2lFW28n8Z3utTm4bVblbTAmUal0
x50aYpH7cYBSTEgS2bVEbaetwfDME8IX2h3AKlUjTL6mGbWHarnmftAcukZXFnKFAbU3Eqxr4rgj
wwHIZLlOpcqqlqHGku8rF/ENj1ojfIcZKMmoofUCgnGAL3XAsHXIfXwF1EZCnA0VJEhDlo1bF9i2
Fv/G6/vBn4cJ3ww/ZTWJib93PbCykM0Dp5ZBwiQGRMxXini2RWpsXJGu0j1ixpAMOzs9kaMR9Bv2
ON7NLTIiRfCM13YkT4Hj7lbONMq9IP/uwQyXJXyHk33z0zhNRQpqLUaZQ6rp8yoMygmUSaGhB8Oo
hiEoofQ8B5XQolZx0ANh7ncYvCVXIrkp9c5idkXN5uxrTnOe6Y/jrZcfd1TxW+dHdZOZUyB2qpSi
e77XhVWmhWPM90ynBjEZLFQo2uFESDgLhgdnv7JTWYXPvPT8XxH6Ya4a736+yfuz0J+De/LjYCFk
pPd2g9WHp8S9nzUHhDk45gTMOL+q7W1dd53mmbAm6KLAQsK9/eIm3eiH6o+6PhyNOZtnffM0EaPu
+a3941VcrLxdgtJR4F5ylWfSz5SEAWKH+JuX+ur6khDSHU4UaMesNwTxUEDw6CFg6JIjAUIhpPGx
c55zE3kulCpmKcma0996VPQrOf1pk5z2P1Koa2RyQTP0AjnOMlo0xtN0oFMd9G5u/xobfZM6dQhs
KJGG72g6XH+FiJCHpStfSc4tLYY99cHXY7vuJ0s0IlTMIf/wEz1uOqOMGyzmL96/lmjVlSs7y0K4
WNJ7C4ZyzCgXodPCOnkERMAKFTrxrV1cW/LPkue4f9DAP7Nm7vShpdJLsj09RgLSCYDTPipPRjPX
21a9are2rhUPUZxVtl7naagaz8xXlvb3IpufBZNJYc1bHoSZlRDAE/uU4biZt54bj3Tfx6gNGKr/
RFigG5rVJw8jmrdzqN/tJLYVbOxKCbFjxQVwrxZviKNB1M3gbVowSshcTImy9hXzYEGO43yDrlan
phg/DB6qs5cB+kABEWG6CFOqzc+8T/LafHHK4wzJ1+TYkQnZpIztaSf3jqewv86cOYxHBaa9GGNH
aG/ZNA7e+Di/Umh9LPtVz3wyZKvP9y6hrTEuMl7qkVMNC0opyRXSHbnYeutMUMJyFK+4boU4pFB+
oj6IpuX6b/HNo54tryvV9/KawLcITiOxlhQeUjhTrXDqSmiGJAhmYLdxttQbjW8zlnGU19wGUUrB
HSPGGezUmxkqYVEwrZhAkDjWN7/6a4F3dEA/R8EoX3DEcW6JPQOwBCDKqpAX4u/1mj/bYDKqZaaI
lvGmt+sbZ0gUZTOC7Ntjn7eATmNdBNIGZRHfpkpMQfxlbE5Cf9wazWLJ3rGHqBpBs0tbulL3vYVo
HItWDj07ULEDLU9bLkXtuLdhG/xpZaozHbZtjB8QusU35xPtpvo33ewgomPnx/dV4EMtHttCneh+
O/MUs/rS3bp1BpZpgfNz5GBu2CHTO0f0/trpwBI1siyM15RxBn9cEmFSWMtNCA7Cd9DxAEiWuPxK
0wVKhnTZpYsKy+wd9pHk61egXCCPfmAlGBiTJzGx98hW5lR0bNX7bTyltpKoFps/yi8BmlPKonQ/
jW9c8pFA8Y8qd4r5PVYkKJPSLDSM11oG9TsAmoWyK4AchjyGl24f2tZtVgDsU1fHUryU3e61S3D+
8ju7SP1N7SiSubgT8NeeD6/Ww4iRKsn5KRT4zWHI7dSHJK6r7tbD2SS6hraNSRhBSQxijLNXRE2K
+Vi+K8G9DVTkZKw50Rzy91WcOkT8+AgKPysIN+o1Nqo08K4ZEjwYOxShFvTzYo484/KbnPtIqXyY
AKKCqAmrOKNabYALfZeb/DqByL9tvq/7dFNnKiCyoIOmZbHJvZSCIS4bJaTBc+ygTU7IidEtIegG
Ipu9e33xuTVd1nlWaQ4zthPcb4uJnrOb0Bf1ZYG0RXNU8On5jwFQ3mAwKlUh9uxzQHaLdVgPJNiB
fp4KJ8mPjDlq6Xf9IOZW9SZjACf8jedbSl3nmu5br3tvUcuhAbvV718LEkTqDWjHCaynQx7rP31i
9GhzRRfkGISElqkxJr7o2upwEn7WN88XWNMqieC1LSAI+4BKPf6+qUJr7KikCId6KmvQHD6DVZVL
SS29vg94MQgufXl+v+k3njR3HYotrsI9akGA3/t6bOXdPmhag0XpdUCjCE68PIv5+KGT2ierAvKD
kgkdf9LJ4t89K/kPa1Jkm/QG2dK4OHML8+xO3jMBm/Nk9+pd+V9WyK/KKX4Bt0hk2U0gy8IZX37y
vjnuKkgWzYj4LadMWq2ok3E629m1liRZHiJGiFIzy3ChRdDrm3gWBCBoEkFPonbSVOPQnRESjqZG
u75mmsk8MZ+bhOigq8rbR0SkV76N/k6mvO3KHJTw37SccHKSeL7VAFJ6jLvc5/dIuDuK9bDEhzXK
J3XwiZ/U6XPeXE3SImeXD0un9ghL7PCO5GMKsoLj0Ja+jG5hozbT13bF2ZJ4lgpssJ2FEkMLU+6f
pqOBJwrGSqOmL1EkkdfnH10i/5lcw9WQQNajMzY61SugPY8XutnR3iC5mS/ROQTyACEzyu42NSfe
ENFutfDIAXeHaake+lgiwskAw8OJQV6PXBvyQmt3oaCR+29KxRXbb9FNMjSVUMawb0cuTrO8RgeY
29dueo4kbysA3BzIz/N4O9o7wZ31saWQHmPriP0OTe5Ma5SMqYI1wzXD533SqisLVICx4ANMuWs+
ptzqV8MdC6ICQSqvoQhMqiwV7mCcLDQCeXzCGt4lZqK1IegSCLe4/I6Su3i63xa0jXhNFtNSGrgy
c8VYLsUXgGZ8H/AsjBkDXxy4J6vIfEpRRr+HUh6bx25JIc0gXC7sLQDA2mbQXku+ppgJZHpQ7aT9
Rz9+DDMizrpHHMpfgDdSue+WUlM3xEkRvnXZhkgIUYocO7ShWgzrfiG73G5jmohkFWKp8Y3+Cy1y
8oztB6mgzFWIws0K4fVvgQJyjhyggg5F/TMXxiKX1VIw8n3w4VgNVx0Cld2sfiCJunXeM1kerSLQ
+ELK1CdykN3noL5HiUS2YWURP7snPy5JSQUtleUJoDHTIKb3DafVPz5f51hehr1AHyfma15m7qDp
oZW+EyUQ22MlSAX0H+AZIWGm5WLZjKmLlwmUYvMZdtk8hDY/4+Qu+ISULJtzJdLAKMCHUvaF98Jh
fJPWE9UB3iTIta8DYyJOGygr7DfMRodqnPY9Cm6xoMYnG9Xe0GQ02D6nC/7qS44Fa7lbKPjcobly
Q4ko98Js23zEAZAM0iIlvM9e0kaftnbP+X4u02ekY+mZzv3ma1+RckXUEcIr4UBIzVyzOZcjqtpc
Fs248zuykWYIntoI0iEwQ2YuMXcEPPPaixB3sRtX6q+Buo8jBceR/xuqCkzccCzW0irqsKUnlT+l
LzGey5O5mxulfbipfFALTdcLQZuRWg7jBKL3lqGv4px/7YpkNnkI5Xztg2enOtG+j4RW4ma+8TBP
PNbexWpE5ZWnhP+9g69nkpGhQQGIJAVPuw/hs622Pf9awuKnmDLSu8RVFxhWIOjzgvsGFAclVwI0
nbdYGqkILkqWbO22yl/G/NEmsEnzIrvrGV3wKuOCdtAfnjhYl3p33FvGqVIqwpuCCeAMcB9CDumj
khvx8OCc5JBHmf8iJRtUnHaM8uuUO90W66p/Qt98iwV+fq6JMoF9tK6mNBh5oe6+o1gXwQgT8Wvi
qpBUT4DqFHVbJlc3zsdza7N3u5FzH8xuZbz/NXYoBYBAAN5Fq3lp2YYSfF+dP0DNK02VsU4f3zMt
RnqYX4qsQZz7G8M33c9vn7Euh3vuEIwapsj9OvkvCdzbVSIkBo5HwzYC5ESTqPMR4cA9HDf9vxFJ
HPpCaYN51qE95DMbpq6m4OU0UKNPOMXW+2trNaRu81D19iVONGU8WoBNvMBSYUr5elqjHxynXEjP
+D8zkEY7K/WPFhnhBdalzhzrGpkQ7wpdVgfK7HoD/zsqkx2C8fHkmJ6gL7W7j85iBNORMVKFUrnz
Sh7fPO7r3nejP9y8JhMdGw1dYRCaimPkgBTscZXcvUbu4SXWFA3lHqVQUweSxFivdgusAu3hRl+p
nRtGC525u2Wmqn0Bc/2dRTZStB5IgmmRFEzH5T4B3p/Xptlu3yfBKCkMePoOMa76E/Ll0BkQT0hn
yrUyybr3sNMRHAEOafzeqaZ2sG7O58YiHpzGNoG3A/Ta22T4x62kA2sl2pGFUwe9dtmBLv78hjQu
OO3UAvgE8YVO1bY7C7Y+tPlUA331GAUi65wDIFavFDO6CHuXXYGo8Le3iD5khB+3VXqu+Z+SsgBc
7DRPLzsf//ULyfz6EX+1rMgSJ1hedge1lZpnbidLZrDEV4PMQfOpH5DzhQw//q1AM+ksn0JdSWcn
ztTHgOQjdYx2tUm5vfaHQ3+VvEYvu+Nl6DRr3dxgYkdVEdqHq+wydJcCHae3nHIKmfFomYR3jPOT
IpNRww5zfiObB1c1lXwsGlKqEWRV3zdbElZ+5uB2v6Mr/8/bCVN8r3l+E2kMpuSMkDjH3/HGTbDh
Dtrq8W6D7Hjp3zPKJFaJ7SYutqKtjqB8k0DvjBj5DqoBm+lEtbYaj7ddGhI9kz6I07oecZAGH5TB
iYdxlxqfYVV3Mpl9WP+2tTZk6ooEApLR5RQJZT1NF9plvXBEmjjX9YsAagG2DJLSMhN5NVbTf+xI
e5HJ/PG8XKW7u9JlLAsINOu7WMC/5gYyGfJPfQPz52FHs77eCwZtpipHvvhdcxkz/u3utvUVZLnl
up/3tuE3oa0wMS8VIa3yWO1tJfxlXzZxJYTXjm2O3PyWij7oqd9+/hwiz6ScJ8bYBApZkvYQvi0n
844D5INA8eunTIRSVRVKqnP0Qu5w3lYDP3oEUA2schE5cLJdw5SQpp1gimZti5fK/nzBS9GYsy4t
rKrQbfb6u9CNj6Fgqc0yFf6A9SR6E1uK/P1sq8mPt2g/8xRC74diSCgR3SbN14WB4QoWGb7HLlpx
1HY/lieqyS8l9HC+SI/CbKe70lOAxxJI84YyCjr3dAfaZZPld7xLSyxd1VVIVCAwRrSFRRsqa9Sz
j1bk4QjASJVAIYwqNr6yhBBX6TRSDP87FtIzFQySN8mrHwzJjz/JI98njVwRlWKb5PdA/2lROXDp
kwKTVl+rWFaXkvbAw0KlNAkYxc1AwnJz3yZFLkTzQLpqy/24txhC1bW73bRh7aMQIcBF4BE0kxAn
YiirdUEBpkmaO+cTWx+pvA1axzFBZSMU/tvQhq02K4JHNQ9XD3ygO9DG6ov9ibPTjbGcSzAPHA1S
UxmTGMgpApOIDsRdboEa/QAffVZhjwA6kDltfiRjEo9Vo6pdhS6qaaKlOOubD80o8vX2VmXvyiR/
R3T7N23rD9X2KuuySA8xnjYGGiC090lHbXu7knRdTCUmsFYFFBM+sn8gRGwTcBd8KVrkQ7J+QO7/
N7M0IrbmcCIBNMUczrZNUt7+tkkx7Cu3uGwBv7VlINaKd7/AC8EeI1rvip5JYd/DWZo2DeCz9G2q
DZ6wMrlklT4/UhfPd9AfxMniEuwMAXwquHZM/B0682CsBCg5ejaZJ9dKL5nCSVby6sDYQGhiBefh
tn0xZSmx8F3PA/zC6HXLPnM78bizhdMn0ZLdblf77OOrAKlwqz7IRji50uOh01d+nE6kZSn9jX0f
+7c11Vgrb9fsdhyGnoyH4phFYDWa+aNl8h2oraYF+eFuKbmBYDzqLEwVEtjR1I8DXvndAu7KTQNb
Bd6XQ/wMg7SJUBuJwaTyHyUAajZf0lC+UZ6bbeDANo4MCsQn2Csck8SBuMMLvdnRlJ50BvJWhlUu
Qm8BcSg/PJXG1U6SL8eXIkjNC0MQSrJZxlYKQbsxcaFsChpWa7S77jQAHeN1BlTHUhmjzwjpLRyv
lPajVt72WjLdwvDSXHKMn/QtAbxTtvsEIQvn6E+WOver2/TPJLjXsb9XpaGjt1tXFKnL9xo4FWY+
m8VvmSTbcE2NPUZuPrbqexrcXcasiyOdmGGWxc+5cSRZjokdAw1iJyBLc33U59sOMWPvr/ATW5aq
ss3KQ4eP/XDXFJLF7QRAEq1sgHWtVoe7AA7ZC7VHsHIOTf0ne8LbXw4SxhJiXVuqXU/RJQ7wA5dd
VzuzWXGbRIfxpPoJEAbjj+UiHxknw7mB1cI52dKPTkNaA3bAPG5SGoVe2oQ4oI0GJH3AStUk+j/W
+e+yT9TuSmQHUtVdMeRdqMRRonXWmOGxf7BKJpU6U63hocklRktxOI0En6uzSWVGS3+cODVBkc/V
XAjZofV2jPWnoaUpBkjuBmBYhcs+ak3s9XEpNisyXmbOo3aez3y8SGZyA4u8T+Pf9iD8NH86ZPJh
92aSdZyu/cStS/aGjBVVpKyaeyo/3jTL0tedv4rc7AgBHo2lSDIXd5A89jsmVn7qemHAZW77VwqR
F1luzcB2U0fCQInQ8ZGeu1GT2DgqdncAZJIm7BQcZZ1V2akj2oB1CjSZxO0tQefiY47nI0SOu57R
AWrV9KlhpuaSyATCRWPddV3qQ6lRsLnArYylSA7DkYGrB/P/l/h9BqbGeMEEUN4hSRO8eGaYzYPA
wir0KpOaBbHEv3nXSVaDIPCas+vmhA+ANnDyb4fKimE/0dKN9YNnol6DrYju63ZqE6/3ZHXzCGxq
YGOiz00016dwEhF3owD/Qk8ORKxi4xmjb5sxM0Vxo/zAWI0VcpxHtaNMxVjq83sGA/PsL6XPb23g
yxJZXKWVraZc/uyzQvnaLp4v7z1WhIGjIfCxHydVNlru20uToXS9S1rZ6jimbHV5UBdzBsO0AOcm
AOs6kxLIPI4ticRy244BJuVS5C3gtl2jZjnUEw6ETqfk3DdVI/ZVTcugSNtTVicN+cjEtV3EEW9Y
WYHQXEFVpFmb0QuYX5zIEzZ5hY8gk2mykVFH0NXWVWHaoWibi1och8WX13sJjkWt8QQYbEcr9cwY
BXCWpq4BlDpa6vaQ3hjOXPN1X7I9ru9AeNKfE+SZw+3T9qmfCCCVzY3rQYMbECxeBjSq3jDO15+4
Qigp4X9Bsq8rO8fTLDtRM/oacwFdaIUdnLHnu9oOt3nEbfAc5pJTMavxLYD41NIvXGZFwwpPdkYj
1cQXnucaWoauf19pT20VF+vqWYEKJOriwLfaXTPmUMJ+LstMIqb0yNrijDLCAeFjhRYTR6AkfQfg
3n3G7AiHthvL7FhOd/a8XMhnBrnHVsR5SGBOnT4s4UGlTiRswjmKz0ni+I91qnOshqxDehB/J1y5
SR/AGc+uLMpXgcJaONGJB7hw8G4Ar61RbiK84W5HwFx/bvudGNhnBQI8ENPXyAzN8pyAQThAVPvj
irZv7LF4xHSeYYXDHDU5kb+EgVctWWuKYJiP6X5phwVVeL3ekuGs6AA4ecHIVwf9thpDooZzLxx8
a4M8VVky/OrcU+mfs+dflV0iEhTcAhP1ZYwtDl9UY3946AKkpj2vSRL+T0fzxyX3ShyXDudLOTlN
qXMNveZcKTs5k6tIySe0mz3lbGhk74hid8Ow7GpQbdVqxmJM168gu5pmVdZaPG5m0WTGuHlgsvjA
TfO4n8gySbqKr+KSkHBNYDPOcA5Hjlkbt/s0sVv8038vfxx73RHXelhP9bXP+svoMmVezUMP3MwZ
l2ow4ED4N3NdXBjn1rCoMrWBVTocAueodYRro9Ctr25nMntk6LhXXuSqrMsQbfUzEkp8M4QVquG8
BeKU2GGc9VYTSTPAkAp5JoQ1+jf1F5QiourWC2h1WYCTnPYreX5cu8U3hHdP//SawZXZBU6nLOBn
qVzqiFtrbWbGO/A00obSpf78PBl57FJZSaLTUa4hso7LflYke+1fJ2xePOhkGA/9HXDvMlIUVLFo
9HeP8hK2nu9ASIp1wnuZDTq5IDj6YYbcouYVhTlIvCvFepGRtO0MuvGalmRG88yEKl4OyKTo9v1o
bltIUSmk479DZnkgM3vtwEuUiaMb45CoufKJZffiKLE0JeaQf3RAEaI4XStXj838McvhdHZPjvjr
9tam7lnVHxMCFfrah9uO2TSHO3b22CoU8kNrVS4FtsCBNx70t1vP6KSinvzOl6d7fuwGVUSdpdBH
rpX1vY1AWqIfYjUHNSHS/WPiC9YrYHH9sayOTbKoeMaP0yzQ0rfKFnTnGoMxvxWOuZFNOOt+EDQj
le7uNjugmoHN9hevmuBqNbOweOm/MIVkoDhJkh/a4rBj5VCrHrXHIK/XGjMWPZfDAgxSLEPKN9tW
WBJmVB41NLatJDbBfGOQOEZcwlS344NiyeXrYxrSCyAM3wUtjp5z53UBH5gVcPeEafgvKrG3ywP6
6PwPgj5gWfF56YSgPwlQNYeVAd+owFLYyUWaCIBeAfsL+uMR4tNpvi1ioQJ5R+QqO/f0QrQLGSug
93zNV6FGWlArqoxty3LvN3/niaE2auFe/LI+odZkLVQENQVDZFAexYba/KsjI6x6KYj16ncMEbrK
vMkJ3mj6dcXQiFcVTg4pMjzJHb6Au3gP1gHuNG8kNxR+cThJYptfZuUkWf+rxBdIxYzK6P1eEy8e
b4mSMtQXvpgU0OQuL92nJk1h8IzXTC5uTlwK5C5jJ+YZkOFacXVQW3rBGGrOJSZkVZdtXG1yobMq
nxjXvnY60ayiSbzwidC+/bZM/UtD/BxSMhCNUe9ygr8JuN50qoAA0SaHJ8vPfs3XSEL2jOURddmo
vHpuFfiVU6YB2kAl7fhm34hC8MAbltSABrMoyTlXECgIdm6uh4hNoA4DgcQr6yBe4MoaEKMCHP75
a6UjcYDVYrRaQdO1throfQSHQwPuw797b9r/wVbOtQNidtdwvBcJXgP87wpY+q+1DjWVEeFuJFNj
2NeXAfnm103EuB0pwak4WQQLf/G1wOl8W+j4r9q4A7orxexpIREB/e+xUk0EYT5Woyl82QVIR7B+
zu7DSUzAj3j13OaTPfjULU8i8CTij+xoHk9+lrMnid2wqZb0NPE93f1z/5xYZ0ZCXB6G01+MzVoM
jntO8fBEs//GhT6JILyWYX9vBtL5N7jH14RVcoX2x+L2b5mzKqBSpIAJLvHIKp3NmmnQvUVkfS1l
CFtX7442P6ZFxnpJgjsD7RECz31IAelOrdmIrSl+qznh4tSRs0fOv69i13P22TRVSnK+ostkm2ws
I6gclwFwcc/438MwJOm7MvF6gXMrD9MBpGoTb7UotFnHg5UqCV1/PEvLJ/swqW2RtYtscc8H6Grl
YC+W4t8b3jC7fRwd7rBn363WFs9HK7am6Z4A0UpxsQgEcRUsQHxuwu1R1lJazBP7LhPF/z1NTP4c
OJB1t6F069Aj5vCGX+23GRBKEZMRnXjfK5WRWjKSrL5z1btbZv+dkFXIlwea+HuRDF6IkcBuHVWr
ckIAkobYNi9tsz5Tm6vsggZ7y0+RdUJFJFZRk7hZg0a9YTD/cezsUyFzhNpBYhTch4fuqinxX0u7
I0Lz2hFcKmPXvJvqCMTo++vxjofyRsw5RJLU1IyYCiWe2psZS3izquGLY7CWHABQVngvqCa3yk53
uohPug+M5qNO/HfIrPSE6JIy/uu1A8r6EiYzJZoT8ij/d7Y3seZJT9PvTpw8bECnpHNZwe8Iq2G4
qASXV7phdT0VQ3tsDI30N81T3yoiWLFPbEV909f4Q9PIJKs4M9YmDVV6OErJpEhiDjptZy37mqAY
gieTtnUElQ6JaEdSczTG81PYaxBRKMPg2Y/9zxIBLROemJ893DNYTPhla/Z7bVhMF0r8FbSfqW6A
Lq/Y8AY2e1irgnaIoGyXhAYorz6IKv3Uf7580JToMVFU8uP5rpVQzvE5IAwafxU4hONzn2rBKNbj
IKh2Awr5mzsipXlhTM8AMNHxLxyzMdhT9n30UEdJAhlZsfHjJEfUPqWbQcN7RQQj4QuVqbuZEoxl
ahiiZoOBLSI9ZNhr4+9nqasHbhNQctj/PVOQLpXbdzbjW+9t4dhzvRCk8wbRMtiT5ut+im1NBgmo
ptOV9dDJnQLrcliOBdV6Xdb40FHdAsWcSuCstfTak+TtnQ4XIsiSaT/EvLoyFZEgnTmEn5pSITGz
erMP7gkQAiX1l4IUaK5xXJnooZ1KaUxX/9+RrIkXsncXDETSEBmrIuiCz32PaUadL/Z6OdGSC2Ch
hNeLaD+s7gvEjrOrQk5UDW409XQbP0x51ZzKFqOtXo9+5XlbJJGH/NNYLfpKwArdEAOVaDF7UpNR
vvhso4P15Md3UMCirwQRB9J7AFqflrNUUDVljkPLe8RICNSiWoLVtVB9SEQbO4bweNNRbSucDuGm
+ufBe2jwev9I0t+hoxJi05VtBw+zURe7+sgtjQHDiRZMq2/520+wk26HzL8d3h1F5w9JfvPOS6sL
pdg1szxANVEGAwqKd0OgzZCiTpjPGhvGpzAK7FLiEXcmUoEa481RwkK1t80XKAaPFZ+Am74uhN/k
XH0UIxTzPJ0jYRDudWzR2UPyjQxEZfHAsn1VX2yONGqFaVLsWqpL8JwSLmC7PhYz3ayGP4ClvjjH
7qn6HdFfA4SeDd1OWkeWX+a3ippdu67hGgN2VxEgqJIJlOeS5lt3YfQvr+TWmSweYBu/NsN5zgJY
i4yt2bqEqgmRBGq8FWKX9YVoZu4JGw8k2Ehwx3/a5AHYNfeS3ok+cGSdScxLbJ3ZQ4gnEvXcuN9N
v/syB+MDxI6FMDMOjUmIrIhxNA99ZBAQsinp32N+/T2OdGneRDzcDiPMKfyX7xKygnWEqakR3B0d
iW64txXh7pcHlFeeEFYhjbwhUZHJDXzhyb8+g3DX6wXQD6O6+5kf59XT8J6F1ma9bbIWfDbqFo/J
0G/kjeYHQC/JU5S0XQW+ONiqY8yjtYzuFY5vbpJbW22d7qjE3sbBDR5zx05p19TpK1+E2FeAqgZF
KxlRKAE62sIfYRaCnAVUUUuAuaZgJt/JDQvbE0SHN7/AQzNfSMxmUC2qi8CLlXEfxVS32Tc87L60
NMGpojlZE90hRSEDkpmUUNG0XsFFbcQ0Gy+gO0glSyg2EREr+C9oQhGjg89UGrEAAyrwJDt6xIIm
pWFGdTTUGpoPC4o1MdCHfDwL0VY/ykk73fcHJGB54aEfgMCUyigd3d0OW+pEvsHxI8tkAHJkTnrx
4jX9isTEMGkqm5Jg4y6J/LeOde9RjSsdos1zKWOJ+e+rP7E10upwrAIuxqDL1rFqQLCvh8Ix6gMV
fesOhsxU7atgOpOcbrdtjZpVqVDbDJk+Zmf5FNxYY6DuyXF0QKI2POjvW4eGsFhy32ak5Mgl7/bv
HWXIY0t7v7RCGexN2JcFipmnCVgrQVFZ0E2Dibaiflz/E/cF4f6GmK+zROAyTmprHStynC8Ffra7
9xFdL0oKTlnr0Wif+mrfHr2IIOGX24SU//yS1wQexmvv9aoAR0hcRlFouYKYLXhSIRNeDkVmgFCL
H2zysE03PpJYrRlPjUK+9wNM7Ql685QM8UqltyOpKr0x+y1UkcgrEF9NXXusPhb9dsMTx6qgcJQR
sec1M+Tvqtuh+d4qZ9FHGVF7BrPP7eclsh69MvSZ2KwhEZzP3PfKesfBVCekfPiTQaV7qmCkWHwj
yn0KDkU6QV0vgh6CocB+/1FZJvzSbMJ0OSE/m780CGstnBulrF9ElOigRstCtwtHxolTbw9ILAy2
n67fk75l0txL1YI6S+LkVUxu4kQE5hR4KKC5VRlj22wrSkwVWYhDZTS2EyA9rMN3uuzir1v4JoCy
Q+akxf3Y0RnIx0p2R8OFAV0o9OlKsgiLIFR/i0HMz2D72nv0XQSsLthd5eP6itjx88fWa0ozzfh7
rRZh44az77U9u3a7sROg9sDUrfJ38iVc1EuRXQBQvzZNoMmuSbf4xLnsuGeK/9FCu7b6C/jj+P6v
er8Pkbavf/GLEDAdflG0JAcqLGqfVQvDmLKoxqateoHFky68EFtwdPc9qv52KQPLnGl0NFBYXH7R
rObgnrQvYe0ONKRBaH/xhMF1+FImHE8tjzaa5pKRr3WJ+OkBuh71xB2UYEBlxkzjSfb3+vW9EMsC
dRrERIfWN7FcSfYw7IlYvZNdbOHVkHT/qw+hoWHe+M3OnDT/Uyyx1PTgsF42m8Buly8Kpg+Xqw5S
3UOo0Kn0bVRNzThnYE8vc5wL+VArwf+e0nxqnoGPtvd6srz/7hxbbQfZjeNXQr6kc9B0Yga3VeYR
PavijUVQkVduh7gY1D09W+fWZu8ljGzrwBcK3Q9E+hPwjRiGRm/MFN+Pz/IjhxIlbkdhYuMDtue2
w42fSDW6/duPbpb5KRoql7ixiPlHDWAZItzWhKJvxlXNfCGOPX56c8LfuO6h7SQVZ4kIkg8Si8id
Yu5K3NSYj1fo9f+gmi5jEHff6InosgiCV5PGnT6Gye7rMvy22imzsLTO71jurCKiTvbCLymm0LtO
te8e+nan70U+DZbtZ0I45lBK2drf1NSG7jZz2BS9kK9SXP8N3Ea8Y/5DfE3xL2XM40EcbJ6vsmBK
iKSePLAUPgHhQOjg46Ntf6pDBfu0QuzbeMJA1CzF+e68k0m3KBPAv3oXq2FSG1HZsj9DukqNwWXG
wQEOoEIdUKKOQ0+0C9njSdMLwV9/eNs1hvoQ+GT80Da6LyObS/aqteQQ/CR1JRsY3bGgApAZdvNR
pazQN1+bH53jHnYv8PE5NKPX/qvBNpX6Mdjh+7PjZBlmnIQnKaqwkzi1CHuSA/zxb6jWuJ/+CATi
C6PtDyr9Lq9xXIZc8Blvd4zSAscdOrzg812QXRU54BpO8BTjAyzVVSAhN1fR2ZzzUL/h4AHzZ5cp
oy5k/H2/R+ROeeNvKl1q39tA2VW9coe9g2zwBIgdQAbEBueSgmBgGtxKdwv8KVHUqLgmYTvPpAjW
JpYs2UvWAACQP09hc0J/zVqPAsrUo9UbHqA+o+RbKFVdVA3/Cd8P+gaOII3b8OvVXvclqyePKfpy
U8xC6FDaNOaQtGBVfB66CthJgN+hCoA6iBUrAY7xT2HECBU4cd/oo814HuSpZsHj9Kj6xrB0c2bt
58x3vGZo/XsYilu4tF1qsGs15+RosbGpA2YbxrvME555ws4rPZCQZEHhTitqd2Gd0YZ81cfwAc4B
lKUHP3oGmztNq+ESwtfeBOqZ6dPNrQ0BU7/+wgrXIU4N1JDiX2h4ZPuh9ZJg7kawZwnz7zjg8oi/
1gPFAd8UAMaYpXfOnkXhbDVjDNYU33LD3NbC1T+dezc3v78IJiT5FvrvA+gx0PCorF83mY6l8Lq2
BoJLXBCb5CCIuit8k7ZRpc2QKPm0B7o5dq4EhvnrfXOzffms/7ornq2Z0eSIPOg1RbV+/NFeDx2m
njpC9F/9lEsxlWB21BVjyxyoazBhccFmMUMUpnH7IEEewI61kHT19X3Bh9CreDFTrjBmHCJWQs90
SmU0bqjChWiyl6YRugYAzabJK8Zc454RhMJxuSEJGG/p3eB5E/sAwZ+clO51iJ2GLHPtPaWTZmEP
brt5PlsNgpIRrJ33cB6rpclcx52q3GhcNgWI9+u43R0KT0q8mjK4UUIT3Q+LZ6oLaDeM7Fq3Fkho
C8uOLaXW6LXmZ1sUQ0C9zF02Rxxxo2hgNPXT6ivXlgYIWo5LlM1jXRDyf/K2RqNOfzkLAsDUXjaH
CN7K4m8AR0DMxD2+Hjjizi/l8s5E9/AHptgznb39rnjGI845+3kxAzOpTSj/y+I3aCpP9hYfW5rU
cM7Bq5D/VgTSAOdnjO/JvXU6zXe7owoiQoe6vf8Ah+55KHTbB+tq9Qjx5ypIWo90LTnEeY9ooKrr
ZRyc6rCCnuG2DIoANH7T7MTXSrRD/BeUjfGimzDH5/ByWlcIut1BeVEIRT1GQowc6roSUGeXQ+/q
lz1/KK+piJFyar22tEIJX5bQh/WlgIjIPLZXllyf8wH/9cLMEXRNP6a9kfCgp7luMue/Sh3Gpw1O
1eaKacYfTf9+kG1jUq71r7WvAGiQ7p+NCvxTqHLMqlk8bes4Y6zH06zLjYTAqidY4gB3wOH5OlG/
u9KTB3S3dIzusslnYZRAfSuikrvmiX+pGR9YZggyW7E+lNYJYP2WDQZckI6L6E/6IsMJeHltpQrX
32UtKwT1jsPaS/iwRtpV9tsqEYOCIP4wHi5X5XZ4ed8lRZTCuouuWEshSpsCOeBlAF/I2DmCZMf3
Gj2mRaQAaRcFUrHq5I90Hz8f5/url9yyZfGE/P62E4XxtGUVM1dTs/pdVdQrXJL4CLTFusE1fY3i
nuqtaiyDAwHhRgwz95xLOWW9OXkb2J78k6962GmBd+dia+zRgsJOJKX2ld14sNq6TXwamHSCZ2mb
g16gas2mHcqA3ETbChgzoMhriMbpEh6o5zme3mgUaMJsOPRfxrfH8u7VlL9OZorX4joyFjl60d41
IB6g4LN+nYrwCPWzjn60VCTHE6fJn0b+L5aO6HLVAz7nSe6z5CFmf1GgCGwOZjOPCN5R0hhIDG+V
SGM5Rm4/L98Uk/33EjXdDvgYN2b4/GdAg/JPkT16U4LXdDCzPH6PxDZXI8Ii+G1kjuxCzn1+2v3z
k2fHTF3HdsU4T/kLdeWdeVAjXe47QR1SB887q7Vp1rlAfsLAYTMxrGQJzBlY1YcrsrXr9vPdGHM6
IlpS6YzdEss+dRr9mtAR0wQmJCwaaMJ/fruNgwxMtB+cMpxSwjM6M1X+Tl0ABQbJIXbYdEem5Pyg
vAO/r2zFHFvJKHyUscDiQAYJPR8vLDfa44IaNA7qxv8fulHDcsuomRg/8BzS5OsFXOd5sEMNSjyd
A6ptcQighkCk5U66wZgWgXOQG5F5PUdyrxNjNq4XKDwlOoXaPb245Y5bUs1cPJq/wxFfjtES86I0
c8q+7PnFebHbkhcDLGBbwCD5aFZVBLrLffuOvcGXQmzj3PeQ/4F8GHxUIhgXBWM58lh0p7cuJSmn
qbFQZ6vOo7iXwB96lzS62ChF3uENJwVHW9gzebRdNtW+CNEXWExZ3uqABpUbKXmVn2P6PW8dJsa5
myQdCyHzcHTGDaHHUgxWIQjlldz1jR1Y4+b4I1i9m2WNg5SfzZjm2f5+E7e+HgTiZeFJxmTvfqkj
3XzEA6Mbc+tcqP06riGrdGhSP6sIcaPxItuyXgpX8Fc4F3KfmWAZXr7JBJFPUBQx6KpZjzOpgImC
cJ/YGNVJHS+Chaal57LIUvxg4v699qSOXoiG2Tl3SabrQrWASghvBC1iwsDFgztjv6lHlbKJmhM3
MuzPqbqsxcFofpNeVL4doTze8tRbLcu7sK1gYm2RbuF5/W/jmMGJEByM7zd+3ridl3gZaiu+1Bn3
pHu+nosFnmLieG9NocB7qDjRP86Qzo4DO+hu+F3CdjmPPvWV5hbQBqvfG/FfyopMW24ZM6ZMDPF8
a1yXrHM0o6iJDfELNUr4NYhE09j64YJv4ClIPxNZn45aO2TJ1W2mMPJy1p9l9PM4qxf6IAFGI/bx
LeSTSbhXv6K28ZAbDy4AizxzOMrFqP+0LF9zujKm6JR4p+i97bZ85Sqx1O/LPmaRyPwhxKjVxEZl
L9+yu2TgI2g9AxRWq8JNLllwVcq0CnPYpRhUJuP9PP+7Y+dBS6HxXaylbfQZZzMOe6xpeYc1kW3t
nNxjX8w+j44ycCIoWPH1Mi5G5jUfhBXzciRz2d0nE929MhJX6rLJEt6spKJsO7jcnVH7s7xf7E9y
Mb3PXcnCufnR5HIlgqoMP+Y4BcJYyUUIPEdzoNl70Q7Dj3lpaoZweQQuRHwi/5r7JYljVnbzQAaP
HwxDrtzHirsSz6XCxZupVlXhYJmkNwonQh1rrv7PZ62WqRvtIcjTAgK+81YSxkQAVTg3+l4NZ+I9
Sqdix8TAcpPgsW39uexeAfXV260wzJx1hfbss6MSTcoWwHHZRCg5OU87DZjo1+k8mMkOQ3aRViF3
SIJNstaJ2Gkr4djBU6J7hZkfxuqusaCqWmlhmM/cCDIXGRL/dUwhBBGnrXRGX52Ob23Tz11W7kO+
rkYsT07Nvois0+KInON8GAudiCF+djr8Cf5N3Nb41ooB6aJBOo1t6a96WHGxi/jagKKPbNcO8VTE
fX0e9DtlWhWxB2Ob6wFEbxMYlQTzhWKJwlOR0Wfvt6B4YbZmEMh36XyWkQONvzOKuPPH1nVe4V8L
89mctTmZ+TPciApqbMxZ7L5EMXyMFOUjPytuMwYvI1BCv8N6JFbCZgsJhIsLzZ3qiCL0Sg/6eroI
sNBekRjh/o89Qn5mY4Vez/Ntw3/1qyfqtiEZuPHrHRdZmRV9I3NjO4nFeqTmtCaBQzcGpIIBL0DF
kyMjLqjKktoyZYlExry4feen3Z9M1o9dvNBG/7HiBnqCngIH0HrEAzt2h1ZJJXpEnvXJJ85nAdvp
3SmG8ERnqw5ZWvPtO8dWUwiHbDrZoZ2pwFc1cB77c54BpagGltp3D3WTH9mrAw34NOKgBLhhfTMS
MgIZjYbDeZ8aJouzmCMreHxeKRxgnFwvlKQGJb05RB0TbmAJMxhygzjraAG9+bvhAC5XYu/UB4+/
8JkEdwAHXmZkInEJ9L0w+/WQkVg27D85cYyA8ipHYf9ECOD2Jlj1Luw8AIDAkpmHITQVPXEj36vx
zGWgiCoCNHahjugZwcc9+qKoMqvJM6b8KFiDkw9zdkDYRVpyusu+jlGCcldLSZpYkwIulqz89jw5
insjtIHQxHoyubnIzQ/+GaAdJA2/sprrTjJbpQ38nQdJ3uwC3Kqmu4Q0+IcRrXYC63Oz/h+JPhRR
slmFf3hLLjFp8h5JWpCuVw80RiOXi0A6Wixl11uEGs0Pf1c7oklxzalNJ+D8fzYNQHLANj6aQ4wi
HnzRuvRttnq8fduoIDxjOXsjCAplt/MptNLWqe2WmE4eonoOYTUQ2UZ/UMemdSpiJmc7mHyqD5cJ
w59R52jUZLzdQwT9JJELys3i55KnQpHwelkfHixZi9MFu+X93L1RreMC/82hzvHl+n+OF2SpATyq
xUJx1Lof2hWSjFyDvSntA+zhxFu0FxqbvSzZ+ATv5oB3vxAWzDXiKJxRBrr2cs1KIK0vOOHPBQ/9
Qg+RtAyEyxBsuCUjp6ejqyARdLiRo6jhBGog4+7koEx81DUl99PLPb7GEPotuBJ1lSYxqHYxYU8Q
ONh5nDet5rIBlyeVy5O2gZ05SdMb61VNqRGTsEasvXl1tHbS4tX6v5FB5eIPhHb3SWXTilmeiPh7
Mtg2KvujF+KxPal9ID2nwZtZOPEFoOSQWrytuMqhYPcneZrrqcbgCeLhIdGoEAljKCkYmaBp3ze/
PSYp/gMKe98vjOGUEEnohAJ/aqskJxnjkzQCfSaDMhmnbKTxUTzRwJCJg8oyXkr/qem0+GufK2MS
TMdNAM7qPA7lpA2F8/yVLGHUDd+yzgq7LLw7JglMitBGWil7SuJ5Mpoli2I6ZF4fayytOscA0ktE
WDGD7aoFwFI6XPO4uU+k8btgb1FWfdswyXYs97goKyczXWW1WbS+Lj9Xqccz2i/z0CwF8gzuX+la
uLSLPMjDo49BurBzwq9KOCxf7iegovfSNZoRfMHTz5rfjcCyERBXA7fHfm9i7GEaDiL5pouFzQdK
do5JxC3CGstHFT2rKNMlvhCVqTM5ExnWxgk1gxLTtKhyaic8qgGTfT0+cXycvAJDFvD94QoQ6MSg
OhZhqur1xMkhu5ENTy/6Jmoo0qlUXy+01owCwxXx0Y5pynWbN9WCjm4rTAiOE/uZJIf9XO1QHsGk
DOAAFtR7mRfdojISKortGHk4YP5HA3gJqCaZggvY1R28+0wiwpZbnxr13ysvjOujrZyHh0ZzP6ax
0gZDgjKu2QXtufqBvCuTjo0VEeGh0e/erSEu9KUpgnbQUtoaG3M9NMcXdBjuEIQqu6W+hjAJ6Fqe
fBE2MXmCJr+taCKXWSLdMaeyeiXqDPG4AMejpQlcjBjkTNFDWQY5354Fg8+QuBm2WN+e2kviVhLR
vTSOwjEch5QG2khu20LoyYjsd2B1C/wMEZFD1eTDBXqHu7yLN6vjNf02jkuVZ6TmEKHxccqb0fR9
YnjVrCXl9zbmSo7gPW5/g/THiyYIIkWsp3/Bwq4YQnIUydt9z0o4S4YlvLSxPa8uRBgw27b6lknO
VGBRGxsSLqtmEtz/eFxUvgN2i5LVsP/rWvDgM/gp/84eTNWOe0Ahvejz1S/tazhjRz9oIH+j9a6y
Nb2ptPcttawU0ZpvB6NxQ8AZMHEKiYIgTIOpqUJ/5iKxBDJrQQGKcURCuONBOh8kSthKn2p0CAPD
WAgaGuIjcv5+ACdy8WSl+SBN3u/AdFSIoAUahKYQK9bo2Y2ohks5N7vaBEqVggqc2zOUmF8npvYT
xvHpT/5Am0YfQ1eciOYOztzqB4L3iqHvugBlvp5JiYuutz6eXydg68NHh6bFGkjoGkwmf90g/DIp
z4dh71CaQl37X31r2+TOqamEa6DmZrzDGYL1XTsBou5d3/FcN7OrNN7v2h00bNRJTZKnMRtFD64t
+OuSaayAEYyq72qbOhiTqRoP5KhiN1mmzkiG+w2k0rJmAMqdHGY2z7cmHGIP/pSnPfRypLA8j1V7
WpvCV+itbvtVRz8M9XprQMscc17J3v9YJj38HYipAGAS6VPykACHuWba/DVxxIkDD6cG9Ow84VFC
MjcKJDDZeSnwPV7xjdhmFlFvQkjAkNJYZrcbrmd8haZ1XKBhZievECVabQ6XXBfrCsoNKrkK3ln1
ONUypl03k0ZvhRgsGdChIQjLVx2/oa7r5wmbXfYxrI7M9ep1LjjWuTZPS7ah2dr5kZFMG5A9y+AK
yi2M74OtWFi9l9bUTnzHhX0TEuMiKB+bW/1GrCHXTnQispUuNz96gvj6WsAqHP4Z/7MfY8aRSCtB
biEpJhugeK+F6eWxUgBQNjq8L4ZvbZOAWTQVENYBwOTaVaV48DF74wNOumOu17Y1DyW/mz7r3/Zf
9WGY5zKFXhKusGKrWfEdwA36pVWY+4cKuzo0Xi0jbNUoK/w2P4IJ6wyblzOjAhWR6ul5ajq2YaYK
XazgDQt/mQnBGVRgkkTWh2EW6buH3xe5MvzkSXQ8cP/q661QT4qCkN6OyRUeNO+OVp5AOlnvxKKn
IbFnLuVEBFL6rVAOKiRnDydOU1OlCaCLp7g9P+CzlBFTMfwbnkqImvVjYcm9+YqOAS7kwqHeXwnE
MkOpbKs9L3M/OW2DMD9bvti0XvVkdvlx6h9E2zEE1rd8d+3kUxVoOMDaIaAZmXXldtj842Q+F9eN
5XWsiG7+59RlnXb42zIAP/5owc9gz3QhaFDgLtGd4CQJeRzFFNZdUR8AgbxRjRqO5DMOhQOaafqu
OWGtRq6GU47KvfhRZL9+EXcQtP7vdXPfrvlH88UXSii4bYc+JsWe0Pe8jiH7Q1hwAq9tdiVLzXqj
znUXMnMhWq7NB8B9W1W3VDFL7x/0wQmnwI3tZe/MM4l7PPnJQp40b0xOYTonKjopM+BI41sfp2Mk
gHDkCzAk91JzptlgiU8ZkvIJOBMgBPHKntPgdSWibqJWGfYsO+Gl6I5ELpS0qlpUK6FzJfC/C0Ff
e9Sizu6dvioOWu93kJkbM7ZNnbF7iAgRDbX8+VB6TMcQknUMxW8F6ATQk8AYd1BXQfNcgpzXlBCa
/dj/764/IPGFJTmY8zjxVKZ6RvmvNVSxpgLvxoP//fsEI4R3e+wKlfrMurKh4OflKY0a45+SSeIC
yZPYnkmnrFl+DQo39CQCvrL/p1GLJTkQemG7KYTufiRbILKELnAmK0SQ5BUQo2rkMGkWavsptQlh
kD0Hj62MoOdM9snnp8WBGOhGTN46GW2hU8k+LK/H1l+9xpEsrhEoWI/sqxSoXhK8z3jyTxulRLUH
rfsGt6fZBd82qZA0KlF8gpWqyXh2MSh8n5K6yWIhSKLrBZ/Fw8jaei6jfgZqZ0fWv+HPnlpTHRn2
5o7klhcZKzowDHsA2oz14pX7iULvati6QPM30FNjFjmpXnuZ7JJFBm/cUcBm/PwC0VdpDPO8Dkpp
kOyCx7rKhNbYGKlYqiXdv/OFN8MT5CYrtEJd5f+qkLZ7vOe/rClHZsTB7PvThTx6CvU6NaK7LEFJ
WLldvqFWSVe0ZuVCnPooblv7o912iYe0s9xVXGcUOWWfqsMktrhXCJBlOTD2exSurmaSVrNxzDzZ
hFwP5Y5DIPvauXbk85xpzSs+DTX34CW0vXrrMJ4/IrEMDQM3AvRm9ADd4ElvgvZMRgR96s3bL3ox
S4OA6vVptoIDvD84TbH5PjVD6p9acx3CWyz2k8SNx6Mzl6PXtxebhrZtDIc+flp6g2zQ3VTPcilh
q2IafLkXT941M2ejnzTNrK6VN4bNYHnbxTR99DFblYdEVwlt7DsPPj4X17nlYszLKz7glMLgEIGl
blq1btVKNifsJ0ycLUfDqNyIvinIuqJ4cP9QtBLeEil7B5oeN6l0oJCYX/51gCd0v34JTvUcqqTa
/Bx7HLxgRFfIzxrOLf6X+qot7h4uyOSbpKjqSGHIN5R/3ZZi/gPULLnENWIWUvsmJDZn11QXL6hj
GqxduVTyBGScHNhDwSExwL1PhVeHagXEsad7lX/x0elb5fnbpC/lUj4GYqMF2uwyMJuD5ap1AFGA
gpsepI1oWGiOA4J2X5kRg4xVTpqbcA5GHMVzk9Zf6d5kFqipX94/WQI2mtl09Xmmmo8v9oNgzxxY
8+hj9nqGMd28hcYh1zQWwwfX9J58zSYMIwHtB/FIQFhmu8Qmo2BZnKWBz4icqzn+1S4njkJH0Dyr
HevOPWQWW0GZOs14WrKNFBoQ4Mp044ONShduPs1/YbMgABBzVH0nYE/A+xgJytnficya+lOo6Hjd
VuTraXsANIds4zQYzzlJW2SDD0n7bSFrmByDCjGnFVkZqyTy3knNYtgq6umR1Skj3g0Ho6Z75U+k
z8fsjB6TDIyJVX4Sb44e/7bsWvoaGsXp+hRiXkC5z+6IB9sCIMzG8sJvaasYf6FsNCRG87y3xjn9
eegBRLoYD81GsHQ/a3rS3xjQvnkhewftecHA6ZA3ze9vIlobIOq5Bxs/HEi/dwQUqTeWNS44/7FR
xdGhUw4k5q0WZ8CylZSHxBFxpflNVhfJd2OoGUxkHOb8pCEc2XeU3sbZ5zi7lIIqoFHvQPJJcUC3
oo+TRk1LV/3Oq2E5pW5WeSsdFOmJgDm2bUPTwYpVDQLmcXkgmIGcfa1MpfqP8ED5/0Y3RC1Q/FPw
uH5c24SFwL4YGdXO2ILbyea59Fhzcsy//1BtdBoNyNkNd2zmgeb+E2QSOcxBB1n75Sl9fyMCbc1S
6whqtDnXmiDTFFQbvJ07UajZ3x+mCsi5GJEiOGNbMrkawl4fLmqO+1sqXMfbDWlDFDMsKr/FpXib
fpdSHDvHZ3sbJbXObA55GH/Ypj3aoLOVJ4CRSLtRdHNCoG48gwWFyJgW1x2oP8aTAU5LYos5nlhk
Q8i+CdijN49vQhFbkPiEINUiJKmjvivTIUht7Ps6yazF21qjmFuWP5WvgrOQSwVCEUd/Ew8IgzY9
7QZfYIHneh4lKVOVHr2Yin68GHgXddCsOAq5+WkvoMvFtNZujTEch8XIO6doS13LrBU7erGhsNlH
qmKnTBSFBpY5GRfrUHRDGmZjcW3gRNnF64py7FuJp/brH0MVMB9C0VdyxNeMqxicTwVmsaqSQoqh
3EtwGo3XZZ6iSJSsYSUAOg9uW97UR+LqWE3/xQddBVGfcb1BpC8hU6WPs4zc9wDEV8m9SO1xpN1s
HX0N6qx/r6v7H5PpQGnkSggtOx6WgXbCGQFHiUQ07M07LmFarX+TvqVfbQWYK0FNYhPKuYHXcA2G
URnefyCjDPX+jZ8qkFdRwbW7fyiS4SeFwj6K+PChYIiAAU7PjjKcD+wt2YZ+koWxAnTVBm3KDEsl
xrKRVfjNPZVtnXxRN8bM52ZMU257YoQx7rXCnq1W7hjA3BYuL96rwpw31yT4AIxD2gZN0PpseW+t
W5kuMmcLeASnYbMK3Kw6W2tQc4Q0edH7f8AEQFNM4zg2IGAFbOho9GPwT/I6d95oJgqOJTjSy4ub
dgT5ZNyH9P5SNKOxmEi83GYttqyBjmctzgbsObpgJ9Sm9v7w4c/f1FhEoXZUaWoNp+m+1yFwF4ic
bzG0/EISPzsEJDM7WOPE2nBrXjRMMjmKENuQGPWkKRlHKL5tGANyBPh9OPwYsFRwTpetw5k9s3TQ
yUdhVfrr/JSTWbI8qzZXVcewS9ynvdCHwhxO14U1V/2IZUpxQB54Gdax5bCUyfqsmRzCbWgmEpFy
im2Kg9oEFZynHpkTz7kD/WjLL5zQfd+N3MWf3dwTsuSNz2cQHiGVmEQ/qJJ8pBex0R9SZTSkcG0H
We1gQ1Vro95/8Yf+YBMlGdqwCmYwbkDxQlRXIArAtybaITzEqIHzaOSid8uGg1N1elIfsCMMoJ6G
Bxo5VrAQI2ey5fbReUmyJVJ65quHtKnwS8y+N/WArUaUpia60ERrDLW/732mzY2bqLCb0VCeH04i
PUHB/14IiW/7bBiZ/1XxBT/karwRfVYwlkYgNGIHEl3dm1cEvc77u5QAUYisF7Yq34OxMwlWrwtV
gjhr35hL5GEVRPzkvNdAwn1CkzZa+hEvEH+BNuu8eXKX4PEwVWxosRewHinOtRmDERDoSYCFxjUy
IsKTNniQXnfKvhKLdHHlOSsolO0H8bbdG1dnY+2o5Oh8NNKBbIvsL7nSYveVIZ1S+NqAOCN1UULF
VwPjHl9OAFQEDV/67DybVPvcRdmOakaqn3sZ2x4MY7jVgd8hMvOhRl0w0YJR2NROgB9jgPTBajjQ
s/0rmXn7TbR2gnpUJzKcE2klbucaqX93sktdsQYRy0FCnlV72NIuOI72iH17OXrl2O/8joc35I4b
nXJzyPivduA0f3+EzuT80/evAAiL4rJxoW85mZS7ypGGL+ITcDZjTN+hDHjItcQ24hCh6MAmYGgv
f3Q3NXFYxp+/w9jgBSv/m84eS+aJFAFwbeQiv7fUV5BmDa/omjH/QbRXuTm6HpiE5Lc8UzyEavmC
m5UGtGsaBY5XppGFnWQ2V0Jm8mBqAq3/pXsQhaID172ClW7yT++mLLEXyj4/Q6oie4YIURAJuC3g
ep1aBrjcgXyKa/R0j/XFxQC2ltxdEpYI+iO/z/uKjQNicTIm4I+4lAfa6ErUVeoLJR7mr6vKRjAS
qVZuuCQhMuGtJ34AI4EwKWf9B+AbHnvqvSUOhsQONU+WvDY+FXVjy8mZ6cVg78edJBW6SiCSPGqE
Y4LzPl6DrszIB9780EnQkTHrwPtaArSYhO75iw8nQGiYXaYJZUm8BWz9yFXm+/4HOHWsN+lOu4oI
bpQUYKdr6WJHY2WCTJbJOcMjeRJEjjHaqi/Slc8ldLf59Y027SI45/dDNfa+JAh2UkXPaf173N7t
U8e1yy5BdoUIzq5vu1fWqh4u9qYIp2Ep1UbhTuBFaG4460jsTdktGzCyaV+RmZWSBakICYsuaTly
M5huPZxJm1QZkWMOIYe9wR5ACKEEidkiphx/Zaz07oZO/DsaV7B5x0WbJpeZRXizyrIaWJDvsvq4
bzFS7Sm3bpOaiM/UYNaOhfTstbEHM7JymKbkKShvERYIg4ZE7dVT6XhJi+2wSPcpGFcO6E7UCaZi
5uaDSGA3ZarqHyJVRbTLJVClui87M/YSSup4aqZO4HSqr2CqmWkne4GlZGQAZEJU/ojXh7pRaknm
ZwEkcmq7OG3h0zm6uDUH7YomH9mJyxmyjPotjUeFRayaTXm6Wj4qTfg5IRygSW5gzcAMSquOO7pF
BEIROlKiBS9UwbPt3Puu75ph2lobXhHiJGCt27rQaAfvLUgNXEh/W1GMrraVwxQUNbockxUd21qF
PNdqATQCzXLoTMd2DrWvIE4SU1TQq2VzgDO6UIwz6bsJaAie4fqFP+3trcgE46S/zynFwdKqsQm1
MvB2HOUX6PS97MzV4nO9Qcg0xcA8sZdY0FH0FezGBY5rc7PFG36+ZU/MduyYj2qOpOln63tiAzjb
/nJaJdeeMfezDg53vF1hdPO2uyUazBp/3JMipacIBbTL/1t9fATP0T5RyK6IsXGIze9cNbPmf6WF
OYeP0rCuMekIBnwbvQSuoQ5U1FHoZR+8Rp/Mx7auqGxFNOTbR+otFSehMxBrPQbJSSBUI9AnVDKY
AmPqxk/OdUBz6NYE/WKhwHjTZ4pL+PvUyH13PiSWByvN5vR2+k1669eZSDIZTsxPyWNMRWJFq/c2
70cUe0UaB4lGYYUfmH6MZNpza22sNwzrVgnGixdjQTstyGJo5fVMR2edBbUKsbbqPefUmcN/rYTu
vYuNs161Bkv3eI3MSpfajtF2L+DotXd/fkfC4YwgMvNt/RflpSRjDYlNxI2LHHShO0phCeLy1f3/
Qff5GRthKCvMM1XCi0jkq8+JDli+zCs2GPX/nFt2fqApjKRp12SJPqaEpfSYqrvlscngNsb/6rrf
rYqwh0G0oQgOwdD9B9TLwGZZrgtgNYDBH+WW46WRP1U7Ef2il6Vd4hIRbkYnqgKP+p2UJOfVry6K
4QclegVES/KfFhte1kCeN2bPnh54uOP0AzKiguVMSqP7UrdVxQRMKx14KLuePew+4QyGEc8dJxEm
DKeowtAp6A7HeTLyvDT82rCcq8UhdD3w+4KCOi0Hah+KHp7hWBCZflnORet+jWvkpzjGkgL3Vjv+
brUmjjmJbmWYZhwhGTjGN5nbrt/AEQtdaxp9hHLhURohfm5pX24Vo8x010Lg0Xk8AmJ6Kifoi7SU
iL2+JbZ4FI1KMQ+9V2wleMPhp6kC0bKYHdr23BCI+UHtx6N9rHKkHAB1J7mIQNcS6c7bPYNsLwwS
KZatBixN7TisM+bazI/J3Nx+UW87sBuwEtaWljaAoUSPdi1AnNKvEax5fWH93tXBd8fFSwfVuRgt
Vu4cG1F15iMZmp2XLBYVW+XI5o3OW24xh4aKr/03P0gLjEw2aLxzQKOLMmrIGO4U4m2Y5krw9AeD
+cdE/a0/adCOb5k1PPF3RcuNiZ/v+1fG8bxYG5iH6yGkxBJzxxuTnAKRAc/Tvl0SAMadnxMqvlAW
Vf1CNHd3HTroUaPIKNSqWtjrJ8ZISUC2E5hWdFjx4Jn9e2edCzEESyAraOWf/OkySqc58DQ/JkCc
wUebfqEs1eko8cH9+bKJR5ZFjaNpRbqxHYYXiEIMo6091qa2YdN13nJEhjsi6xULNXL+feQl8vf2
ZwbkmMZMcKwsM4qJCTZLBzzvb6IBRxZCFX00PvWi4c268RIMSrUwLPlthNLaFB92noiS9LGq18FT
RgiUPjDk/aue0Rl5m0HdFY5RS8YP+8VrIfc5jzDT1VVVCvNdloek8ru/iw2KHZ5phnlJfwUcjRCo
1+qQ3Lq2P9HEfRw+eCueIYN3tovCLM6wcLxCbGuvklkCqbcA3L+b7Pya1jnwZXNN5JMECYL5Y9t9
7X0EBkIOgmuvDzZyglj61Fa7r+TiiEwRK7zJTmkd76ksVdpsCX/sf0uA88BmqaOp/7EeLg6PHnTP
nNbHyC+tORpNOSCgBNcrtxzIvzgswCeiIcWUOjLyjLeV1bqKau5zuSDiYedeVZ3g52UQyeTRga2F
ZvtPe8fXh3R+XrGR3q11fLLAxgTKTPQnCRUhXB/0ZXMD0ExuDMd24qg5dllKgpwoT/sGS0qbyirS
Wnp9Wr7d4N4Wxi0hPwDFcuF6lN5H1nvQjLycFJhnUntxr3mm8+7mTaAECp0iBqRwJ59DFc8UGxB0
tfvyCDoX7++OsgrguOT/j8L3T5oMJ2Z00Q2V1SgFkLId4QauQy1rXqObuVOl+gkZR/KISJZKH7zN
yxIKUjQmlovBXDIUE9tljmg+4W+6DfnVOOZDusCW+p9BIxD03K2eG6r81SNge3cSPLf/ZH4/aVwg
pLOaZod5EDH9m0Lm1ysvaqRLr1yEQSHy+WHtSIttt8rX58C6qNF9bBup/XWMe3iF1HbgT1zuzdKc
7kbRQZ12sGBAjuvzN/iKiM/9IL5pwkZd7xPD6AdgKpWPlRbUXAaBypU+VY5BIvbxtWuAghXjWLC2
xVpkU3O6waR67QszYNxx5xTKgOWWOtcoX/NZF7RCtLWW3hmy3zYNHaD/aB3nIZs/jmDV9LJv7jCZ
fHI9yxXf4kV7znAvtuByRe38uHG+4ytHWSmIxsySH+ukz/fMTLEjV3qJUnpUbZzPv0+CvIum/dkz
L4raIEKS9tZ2Z+B6hyoy+o6KyQqyBxtMq+LlfQ1NQnjg1TC0mbyOPZgQf5al7Vnf0S80NmbaNv6W
MxJq8JGN3jwl/IGBaZKLWnO3A3TSE8PMueCCD/jvQV9bCiXKG/kAKqQqiSK4G9srj8oh6TtTTs1+
nFb7U3dVz/oLdRuN2mqiyq6tTl0xRtt+gQ0JdsYG95GJvIaj64BPP0F4chtG4gstVCFvn1HHcn/c
L7tvyaRciqtbCgu/+PLnwa/OClAxFfRcFimY7rhQUI0ajkluI8BNcUoVCWME8aa+J9tN1vIE7405
LqnKhnXp9fzK9+Zoun3btFXjEWtkI73xNY9WvOFFS9wIWQDUJG89QY+K4zddM15r2E1klSYOrres
3sQyQwm9Vr6IteUuWPperdEPiJihZKskORCNNziJH9oLvGJerPV0PURouS/g9pxOuaOTtx8Kp0p5
KYEmMeN6z2+33O9S6VzAWpWw76yxJFN9ldn0YNpsFDr9rBzXD2MvZphuewFcOjkXQhhIdQK4Nlyo
FGmvXD/gbANjbZ/M7jRgHBr1DlGg1V2B+QreVtLHHOYNurgy+CjQVcKWm4P/IaJR1qXi61QKorHf
BaWPhVKg74i2yCp4Kut0lnS4u8/rZswq/cr0TXhHA0E1CSRrvQpInSFfD7fzzxmCqjiOX4qEze0t
hA4rpl9p8tat4++u6DuKK/5bR1tPiiPEjZVzhpgVsB2Fw/YhMVuv+Jux7LzNEpXdxZCk/7U0oghW
J5+SnzXsc6wHoQDe9ZY52ZLaYSKBWMwNq3uJbK5lJTDBKwWPpy5hOji2NBazOdkVkZ+CdjdzwE8z
thdJ+oDW3cd8h+96MU4d6yK371EJF57ZLu+QSn8M7qzht7gmxmLqYaZIMmRTer6CBcpkAWP3kTuA
c1yZe22gutUVrpQkeunHwR2/HevrZv4nMRJoe7RRvoO7zUCxOLvT6tKjrC3HsIFdteRmTvSaMyiJ
EJDQhXVhKUqlDU6YZ8VYLckSiYwzT0jyKX5J23MQNQnzxSrRucJAC2RoDJUipgluJq1XI+U/QTAW
flSxQ2Wh2vxFIXLeWNM6gzlxJ0alk5IZtIhw+C2qh4wL4TH4yWdH5agVI3mKiZxLabILQWLIarGv
vTIjRo7oMBB2fx58MxLw8f9LHFT19EeVELOATHoX+PUTrKN9Vq6SFGR0Wv0ARdNUK6dDWypFuoPU
8XQ5QO54cFjyfwDjUl2qC4Soosa09ocxqCacD/3W+r0Uryr25aGCoBZcdvvzi+uYlaqAewIqnqre
e6LMPVYmdHJ3sMvmSFnwASv5IMtWWkWyq8RSp6pNm1DW+nxPFqHb3+wDQ9qvTS1NXBjmQVnt9DUD
mjtS8aj6rRwY05u33mjHyutMFvUSEyUWAuYRvQL/Lq5LI14nBYGhwLfoCTi2CZNRKsGEbzEA58mW
eLBWsienHlv4+NMeNNoDCxaiXSF5Unj2qZq/wKKEpjs/8xmr2nUb5CjQzF2+PdVR6uhi7iWyvFAO
wwsKLlOjXGGbfpnMILdtzjNcAqcLRuMqk2K0tYqkfg7Gw7sG0Ig2hc2aLM2FbsrWBYTv/0qFXSWf
An6xAo6OvwYxpFaR9RLSUQj+PUkECNjTtZhowbfzzveG76eF6OUapu+UftkfA6Ubaw9GjBTA7o67
nEuEgsNRkykf1wBRYU/OgDk6V7CSbwIRDLCSlnDfVgSgTBsnsaDWGF+6kmQdlHCgJmfJazSQWRmG
0dblM6VTV9lkNE7fAHrsBm+cHxbeIQ5l9QTPhpqhLPzI4cqM8aBxtMWiLocTvIDLadlj+1FJ9DsP
Fax0V99K8zpxVFdI+U6jYnDgOwIDxaJmWWZzS2+G/rt17XaxLv6WpYhGeERzmyIqQKdhi3EvtmgK
6Y1aU+OJAmNommHpmPdNqEaIDia5htbeWjNwN7csPnrTi5fbvjwhPvplSquukif2UQhhkKNd9Y7M
fwfFWG+lCnNmvS6J/oYW5/ZMqzGRsHhFzOtZftoU10URcLCVNXgB644hXe4suAAUqP2W2W2kEywS
0uG3cRxsmwuaJTrrwt7slNQsXzHWm7KnmT3YAsAn3SpfZLvWEDGxvgbc/FI4sGM2FqouYWfNIKNw
3Y6D5GhAuPQDvuLVM6XIxOYvmDX8Rfh5UimyxOx37ZB8rw1lw354htIUQT9uzDMpsfp6SRVpe+M6
ZJvis+GGRHy+F34Guq0Nh6uK8K8Mvf13+buZuVh4zEfkXaRpwuA4QcVio9TUW0iWon5vtOhUlFM2
kP8pMClBEMDzgJnQxLqu/gM+Sg1QPXaNJIxNAwHCDj8KTQlYluLYnzJUCj4xajXd7nGSvyArbbqj
gllDFqxE925W+UCvNw4gCFntPYMlo0tG7t7pipWM4mhaARP3hoYTO8+yA0gavj/E4gZA4ILAHhxP
6Tku+8GXqOI7v/mt9qlx87N7QeWbrdXNsGJBy8byU2pZZDMtnCSy7xl6i/8BEypxw3FydP7X+Ak3
oN4Y1zFm7ymokMlDnc6nP+iVm7zqaOKPd54KADmx23mMAo2pl720f89Fj3A7kDpepb/8egztRoT+
LsSay3NfUtcStD/qEWTNmrij9vX2L5l1SZ4ZII3SLqv99BfOiYrcpzuEx+IVU/rHsvfM9sUr5srq
W1lmfjHol94CohKcWxIVGcCGY/L4gVDZVoA5wFAao+NdD/sp6WdOaZD6SQNCg87QJKpF16orNxZh
bmFN6A1Q4KldWX4JgkFY1wPRD+eg1hRDjWOqeNe+YsaUuvd9CL+xGHGusYYoNu24CgVRtv91n1Yg
4hKldjdiIQEYu3MyrSTgpuF9fmYW4a6RHuzGSrqNEvsK+TEhlhvmygNERra3Zkf0xlUmwaIIL1hb
DrnJk8nXM1h5gXwC1d6D/olykBJC+8uImWDwTO7iARnjOhroNMMUFJjn7eELF3QcjLRPUlB8RhW+
iPU2Diegca5RRTYAtLV3yMruGYT96HG12CFW9Gso8ebB3D+LgCwXJqAqKQvvtNcLRwB64xhCeAT/
mduVqTMMEyw8CCLjalOXAxe4ISeI3RB6bb7M9SEqJcbRmWIfWQeNWGRVSMBFvDXsAcTjOgurvrS7
OXnbLOcVgW9DJRfFE1zyh/V/Cho8peyNoKcBEEVU8bLa1IfTTTOZ+kG+uUY/OpO74npU2fv9VHtw
qWDhNAlz87MD4LA4m/HsNfEsmAwPfl/sMXfCVv7GM/4Lsa18mokM+8Whli0qzkK08Sp2YYkcPQnN
itYEJSa8W4vEX7reXKgj4OdVOgYGF2j8SRmNfPzGnN9kPzDQsnsT46lPGg+JHzWyW4HP1QLQtU0s
NHctjXRpwL++NpJyvZqXQVBcXsklZyJ5eUAc6igTLacWHuIGGoMyTmJBHoxa0fVq+Vcfn0jUcon5
U1LY2DKwhaNExm+yKaOb4z7qDJCmaBv2HJyazKFuQdxb5BxhaEGSNhNyTjp7uxe806eQ5z+a6clK
unnf37CClFOUZiP32XNgJSasUkBaNVwQNZB6Tkiu+llukpQJT6eSptsJ/Mqa1WJBO/JSRYMXwfD0
orkvXMFrvI4igKNg+xEPimctvSQ2jb52KAnez6rAeWSnjGzlh7WNuwKfER/Sy/NqaBSoVtWHzZfU
9dMUnbSv75WNBGicJA1iBkBAssuKU1u3Ze/a8+PuuGkObLf0WHknVepMMD9UO5mE7Q91k/z0dees
ysmH6FLaRFmyQjOFi7T10TwNQIX7UHMG6eLzamw6AF4BhIWqDCX9GehPAwAT1YOh5PpefbRh1F19
RKymh+hKBuZyxc0yBAlYiK54ul2inf2xBN7WL8fWCjkeyxz/sJqienO9Y2+sjD2UXqq6dngw90nK
Mqjmojzce7y8EcK296QVJM6b8VTkQa0KBDvNrApi2UL/1mQ6YxCVGhCquz6vuFuEKeIMvqBURYju
7Hr6z39vQwsVAXFHH/82UU5uBD5GMAcW3ZEvOwMOJaIK6SIXpipE15AZ4wmSqZtoLM2ZMikDu0LA
Bp//ywd1rOxya2xV89KrFZqy24RmODB+SL6fl6PH4ZUJ8p/ecbna90NuvWfmNVudpFlC6R3Sbq/r
QMlR5ZLR86ZetMFx9ItzM8h6pjKUVDNOa62FOYhm+w1IHwahjPz9S8RLowShm0nYgfE4Xgs8sMJI
4y8ycHiZKyIMo6ux/TodRWEergztDp1PdaZ4W4IXHunO29etH1TsKppKbPHjRziMRM1+fG68gnz7
oe8nGXfV10i08ihRcWyQyD+kpD+9/JPXzm1z6Xr/hEVxbGa23QdTYKh0vDCcyfNsjEJEBfjHngca
hHQjiyTk22Nrr+10aWKICPuKicQeEeERpg05hgJuTrSRFO6g7JLHoTiOTKE+HrN+wTNXlv1skzf3
pMaLHqOECj94YJ8+pmMAKLTkWXBbLp/8NLrSwyNy4DJ1ObbisTS9bv8w32ZkaaOp9gyDv3aQLHr1
gS4zLOavhqreMea492Bfu84F6PbEgZ88smbI5UPbKmXkHO8ZL439qdR4HIREjdygQjnxmD9tvtqm
a+QlDqjtr0/26spYbSMkJx1FvLYaIsA5kBHt6Vi0A77PCTIPNpKYvP9nZAVns+gLSS9/E+Z6IsEQ
pfF1La783CotY+6IzvhiF3Roa5nKfYUZWlTiK6Rrtx7665D2P7enG3/XoP+nYROwxR3tmf8VcNYr
P5IqVBrMh20MLED6gomBR6rS7DX33nvjTzzpn50+vz2X5RrHuJr27z90q3pjs+5IXTI8bNWmCUzW
pGVTTA1U+6sQLYMdmCpgeb2ESPHhEDLxYZQUuzxkCSGTrwpQSrn7R7LNPTOJE6kxfREHFR/LW3YZ
TiYKJWzIJu8xlxqzkEAL28eDHQDW1vAIg5m2+K0cDMRpt0k5z1wuYaI9ocMfMxMwCRFjGRAuoTOi
aM0mT4TWOOjk+RNcu9PJlZr/Yp+HtjJ5FXaxkIvjTS3ir+cAvIq6sVqZO6czOvtQz39wJ8IJ5Dx2
Ev+alVO8X8sfQNZsFQRPUMfAG0Rs3T4PD38xjpduTMluDUGp/uomAhH8978wEr/jhju21xSVoqfv
nr0JD9Yg5xDGEL8VSahXPTkdmNyZJ4iMbw3FY/c4UJ1k7a57JRoLDuDwAJwGZRK4Hx7F3KLWS5JH
U0y8ekC1xAkBGOri/pJHtsgyP1Kgr3oChl6iAi+GNL7mcKr88Vz3u8mILQW82fWVkadiMFbh5vL1
l20nUt3VOyBtCvetsGVVR35Niwk1VyPkrf1DHIw8ztyUIVaMKhGKPgTJ+XPtwg1XzUzRHWdaXhqF
7UnGYVlTWGSLEs9D3T+CPL4vBDRjix0QvO7V7f1+N60NpwDOdKbjTIQIxZDLun7Ukp9yGYqFQZby
tePMcqoXTTI96BTcuTyve5Gz38hbYBpQ1hlNNpEDI/ytROkiqyuvvd0ERssEIKJEFnQ8BcluBGLW
LWzazcIKXsXSM7D7xzKFzFCpqmswvzxVhrNhws/gyUZUknYtjYF0iRYN71CfHcQ3FNJSMGEGReDl
13tbcbm1uCbv7tsV3UD7OR8GjLTmE7hcqctNINMa5XzqaPlsrJbimeupASHG0LSHeEgzCCR9ymlh
B81/XRzXLtfn7aOa7A/lS5tWZ6FqcV+hx/YATwYU6UThS/1NbFMuJxW0uAX+NE8g3ti8LUtRvgL+
lzfxsA8vPKui4eFGECj35SohMwcxItAIpUEzwbTaNZCrGcoxl1ibmsa3kpg3zNMsKfiUeA7WHtiR
qQzdiPxgXDJkBn1Fs2/GSXEcvw/dFeVofYR/boCHc/Y7Wgtg3JdFsU2LoWqvBmWUsTTLP+edvCbF
HF3TNzXrel669toE98HXTsit/OuhifWN+nmzR61S6luMUIU+/bjbWolFkKaqVFfPSGT6Hs2MuG3p
DOu/2aCuNZrm9jGMA1Gx8trrOrrP7UPKVFRWw6ZKPUmuZdKUio10A6Cf+uHspao6FmEXgRF+1wgH
FRJrYQLir16+13Fia/ruA06LuRZiQDyv2+HNLSNyGWShzdKAtMHgQb+f5aUg7U2d58t/4926uIaP
OJCP9eX3ihS2j/+9cFLxEKyR8UicXG+3aTxS1Ptox+fSX7W/lK+M14ETWUzNwtoEEKWKHcEqtCyO
HnAz0Tfb2tzik26YQg5mN2SjQwxm802q+fkqCLkTpWjDrFagPyh5ZPBLRVR94QGo5o36kjNpvYQU
6Ch+Gr8bRvxTh137ugmrITJ2Yk2cOFq96rE7I92yFJd8mhbIf87Ev6a6qF/y0Bbs1WHtGfNO95Xu
i6KGAxR6KZrjREAXybEcpJdpqeUq22Agr5TrAZRlr4ZO6tF0a6FnWDCIeMZnIZYnHhnwvJ51i3t7
Vx8X2KB91Fvt017UuPLpVCXlBblK3NgIy9/xg4q7u17weCYM3zcaaWfSG4JZIQ9uACMJcpmkmgJZ
ZBYqOGpbMF4vKQ2XmXT6/Jg/0u89pZgTGHDbCyXX1odAoRQqqYhR1Apq+N2t+LGL2S96cvQXUdkw
LXNEs75hg162F993reXfdwgEJyfKRxJzsJoxzQWIfpEPA+qlpntBBttAG5WOf7kbOjOHM+RntU+L
qjdmxdbmmWIeyZ6TugyNVON7jMaZD915CJz6SRtJ+T0w6nHzmeEPc41uzFVVU58+trVtTlryqkhy
AfUwucMITZ+xVhJFreZOl2de1LO/7fcEdkPh7BfCJRW0O54DolZLsi4ieMrlVMxAllitY5nKz8iW
Jad5nBNCyNIzhGmiDAQJxL3685ziaU2H2cDJhfd3rJdVS/lBinNIfRas+aSS4H0+MO43Wqcrb09C
tTcqS9EcU5tgDQVQAwsTs8t/LhihxE+Evd2lu94hHJ789YFOZ93HqPdVN6UVmQ1ZJ6VW9ieVSmKL
/xX3Rz3zOfM93+Dy+gQhJTVu91Dujc+k9xvm8eevZubijw8hEl4HxEd5Of8dJDo0bl39/PTdvYEX
lbL8Jkh/npDY29849a3REPaKuLq0vA7GjEKjpfIPCI9ur5OS+uH8zzh1rnIf+AduhmpY21fBdn1y
GbVZgzvCKg2sj4blAb90jRQP8OoFh2e5zPFtgciQkciL1WT86Iu24ZrHPsfliXopLc04L6b7Oaem
xf9RtSJqeGt7j5AyCA3zNdwzdwZO1pBqDXYoMB9FeDMR1tFpQLt2D0UvBITxPnFJ4SZsQ1DXpoJi
g8NwZTsE3bcoC41mDRcQjvcf+f7OxF0JN/u3sQpeWNiyNZAZKnxHm4psSZ11rfVgsn6B/zQ3IO5b
czOTa8I3P09yLUtwmRx5AFHiIr26hSAXcG9V9hDcSMHWKXSmaeFRL8iGddW7HZsZAKbncSh1hZrn
1RFWV1DnFjwm7KNx6GvRhrqEchrg1uSqygoVg2u9K/CTw4/bccmcQcLTVX/tERXoufOap0eFoCcj
VSuACTeLGCkO+gaScetouQMZL7ILhDATlT9tpnlSntfThUIXiOrPZMr2d2bZWf3dfPxoVvxRXKKV
tvMpupzRTH6AdbP4DPz5OVCKN2tWiQPprSxRSov0TtJ9zZC9lT6FmC3qvtE5c2kJbGujFmRklMkw
mY7idUlNGTfQFLAvuq8IY5Okt7+jLzXe3/7BviutTTtDeqa9HhcVpXWutpvTqMQ3XvNLEEAEKTQY
dnARbjKikFWF7FV1aWY1Mpc9uA0o15GnBtzCxqdKZZP4OcDbHXBaiZOQuEy/bRMBdZIRrhqNcxhJ
W7PKq+nfvPGyzWJlRtixpVGQ9nJgVIHr9MXwPSYHXFJC2WvJoWHV4SHsl9D/K24Vo2pCq21XG8p1
I4OQR6cM64PtL90z9ZybWUiYJ7zN/2BGeuXkU6WdHCS9125UFXFkWS+S6aUFUvZv8YY+D9lVWLoC
Vu0xxMsO37Kh6pFK4iw8oZ6xj4uR7XL8MN/VJxyU0G3se7rgjreNZypKoSa2hVMWPUE1LO/SIhTG
6gEJ4smRZapYkrTQHAkuy6H5AVLt7jbHYPu9yrPu/0Y3IO3Uu5jE4VUZSZQe/58b3wzYXyrTBxCI
d/tOMUY3xUqgwkgL1kQ8bKcSowMFgRJWTwzq4V1zciWo3s7mu/nyHnwjcDGW797gJBzHBaekyFZ4
C3DW1pWEUA+aOYifrExNaqOVN2QzlmMjiMNzJEkJN2HuWZGeDzptDMlTcF7faaGd3PyOswWXHZuq
ZlrnIrqW92tN7HaX/fDXiaNxiLkxSktP4oURDlw2REybFmOphcvIiVlVtIthJ23/TnHiYONQFk2A
IIuypMZMYnl0HNZ1rqokr1iC2cwjAXYFtiqAe8+2NjUnLtCDM9M3rtS6uXxORk02D/Ndi3VTGUBK
HUC23vXxs27hAGLxhdCI0V3XhO4+G//TulkCS0xZRabYW+tnoSzB4DxoLiQpDOK/kLhSq/7Bl1Mk
01fdg4QD6GKHjRYfzFdckbcQ8sfRaTrabhIYcev+OtFaNZVEzemyAmYWgX5+3Bc38tKfTeUK3FLP
PSbYLXvplgPIiOdcnacd7X1+A+S+xX4rqnVS96sYNyVj7IdMQ2F8++QySFKw8mqpmEo7uqehzddV
nJBMag3nif8l7w+Uxx580plS/GMp3hiZM2n5sQOuxoUXGR9JzrRxo9fNrNUiNMr0BZCKfjU08JVz
SwUq+nQ7GWn1XM7hhFFzV9QXHDj9VVJq5GRaS143OwoXQrdPCQXa3HM1lmPcm8sq5gBtakA8aPhk
nTmOUylXwmXhx9bUpT4BpvFh571BexFMbJoMBqzdKQkcY32stxWijCsBaBtDMMWLngb4Mbby9/E6
Dh3Je3gT7S61h519KlMP0sLKtN9YiuMmMgC5TUDBntWSlu+c9KlHar3mwzBOvwG3UfLPDN2nENlI
SDvFz47mOJIlnxXoB/070B7ys9g1+XEcJ4FVYbaofMJuK2aMAyVnAnLDboiuA5wbjFQAPgrRBAwb
/Hk7uAMoForRf32T6mIZUV2SF6KsjR9gyn61UYfHC4bDDFX9uFb4tGtaub6T2hTqtjTWDKCWGRR8
aFkE1tQ7lENrZb1x2SBxGn4nmTnzyqo4fP9KuF/nbvpEvwH4xyFUV/iFNxGGnOlaO5kFt95MuK+n
nH1DP9T1Egf3j5vwbGv2oXTcedbe38+IDQhaaeN9LqnesMcx6BuXKXQbLwuTFjdZj2SK9Gm1At4u
pROR1TWLnDFil02hTwIxxvvvpIX3oaGPwtmjmFHhtc2PAtqnBicVtMfib8qHfyz7lri0GU5I1CcK
ul6z+FUXpc/TD5/xcBxe9HpAOX2qeNzntzpAJ+mbbg73WvJi6LRUSKMkLW9PWdHKsmtwaEJWr1ah
xvaLrN73GENHbkgqoCYUrbg3KhHtxMykuBnrIHst3GvUWULfWDFpN+OMEMnhED+BOtfDTyx5bdMe
DseO6PHDF/cp7dO4VD4YbBdWSqZhf5Iu0H2mtE4K5NjzSuTkEhQ8TM/yub42jcGHvM8hw6iWz6Ek
GYMZwKXDf96j1buf7ywNrS8qmW3ROwMtob9MneRX8+5UAcbWORcCUou5U4oToFSCERe6cW497Xqb
VwSF20bIxp9ynFqWAlij5fvT3lHSZp/85PJoEDZ5oPD5xL+dm+1DVYh3I5w2fjusJlgAxf3fhpGu
kUnKOE/gsoI+C4fjdJsvPtg57A1MEeIrAwhVcwKblQ3XpNWwfUQ/q3APvxS5b8gZ4Ui8AwlSJiG2
GC0bwyIe5OJnZw6oLAImIaWi0UgyUwqK+JCxiNGttxVzjOYjCePJpzj3mT+jZgcVGgrfH3YEM3h2
5Z8oD1mmasGwJsD9+TNuprrGvb4goIpoTAqfLzp2JoS/rkTHEcmSo175zH7hMZXmGmpeKK9/Xus5
ODU56Yh2VVeFx9sqXHUyjuINA/54stXFIUxy/RgTWA7bbIHsu/IOUiyxh5puKekmbnUxiaHnGHBZ
5MANtVwAoCmnhGlx+KRXzCfGwGAI0xvD5MX5PzsL1tVNPpNDQPhnjU6JWaR3orouD8CkR8HyFEb7
5rgL1zP0aA11GOVvA3ZO/wRFrM4RW2rlBvA7stdy5eeFmm4rABFUWH85UP5nuY1taS4j8Pj6P5w7
buo9GBTxjsCOVm2+6/9ADyQY7+oU/tEMG8afwMKZluHewKtdh8MmC2LUB1+BYjYviFzip4T0Cd+h
RMH2m8n04K4nHj4OWw4hs0Y6b/8W8bYlhnk+xBkb0JUzMS4nXh8807Men2qzy5GJphqrZjgNgNg3
DkgjcuP/R6xPb4UCRh9bAxHGhaZgRxJs8W3db6HYI2szkJFO0Nad4D1+6KFe+RVfXyLrmN7akVBr
Oejpymv6PKhegn0Pb5VTSr/i9N130VJ67Ub6i19ZzYTA3ZXJxZZfuWuOKcOkhKv9ZzY9pvRZjm+w
RZrX/wsoYJqt+/IGMxFx3atgeZ0PecMDwdkk2nsgCM+0RnhgRDqsE3ybPnzD0Qmc5P9bbVedrSxQ
UgbNDh40IarXXdvVKqZq5G/YpD5bLoWbYcrOwhFpfpCYJzCM3nCtCYsJthq2L8aO+JkNJd0B4Wtg
Ocq4WdKIia8bZJkKuEfkU1MAAIt0izHnkzF0rWSCmisecABsfoYaFinqf/jTf+BJt/xzmwb3lq/p
zJV3AZrU3GOdFt8G4g61ITHrZ3lHPYiYpMG4GUIco6kVC9YIN+yXAq0VHUu10pd9QNMVXMEkJbYu
derVMmWNYnmRujkSwnc2CXrk1EZL0PbWvVld379fbCZKWqfUfc3g3PXxqHszdDTiLB5tTf72ZbcE
6q/X+uESLqZLsz3d8r6S7xI4TxZ6T9ZpxvfZ/MSlVWKOlQLM6Ed5E/bBfwp2oqZmYExyT2vtiBwG
1kDeAjI4O1WSljH56Kd43FRdWBBQXQlSBRVS46LB5zjg0NS+ps/xYWi/15gUvL+UVYpTX4MeLjGy
kK1e2v+v5QNJWD32ykjA/po7HRAY/N9nnQpNxL3FePaDqyGB2NpFzIh3S/i7gaAYYvY5BwT4yEgV
OCTOyBWDle2lxljLzrNf979/Pk6NG4CWn/2B7mEniHrcMR3FLjNIaMS5mqs/HrQRAGwej/qAMoys
ImJ/28pQ5sfBi1u2EdP14dQSqPIwPYf9ghCdwvBINRVhP1YAW9Wfpll/zurg8a4O4Tz3FuV2k1TS
oF886Z5f/txPclbWVmsPrbuR6QZFoFoXPL02izeikiuGDmAlXrLaLWY7B3on+UbupQehBwPPtxRV
VQPavvotOu3cWMPwSZsgF5MzVhxuvX8r6BcjvTzmkVr3tZBqrLt3XO0OeUmUl/AviiyxMMAZMn9Q
T5Cjq+PL5euwgLorkKfi14PAqTebFsVLL9IUDuqXaF9on33KfHgX72qS3yc+nwLchwvfRdudcmU1
v/uzfJsn3yXic6DwI8rFSANL/b/XCPD88KPrwxm4uBUSJpuQEH8eFET3/ND8PfcOhX3J2fG8jAO+
hXg4U8MFsgYJNiSErfLsn3hULSVKuvpzDFLO5ikt/GtNjycTv7dziYZy7xBOGx/U6dNaZYfwOhRu
qrkoSTMK3se09ucdjOPSalGuwpMTlZNYwWTEsEkkf43Lc4ALxAscpEVeknVOe9H+6l/WFvdFxrFT
l5nWxKTorcp9Dnf4R/j8cH/Q82eipAc0c7qUtEosKcN2hV0IR7IBa9Of7sv6HSkfwg+ERvNaivV1
VpCoO3yRJyLL/8vrsEKCss2PmmN2QyAm71NjLeYYfA0+taTfDHl1VbwGTjB+pka/Rgl+Vhmx/4tH
W3OLIFuWxUGmqAnt6FggOjme/RxdZT0gO9I7Jh74PMuos2eeNeQvqGTx4Ot4nwdIFC1n9LAn0D/I
qy9KXdF1oxJ0yA8c5JOyH7JHZl01DaYFFpnexgzo6Jr4dUbd3PLEJRV47GrlvJuRAcun6CXXCHYp
+dZvLSUUqOuOToIMWZDXi2L5vpT8vIDWxdTRe6Kg/ftOxA+jotH++fjH33bRV7nrrnvg8WklGNp1
Oy+6sUO3224rrZ/VA1a+7v/C5QtgHR76fa/zC+vkkwkVqi3+cP7PeQgFBzEmWDYCP4NfJsYwivQ+
iGcJ5BpY0ye6d3SsG+9uLjqzAB+43Ji1ft4oRjLyL+ub9ipZ8tl2ykQ8/v6VjFrbCfbzaGOV4Uza
S2EGY/9mcjuCrujbLKvdvQLnQrDr/8pAPEJvxE6PxaeShKdLcLyQHuOVxalqNrkbxuqhPl++FHAg
3SXIVZo5XRfWNmenT6Lvst1TJGR+XM0WQsvXvkMQwp1Wa6iVStf0AmLOr9PabyPozvvS2axxwDYm
QZuM5uHO0g+TdGg05x385NLV6KV/pIb3IvTzd6k6ZzUGeXUMTUY1zcdMK30UEnvZ5T2PXatMneLp
85F038ilF3xaz4DPkSUcuJgq70boi1rOw8qeaAjXtqtO9mMcCyS8sVegS5FelzI2vKzDPCUpUBly
jyz4PHiOuNd0enP4zszY9HLkPumYnhuMLrCHQVJwH+F80P9Y8d8ZxsyoVgR3HBWp8l0+lVet6kTM
EK44j1D2ljcDffexsnR4MgHM0vW6VHSFlIkDwAj348a7FTJx9+/mkTnP+xmDNFdJhtWEGEbqO6UW
PRofsT7QScpNaGluqRUTImVG84dZvNTcptK4g83zGovTXV5PuS2VS8UVHVwqOAjMzK/F04ZGsSs3
RnkXm90PHfLUrfnAPsPefBwPVz6FL659drJzpF//2u8RYdh2I5894IF21nsLIQdmaKYhIJMlERY9
QZwT2i7sUraWggOz0j1jU+kKPNTf9YDMik27HcXd6jnHQ5NUZ1RM7LtnY7y87L6qWm687WMOQYGo
QzrYDA7GBTk+nBByDyOXTbIlqFiMyNB3zZ9+QzSrWXQ12ceWaLwyGiGLoQLX/RectKrwz4ywu+Eb
uVUYgmVVi9kgax1oxmXD/XVWw7ykGpX0K8OeEPewafQniwCmzX49kSX6KhEeMwkbz0v6YcTEz63d
nRSgvcq+jeIMhUD7MmOobYfzKK3xDayOEA9T4HP9RzRwRKwfnbCtlkcqnUYO3RTUiW0TvW8/0T5O
A3BMJc2zwF1G+3s4qRE05Py1VLmow9z0KF+NRtnvynz1a5HaJWd26YlER91W9RpjDYwt4dhxiLYN
30Sa8oPDnzJ6qFZ70lHJDGgqjUcK06BOqpvJzqPXkRMRDqwbP6MI6+/+pdFkuGnNGMhmguUaaODM
GfpZRkpk5dkpY2XC91rZwI72WLMd3VvEjNS4Pg2Kpj5iJ3etAPsWx1vT8+mpls8WOqdCthFtgLBq
PSgMi2J5PUO2NblXBhbOmG1F2cWZGdQK5pxgWiyGn7nUkpRHRSmvpr2KmKZoyc0a9ViRatC9M/GR
Cogu/tI13S0aDZA/ZirzbFP6JuQlmzZ9stVc1DtfKtI9PDwbAheJMlKRDQwAR6Rd8dh9WcShgO3/
v4/bX9kMIAZbBgwJHrRJMqufD6YfhRLb4B4grgYowoCwhTs0rHrnrJmhJAO0FbzMO5tFhcm27V0M
tSMZsv5VpapqTVTGd20JB2brcplT8o65IXZit5Q/UVPvjdPiKiQj0dshB/sjfSfc1Mzr/2954MFl
BcTI2JsGEJSNezjdprQz11ZZuY5SbVLSB4cz+16V4gp/LX0JAjkYqYKJqUE2UhgVWWxh5gceD0MN
lE/GwEMhlmw5oAvnF+sHLb7yJirsRlBqLpZmibiQG1EGTBGOUPzQDLAAYOn/lJWeR/YyJ4zQpHvr
PuuVTh/u0Yl3xfhU7km++e82XOZiJqafAT53q2zYCGkwUSVH1LvkKhm72IKulm2T0NarkuS7M3Z0
6e+XJIsoue2IRH4QuEd0fSrDWtiz9ny+X3alLJdUHKPsbnG0zwiYuFE1dZhwXtOIPmbfGkKi6f06
EenETGzwqixqoBaPu27F8B5Ov201/4kuIYdGvLrW76C7IevgASArOdMdG0TMBBZtvPx8B6+/DEQr
Hcjjg8cnvHnqd2X3yMRVmYjEngxim1wAoIiohi/sVoSOqIQ5qrDREn38bZbhhsdHu8igY01FX8Dw
ybzePqOrOIWJUyvIp0Kj4+XrAdGkWj84iJ4ka3LU3dzE6eKyHkWjLGCxWy2wvgCl30tUmurKRWEU
rWJ9FhQaFC6/UZE7RAHM+aqVwRjmAlLGGtQ3+oL4Z+cGjawhsFcazqoMFy3HJJEBDbw+Bt1aYB9D
Y7qKkuVHpTjYjwUH/YmV+xYNMukXk8vqhV4cmDsdIPDqYWNVh/jwoTr5fTeF4yLSTjg/ftdnYzTo
QyGEGJU6IblvgBZ87XMrXsaIErXQdSWho2jWDChiM+5wwZLbk9z/UFPrfC9SAs8/qramGh6hwaK8
r5uxNpQGFBzh/Pleb+o15pVYE+5DXIsrJOGqgH+Tg2LDDt9Zmz0q5gLQ20syRjgn+zD/U77P2kfw
ohD2bk2WIgvcp+K3tYrXVbknsy3pKC0+Sz9t6ZCV+9aTyD3ZRnx1RY7Rzpo/WeMwC7iAf1kl9pDA
nzcrgrK/0rLsGyJKZMosR4uaPjeuFeY5Zjx87T3Ax9CdQtSqoG6Tgb2i6h05YPf/WhDQJSQowV5n
P9EvpGpIXKQ3VS7W29wvYmXA3uczVAwLxm/BSehoZRsPoA3OVo1Lx2pZaqrLF1B2IAxca/WJDpuo
dK90pHZKQxKGOzgcFxIOQQp6ZKDe0ppMSWPzTDNIXVT6pzdZiGcaOUP1gYv3wUDz3EaOceCEY12Y
J4zhZHcW/OqT974Xn3ecWqivAuQ2QY/J53BNSuEsPHAAuet+Qv8/MzRqLC/DkzC3wDURKso2JHg8
Q5tnrVBIEHgrOxaBS4Bdnulmc0I3Z4YEO3PR6w1jq6cY7WNYYKO3s+Y1o4bwMYYk9yfY3xlKb/05
54607mlbWeqiqrFWS5/0Ucynwv5/kZxD/62hLWZzpdRJOIdhaE70HVqo2CCD17JzBQEfclaDR6hb
zRjXaAHrWsMQ2nSap2ChLDAuWwjn+GGL7VlLJf3moO90AG8WNOY38s4D2o6V3VENQQ/dzga2KT/n
LvcpGDEVh8yLZoBku+UmzrCZCcLR5BqhpAFEmJ2Bk3KgnqlG1Y13BAMA1a2FQ6zfFCEX2T6hwIln
+9wOQdusa4gwoiEvtGIZFMyNfcWWYCFr3oXuOGJHmVRh+io8WRMUN47gmcTM6l5stUAzSrW/Qg/y
gUerAPqS5gPRxluj0l6/cbWrAxCOzQrECSrla4TAfCX8FKMGBjSbj0HBk2F/65+tVUNx+mk12Pek
XB9af9qgVjYZW7UD73+MGgbFkYiabBUP6ghbQUZ7wmp1/ccGnrYkhNNXGkBEqVnDEyKnGJPg0o9i
fX0BMo7uOI9m0m0Gb3fyRU7Y2PcsCwLnwt5p0ZInC1S/VkJZ7mVE9ASFULzr6qMkYXt64zRTZsbj
22yof6Q7dKDcmH625XIL+OOFfgiuAWPBOrVSPG/GD9pMdHZpkwrzB6VycEjkRpdl98xMsCqW4hRC
KcGmpYRCU2Vwa1bwkEAVa9Z/lt3Oq+GwaowmaChk/8JISndF5EN81PhPXmOniWsTjp4TyfAmL/0q
NswO4SZ4KN8DP8XEwb893I3EJz+lNy5EnAlDPJ+sEc7PfWu4PgcMjFOr9rpgEJUsoOqWvWa0RHAF
q5H+cnMrxmjxGRUmdL8r8oV3LTk6sokwGFxITeOv4FKlkhcYVbIRp69Vd3QMYfbr9uc+WejMnLg6
uAoXew650vr5k/oNhQQrg+sQ3tIeWYRcFq8DRxokr+sOtufBD95U+tP3ZG4oeAnai0rTzqLm7YVr
psVZFRZ+LfrF6dT535ADphuygRrB/euWZNfCqPIJvz7RZRYjU5esYocsVu1CyeiTkbXcWMRvsadA
rvwNfM+cJ5kicYKbUG+9AZLETWDWPdJBwAhAnR8JIA9Vy59XerHg+m3IEo3R2tzV+pcti1ZJ8SNe
1+soWBmfVeuO2uHQQpdPL287Bcn8590ERN7vZNda2YmHFzAxTuglGxVrFYiYjtkHO0BYiC5d1FOF
kfrceOjmkCPq+/eAP3/ptSFdT4hRiB5IKrQtu6jLh5icOcr+Zn61cqT5ToMi/Fv9D7ANBRhtIaty
QChGsEHoheK4wh4pL0rCrSYWRs7JbPjOBR0XEOZtu6uG4Mdr7qu1QwAWU2IT4F4LoW2Fd/STR2rE
+V7avTOPiUth2eVjXXXuLRaCPzdEoXLiXRk5rEG6ZLuJ6wcstyLlNfXifU3EdGxs8B6NIJpxu/sP
Eglwq1COjMb6EYDXV1ec6vwuWs2rOGgjXpuI3DKTExSp7kJv40OubrdWA5Fn68aS77ij+M6pYRQE
DTgr7zact7LPh6GGaByKVrk0j6fcjYJCLIxEY6EI93+gOn3rnui5ydOrSxkA+HvZ5WEUPPz7aj8k
A9F/Vy6NgjJtrtviMPE+UnGzjhi1cO6AR5UtruE1DuKtOPL8d2cgu08MIBjn0F9XWEqlDRQt6FpZ
AhrBMM3T/UaFOR4+UgbfRr5uskfVaJw1vznz2lWAIzqvjm29nXI1WrOKXMBYdonjKrCV0plVom7B
5hc28xQ5DnSffEtTd1fhdgJVlKXOhOee1GW9dM89Sum8aKD6cE0LRS/VzFTQe/B35BOfFsUwMfht
RgKtPi2hz/r/snbj31gdzHFEIXlhuoye0KwpyHTJAPbS6YQAMNnNhuHqL0hQN8OOAtJ/G+/pGkBw
EtqHPsfR890UtAOiP+lLYF7qXMWx6rIIGIpy6bJB3WH9bz6aiqKOF+vVdJ3Hemmp5iYVlI8JyGqL
PJCew0oi03bjoEgv40B/5h3XZjlSt+x65IfSM9xpIWEn9r/k9uve6LlmHzjtI3r0HtYJfCrX8WZe
ZdeILxjVtsy1bQUNFOLHbKVR6q6JHeL8hheEqTDqZY497kBvuhykBAt51gajCmdITEy2upSWW2Oe
KsYTWkpplhtyab4M28AXbI/PSRBhJ1U97IIRUat6LVy+Ir4rL9zG1sTrxBhz2oUBO9KEQKDHPdUg
c+E/xQVY9EZ32cn77eYy78R8Kuj/FutQkWW+aJjgOOcscklOEFbrNPKpm2/iYHWfFLiHyL0nk8Nh
LuHFEWZPVpDvOF3UR5yvevakPAGmnInuCp62PWkIPxtMLJB/UNDpUCAksuCGuhUvorHIVtM/ymlN
djg/5cCRkm8kReL7MTHElhi4fvYO01+y0oXH4ScdqCMGLFRcW3KJbUA/09ELRq0VAs3BUnsRFSA+
hyWM+XWpguAryzW6oHoTxUgUJ/RR0SqlGhdl8CbAU07z0+7WRsRsUBZwiQgN3hXHed8uckXzdVut
G69GkXVk2uLOu+V0YgjI0i0Va9LVX1QmUMCTZ686Oe/prBBO9g/ZKtXRUHLT5AndeR6PVEgpkWK1
pwFwUOaE8x+faj5P3EZqEPW0Ot1zo67m7d4oBUNzNkII4lz9qpYtBZkkqsvHLyYYZPpZFMf4rbW4
TCahZw8NZkD48sjk6DjSghxs1BG+VR4zTvrJUptXGnQaIbfRufEHfvEOVsx4SXkE6EDLPyjq8I7e
yxtooIMidY5emFtabFNXAg3GIib5OIuqSQw8np/E2jTza7sCJcJOJDN8tZb9mbl6xqft6uwNtvMe
XRIvQxQcRPm4pdIR2/LO+LNLelS2EwKXfacD/XXDNogqBEEsvUwdIfd/LmFC+jTPXRwTilbDijWD
y7qPc9Ze0lXT+S4z0aI9Dd6/A9pJTfMylYwLYOGZCbH8RbY+7SDFS4lzqZemPDD3If5adY39IfSx
3SwGFDqKO9Vqr8d7Yb6JBt1aFSELfjCPhrH/aMoCBAoJD495ArvKPwXmvA2jWuIf1Px4R5dKS50D
T8EeIqGZpTihmuegjYa7kDNrboHwhAV6VeEAZlPihU4x5nF+X/wTrUmlFuGPU47z6m4d8PNd6JXu
EgJAOegzTr0AgtsVGDTRzUGfU6M5lrDnTUbfKyHcfiFjIwYAFjM+7qc+eQY5jHS+DCPRJknRi/DM
+9+soF1lhctuRdXnfguUdtal/lV9reomeY6hNVdrGVlUO4sTk4QDR8d6SSJDqS/nOnR8WN+i1/AG
6F9Khw69CYUsHCzUFA4R9OFqsG/4ijesXhpFzKsfj6YTr44Yh/AqLZ8RMlW7lIL/X6OKkhdx/dAm
6110t0zkOYfZ6/kTDeXPL5OCIocubFMYZzTEH3sAvtYSbdEObcz2kvggFAt4exELutMitzsBGogU
G+SQDjKBG7WztURN72lPjAMMstwuR6HNedc7OsQqISXd/Piv5arshXE6Ov2ycDPj6hTd0RFGdBk6
36QY7NzI/zXL8gxgyScqjUBAOBfjsEtUkY0EjRPB4J6aUBOWEPD3KACKtnHtMWwCCESRB2rySWa5
YVUXucAT09NlNoc7abu3TygwwNPTyQWOodXYPTLVkH7Hml9nWo5g289JmtYlWt77ghbD1O5T0Wpp
du4Ub72dMyLkX9NifkoHgjKqIdRiogtyUgtinvld2qKSRrFWvSOlWzZY5fAj7wtlyMM0lREnK8j7
Ps52vnsxdAX2doIHQXWg/zXCTIvz57x4rK5ZqymhI7XIT2EPxtGMuBUHFu98xLRK16rLCiYc6YFI
ETZ8tbq3R7Xw+U/AS8KvFiwgWMTEGQ6/nGH8hgx6Re0qoZucEQveZfnBq0G7Gnor6jZM8N5+y7qc
3jltf2Cmi62LFZTCwVWZEJHnYgQiXj5ZR0mCJIMAVW+BJsL9Rewpo0Vs6RXC5tqtYim+Ea+dlgcL
OTIq115xI3rQIVLGUMW4cfZQezn78v2lrplzpA1eKw5lWhouiC2WsKWvlM9q0JGG6yWsn77WRF85
zoRnwQzoDJjRqT8PGflD94WHoO7sANClEVsyfAG2NeXgZw5ylzo/N5IaiR75DsKogtJAH3DgeV9S
Ppi0Ma4UIKXeNlLh+ebZ6/z/lnSCRej+nKGc1o9DSsacbPRSjjzqQRtRGAiMWwo790RjHP+TNUW7
dSbW0pud6rRCB/clyVHGlB+Sh1VPTh0Fq/z7yb5QGli+o9bDK6ML6/NctZtQ47roG5RsK0QhuT3w
QWTiW83ZQm1QNhZf7OcKWaDAZprSbpNrI/VQfS5KnVewWJqYbSRmNBjiLUfXvsmxcVrcgjRYkLVh
ZyF5SUkMuA305x5lZ7zyVA0SZqZVtYJHwjrbzHGaPcYjEexeiauxJXJZRheaIyvdC4qiYaVboOaw
TsnqcGngp2+uITAPGQjNvz9xEhwDC7astOplq5wwJuCDrRRpkhDj4tcqNXWVtmbpNDqraiXRkxWH
Nqi/gEFICrdW8wKNuco6yXvxu5mus1S/yBkiGO2XIV9ulRx7qQwr3U10SWjAyNteXxogRiWYIXMi
ry+Qkw1DmBv2KHkbzcdgFu76vcWABACEcQTajnM/V4GTZsvznAosPKYXGXBBk6mB8ej1JOJIBFAb
ngIgxU+h49HG2a1l6BvY0bO4HxgwrBtZR5yfVYa+mauEY2X/KJaZjCdfN3sI32hKdnjBsMe5Jmgt
DdJ6rkaLuqtFsXn6k99fe36XdAZSqOGg4o67WGbxeEUe2lieeO87ef340XCzW33dlguPD5M2ElmY
5G6LyyzcEhqDiNzmKpBA/tmDqE/coQEow4h6OEe788dKFtrXN/E8gteTBMXu7Dv2gpRdu+bJVBQ0
tFauTD4WYAtHSb9zWEP0TcWRDXFkybNDcDcirnOnfWnp4D+kpunmcSTXsfR20bBL3jF4IoZEIZyY
QeIIPLpc6KogUc3K7jpDy/eqWxSSLp6xLBOnSd9ZUjTVKYxqEPKTOei4Kr+dfGbxdDEcthccm0AH
TaRjNHTlAsWSolOiixa5FQ6S9LxHDfvJRqLV2GHYJ3IgmRlQICdIRvQCxKsQYvWdCbPsBrVn8BJL
0BLz4DPn05uZ4lZpoul8jxNgdzkLZPk5mlqjGYNwaxlH0bpcBpyUmhNzLEP5pKLM8neSkQMyyHcK
9vaVwwIPJkODeEV6FHWYxH+WXb9YeL8j0YyXikgzjXF9r+djyzoLZApXz6Lqb800Af25WjHwdEEw
Qf4ahnfib54EjaZBRXc6dMtpxYaBgHPTRLLOaBycKZ1t8dyuFPCV8Gv3IVo+vXqkzSuMAucEILfD
0+a75IEy5JD7AvCvyJQVyOS2hQk1FzY/gWUDVQibz+5WC+qkxu7n9OFZ4EtNq2SNiikYF8EkdDuN
10gFvFmjZSW09bdtiaqdfGcgbv9MTnPsTiCCBv10r6Lbd3/Mb/o53zDO5NQO6jdKw6lSUPDjIXfj
3vHcgI1wwtffSqwU9UpwDg3B0ZcgKR9Ike5j780RC/eRaJldQxBaCdohYKPQLj4xd3YCq9v9NgwK
lKkh5cZNxljso1pgCK/BCkYg1Yrk8slPwmPFVROI7TCuwgt5NmtlY5Mdk/xA7dGIqxc/oFJbFg0x
rSmyz30vZr2W0/GDQiOT+OlNvQJr99ve7f/Q3jpB/JqQFkmK5zXHXQ9s8m3SplnlxqF9Luo2IJf6
jvOE/JYYTNtyd6k5EgS88849BZEPdk1NELKiK+3I85YtVTaIBn4KH+ej+WrGcPiftwghvDrrtOnj
4usE4QFckASRrod//oPj0kM9BVXf5LmuLzAyfOt1i3Y/YhmrkPFNZjBuK9MaBUhIrko8JwOS2DoP
4kV78uT5wGxZgYnbs4C8vn782bFV/t3ZJP7Ni7wDx53H2ZizWGMw6MXPPwaZCsPJTbGM5dcbFH29
xRUsyoB6Ae3ll3Yd1Zn31C3PZ373CIB8CCUUNxldM+mPOUtMd+InyM9oL2MFaqHv2vSmKRkeVESr
kxggl++62RRh3Bh4a4YB1lYKWKS3ubhMyYyhOXVswUQnBg4yleFj9WwxS+GovXLx43sbCckpnx67
ZdRuwINInBuKSQxu63WJ4Ed3AsC6bDNNBlAserKhldZ+WBLiaL/fLgqLD3R86uBbMinukY8/kYlC
7s0g3Z6zvLJ1d3PvwrmnVPQQLVMiDdG3EjD3qagI2Af4VZL2SHynPwa3OthTc74Vmzhz5Rultyop
thZP6OfTuOxO8rwMQ5gUfguFyPvzsWntlNFSSesZBB1HITm83ZjnZd3fAxbHTqOdvttX1EyRxQAb
LWB5js1tHh9qeMeaqd5Z2owxUENpA8vXapjItYctuuhvk+PUfHfVXJzGzhIzSV9sRKb8sYrlqk4Q
ypis0qCKQxBFS8JfOiiHqkhZEUawfV8ktL+S8rYBQG2z04vo17efVMwwavkWmyie9nxsJiLUJh5Q
gbMEuTzq7amWUaioP4dt4gk9oQ5CZAj/4d0DtpmCqqTMTr2mEOaO9u7aNLN28edifrXuXeWWma0U
9NAwr6vk8zn1c6RQilSEjKdwWYJ4D9cauNkPBEPiUvfM+uDaVHxTkh1I+Ts220V80uOCn9Du63wJ
Dze9RoDtrH2iG0YyyAxm9mEDDvRiIpO5BLV7Z3T9/95NVcIGtAOGj9VrILGv4vusDHaIBazTPkg3
ZVAV2yWgFgwHhd7rhIVt9bgPqONJHRgNoKDA3qi15ck7epy9/oYFscoOmL/k/RyaMSNntKIHMkyS
CP1BZzDiNHhnKPdLK5f7qxDN+POCjnwz5tjBfprFYs7ueREu5Qy+BeTsHUVDstVo3J50Mx17qamP
wbH3rqW6eR6zVSnbTN5aBIVT0xYo6rf4UE/POhyC/hXMBktzHQg9naRnJ1u7HOulopOJSS2M0sO0
KPuUSI2VJd40h9T/X89hnIPI9WvypSwReqmd6qKKSqkJgxP83YmjdguVEmKONDIwWlSpbkLapZZl
4CTZHvSzymxOTLI9rPPsAHSQhFzdtO2h5mYqzp2gFeg7Fl8iwgLj6MWGX4rnL+AysV1xnzNGFStn
6qtPYqIr2Ydj+4QJq4u9E6O3a5STHApSH2JSjAa9pilp/bN9xmch3z7t0sh2/uC+DwihrdhzsKnR
HDHS+h4yqHzQfHsgEvyLTzNLe8Smn1pHtYuj8zKoPoz0Ubm6KHVmfEcz/MrL1XuIGg6AOwJIuz1H
77dIefoNZbpt70gwBCnX5jCJundv7SS83kesY+P6KQYxqKjWh1Eri1i/x46LVNyD//sR5T5Gi/Qw
gLKSiFEOFgo1fAR83GAq9ZscYR67C5iNN7JVWYQHmCD3d0Mp+Js6lO59Py4Fwl+71Yg1B5N5h5ly
8ur1giZsHDcLyvEjlYbpeNNGP3SxBDuaODzkFwWpcyuF0Mro4Fl4DzrqhzTP1E0IT5uggtUUD7zq
NHoYj6PrkJXhwQwQ7YhSuHVKeybhyyjiJFw2it1a7Cn9SAlVB57TTbQQv6qjNbcv07EQWTStXnQ1
cyn8iJZwIj+kmsIsCfuqtc1fRlEaHd/BrTVP1i1pQzN2svXHnSdNPuvT2h3tKGIIFobhVS3Ptf39
3Fal8EzFBDCKh4aqRGVEe4QITsLeLDPygGWmDsUzubF2LkvOPiLz0yGk05n09H8aPSwJXq3ZWbG8
mnNisuNnbWOE6Ww1v/lTAxlpW7MIWmZTvYkLPX/sE0No5zlouGyECZAeFZgC4TX0BAg0J2Oes2sK
+fP2bIqwjxRWG4CtvwG6QrU5XhPkNM8JoP2v4eBlDV7gDymlm2t9jm58O6WNP5IVUBieezfB1Boc
miC69H6cVOLp497MxKrc6ejXJXJLmTEywkjE6kLlZIGXtRtXEk1WcmiTjUfJcMU32y131Pxs85gT
bBLWtaAijaj8J3nOE1xWaeAue6fzvUWEqQK10G7zoDeQOCnl4NTjNfwb8dyqAzAn/+cnMqx7iJ61
ggPPMVoasEVoFgtvvBbx7LtCc9JrHrCukuJTkevYFl8gAGGBrwLqLeRbwk0ZPxLEnsaFzbZ070N7
mCcqwUT/JcbJ/Iof4oA0zUhGTVloqi8n1i/M23snfp3EZV3G7bQP9RbO4dMYrt9wJdZVB92VXASW
N+2tY5RSFaBXTflmMv5wkn8GFkZVpcT0kAgiEnt1maOx864L4AE/BbKFOk3PDYyIm1a2uSBp32x/
r56rpzB5hI+DL7uOEHn09IqlA7HEAx6lyM6WwfRn4PZIUbIi9kKbmwS73HfNRS7tAZsGqfFxSO+/
PmHib+GHWveTR+GcHukWh//qfLUAahP12fvAXxmDjAZr3grDBgqVhnxbr+aFrz6a+ocGzwa73oHl
vJIedJ1S5CZJnLh1mQCvGRA3zlCKdyZGfNMD4X1ADGw9IS/G6iob74GQC22nP3QLnDSvbR3LqZxh
7/G4SXFsMqfEPUgxC1GLI3x4sxh3EHh8V3bM8ZRA4adkJEUK7xpcIU/yODj12uwqx/McyoYM72//
+QzlfIcHhTvVr1ZyoJ6UWJZdtiz9lf9gZhld0KGSqKMCckEaI3UGWd427738g1Mx4PDAJQ0RMvfT
MLgeqqUNzDPWfqYH0CxKYzKMugdNgpGNtK2CSu/EQXAVQteqxJUMW2pxySJ010qgIL8yx6qACena
TYzUbWgLJoZk1ik1vBJCq8MUbazguOiFrg3PBw5cWyj+vhU5N8UT6oWPrYZA52eANlJ+ggrjY/YG
G56cwZZnEIsDtqGO6jr4dz+T/Wr4pCLCCz8r8ANiU10nEK+sCJ5Zno+F+ueixE5j152FULzAPtIB
NIiLXVu/C/nX1w1RpUv3PdbGYdDre3gAQ1iFvNcl+/0OAXqnI4IAUug1soUHzzyJpeQNOxt9C5NP
D98kPTtSrQXOtmRD9bWdCbGJ4m2RDVueLTWPaYklq9BgRzMyR4tSXHx+w2HwFNHVVpdb6c3o0UXg
NUF+tyWST2Acq15gCPBr5NAiqsIMfdQsA8FuoI8xvMvasykTDChjTHBIrOAGT4WHJlqAwTbFQNHY
GdCPI8usyjN0qq6AIA2+TvN9CJSjefQLmPOenFyn2yzlXEa35LCpW+LP9v5I91eQsSlx7GQ+nE3D
T36Yv3NdERRjN+OvVOSFUgsXgCbB2TZ2CXLxjcTzPM1jW2no/82qeM3GfeYGuhijjnKeicMG1QR4
zcGeBvwdLej3f8HM511O4uJ82jTtxgZjgEEY1iXVZCWLfk4lNKhP6fjT4Kt9hagmW3lbo+nWTTFL
mXP+3c2ByzxRzcTmaehL79FoEvuZzJet5pM2R6WHrpchsggDPUiNC75au2N05xy8BG+5gpC6/OqC
mr5NAQrAFad3uEYe8MRC0d/FN4HedZLtkAG2y4hI7tCjTR+a7ehoRqZ6hOAYSpyoCxa9sESaC8Jr
xlzgkGZeEq0g83tR4re9AW/zALsTObztHXQmsbDKMtThpV14T+/HmK/Ww2vUHjAq1KHNMixYcGDy
xqGfcew9uhW8+ft8yVLaZKiL5o2d9l0ELGqrHhV2/FUhYH5zvQ0AndZt4KFs5HzPKQH1LncDGkZy
E5SSWTn/2W4rrJ4/mptqplWvUPrigbdwGHyuuFPK00GJtCDQVOhKMc1J1KJ31NPgHyWkF93WEkhm
BFTdAeea2L5RjBckxZV2u07bN8datWPaZSgQiXAhjGoa3lDNbRkvqcp1KPizHGdr5R6F4UHr5Q/a
+U7jakNbs4VAlvLDTGJtV8P0pmsZiIM/8LmJ6pnLC9a+H1H6e33ly5039qjHv8catwq/++ISkio0
mkteQ6W25eO4UM5yt/QR7utxNqSx+oHcn0qrHx9RJ+M0Yg1SRXjtUq9MD/lxmnpt+mFrHUDHdX4A
Ag8mFmP3MEtMPhykvXWC21JDq0gkmAPA9beRHsnjIhZBblPF8eScEGd1LkfmoCyU8z/D/r+8cqQ2
D4YOnFj8YwAsPVtl1iTchkITA/VP142gkpRm77deCcBZ3Gs3qznkVyf6hWRM9u0sHUYxg/1ymljF
BumG/MKL2qBQUIJpAVnQysQYq990lLFkg7oElD+1gvfqgUC5TegR741ivNb9pkG0H+4DzvYIyPfC
KvdbG/W+GUV/nUYgXfeKjfd+31qNY+aqZTatBWO8OLwYgC5LVn9qvMi+gYm/Ltipw/7xj/ZjQq4k
E7P0mHcKB/zxrRywKsOhc+DyYTbebHh1BwKwX3PdIeweEkSCgQIJUuxTE4tZjYiQGr7ogIhKeqyk
LqJxc/eUhJTi+MQKJP0TwSl11P9/Tt08xtPZJfyBotiVJZ3g3UKhGEIOorm6e69AGS+D1cb45Uz4
NPXXFFrvZPJSRjxvosrrdasv9dZqZZiTJdCplqge+nfNuvxG+Q91s8shPc6aEHOuxDmPgxvC13KC
3ZWYEb6pMzGstut5Lg7QfxRnT3HgK5R6Hr//A5/zOE8REw2Zc7bnUfNvW6kfjfedP2g1L2eutdQF
OkkaO3s0IM2CvmjSBUCed/Tpqfj71FP3GtC7J8gYQ9JnZLdIIi594jUARkBy3lZ8gcWOSSzeRV5P
VWdqf0XHeJrpbEFvZ0uzo1bwEGcbYU7J5ojAOfH1LwsPQvl7f/vcUdRykHvi6Cd558tPl39BE6QZ
ls0/rwahX3tAjU38d1yOiTqihqWyQL/phY+wImSQhS5tL4WzapXCwuLRDxKQfyhDvuQjOPlYTMlb
c/q47hSGFJxUL+uei2vOjfTF8bnQ1aTB+ojlp/r3v0/Hj+9N01rrXRGnlohgmLjo3MAz0dwAmkGN
Fou4h3i6ZRxPdTJg5E9vj6Hhp9vJ3DVYqEB3jzgg3+ehbdIo6SljMF8IW4OEiSTRY2TkCbEppUr2
DD7OYCXmHrGpTxGn5+oqayv5FBZ/dQavx7R/ol1pQOK4Lwughgu8cfu3t/iSETUX4e/Jnni2vdev
47x04iZNPpz6diErvKGAIcL8U9ImbFaMpCTdMWNzQw5hyqma9fT2VhPJ4a/M6RPOjH0yngT51nqL
n8Lxz3hB+pv3wpTu540EP1FrKXCsgyQkj8lwdVf2TUFQKgEqZOxsWwPUnnrwAvBgxme4sP3+JIkB
Mz/kSCvnmKerK7Fa+Hmq1/M6Vlq91DueFnNVD0amttApFm8qZrQTsulfQNfZXxFMfsvFhtObo2pF
FWwNBs/q/OLMqWxEOiay7B4Oemm8iKaUesASwcbC/MDDjqEYuZXSpx0tzEKjz8PFQIpCuyF5Qldk
bophDtdUpORewCqTS88WflZ5PEDgCE3lYuUDeEYqmlnc/3yNz1cyoangez785vBk4+H3SALAEIRy
KVU2brnQCGEQOqUSni/kQBUq5NdwQZs1UzDfolLQKorF5kj5rQLlHd9LJ6iU55aDkaCoUsCa4niM
Yd9EkukM5IBsHz8xcePOaL7MHmNLW8G3R8fxg6ItHKUuC9DLIh1VDBzAFT1y9TVql1shY4RqI8C9
SCcO3vZybWNiItf6xaGRLxyuAMtvKP5w6ufgJDQ2k5slAqjsTQMlAVNKaaERsM/7jP8XePBa7u3p
+tY7b2G3enwQ1OCmc+RTYYGrQOO1J/VxIcBgYPo0cp1IUJC85hLilymZMyqNXiyaj6tSpa1sDq5h
yAe6EDbCiN7sQRbPVjZOBzbzk9UYpliIyq+iibzrHvFXL3Ym1nte+qxsxMSNcw2MAz3lGJabr3gT
/JPVv+rPpuScdxExhjoQIN0U/X/vhIGi6UYE2n9EB+PMYxB7d8wWQ/1uSw3Om24tKmVLUqTj3Lzv
iMgGpAePQ2fWU1gmerbu69/+i8GZllZJwnH6zIY8BTfbhNzHOqYPmxkyK2JadQDY2989h/gaertx
Ch40ylBzBW+8GNvuwkbki6bm64b+7lfFHinKue2FCxc5EnOh6IMM6g7/L69TteDCbnTYs7uy98ry
vQmEl5+vnyJsbaUWHYCBVab3j82TR/pUT3IRcfHQLJ3ub8ndojOvoLs879zn0XdMnsdZeKk5WCri
hNG05I2pfYSvsH2DPmLWWzK9NgD4aAGzVi/5R24RyNcse4DAYw2dDWgrQS7ktLpvEjjjSYp8P1+4
4t9HIqIkexvSZQRZw8E/AMmfefhbMMt7fMvMvER707l3p5T4j+cS53h5L5paF4f0daC247lHOM13
RcghYZBQswirBJNwmhIZrsrILTN4EH7u50enf26yGrBPGh2z9m+N2KPKM3gsBq/4HzjMvZaSUamn
3Cgzo9r7IxUiz2Hu0oGVNkryDwT+gXTIqS+p+Krg0p/I+/zMvk5cByGNl5XPF8bXiBJYc+0VCaZQ
kXmGZpV2mqEIdnwkeKxDvFcO4SHlneh7pSvIA9J/fiBPaQuAN1+dze+FydcvmdQY6KZggEecxgXh
BcxCNbHvmbXaPaIYjPBAQRBYf3kcmG2svzhLrD0v54CR6jDBZNh89SlKbfuYc1l8nFSV2EpIckA7
aC8m38LUh9xikC39WQBmOVYZsKwHW+poUM/4ZHdfZ5c6zgnyifhjAE0Sgvo1VFAAGD8Q2Wpnm+9b
ckuNl46yIfZuhzDZNQBSc48LLhAEULIPDTdh8kN+1pOxqy4JDe665FVucagxrB47cAI9txpkxXjl
XNdhFosm3IeqYryffQFY+mRq8xl8kVdZfFebbRRrAi3gMocVgtyhFpbrSdgFyATnhRhE+o4AvEOF
68H+0MYeAC256WMf4mtJ6qCPkYYkJ9uEu034XClc0ezawR7cl9iFDuHKYQHhFstWxTvmGXsbDNaV
tK9O33a4oQzZ11UCsrQpUZeZ79EXWzo27Ko553EdOSveXebeWtD3bLBh3NJowtydvXstaAtJUr6u
K/vlCOu3/IzXMl18jse67e4FFRtcR3Nn1vzmco24+4zuVgS3gIRMw4dMCADEBnoKEnf4OlGpa0uf
kYE7RQD50THzow//nMeSlmxSMDNRfo+14VgY90fOqr0ENpGBhikqwatbWvE6lTVDeWTx9QGcLvia
A47U79yTPn9RMcZcKaw/7Iqu1wA0sQK29yBKhI+2mkgaibwmAikLoR3eTq6sCNbeOTPLjraui5j/
QtxBhldKgE4DXEX1ScpXGEBs+3Mqq7BiPdfolu6lIuBixBx1h8F3e0aYfEzpM6M/tRqDBaqTMYAE
w4jY1tBBgIL1js2pmXCDvg1jtDwxyHKHAMhXK1FCs28ydosxao18AGvWIaNWi3QnoJOjbSKOU0mO
MiEbYvkSKoVOG3tsFnBNOkcQtOvDYHy5PMTrIuXCmhn8WQ2Wc371y6VbRsszsyLwfpYAbsB5bQ4p
gVDQoA3PDMI3Lqfnj3TcSq8mXP1ZAnmqCLuDrm4PevhY7Ojc3Ytn311XO4v4gA/5z1L8b+ozAR03
9zN6gLe+bsdYN8dWZXPRgHRHMLjqEgg6JwesuWQdGXD0Sv7kc9OyAQbUfUpkGfMYsB2xIzxTQvwB
OA2weZ+MGJz5ru1rvmkM1EeCA0ZA2P2T+5/HszJOgs6eJahcVgG9bNlTZU6lRXuU2f9d1K8aaA99
7z4XUc1DHXecY3Kme5onSXZQXZ3dG6aTRJqG/efG8z6eZFZY1L8T2nXeHg9SCuQnTOvMoSEjfxcn
mSK8bnFnYks4VUoF0bULbZjQ0Q9FnliZ2m5fJeqXI7Gt5zrrqoMaxzqBuW1kwSXWKxQrfgyjcZl6
jstX8/xUeKS7cWKfuXTbBdHkaXQgO8RI+TiCOG+xkPp8NHXjrhhPbFbOe+5KG4Qq2+21PWa4F12k
yVxeo/CmGI4S33RO3mQrxB+b9BXVcfFvI2hwSoszn6blZYzo+SoagvKmyCPN9FePSiwdQ7j7cog/
3yln4+gq8Y+OutpZsrldtdY9f3LOwfOxKoANfP1OuwaDgkZqNS030EaCcmF+P2Fjj+uSpOK/euDe
2CWuTb92++BGMfN42fUv5D/Bu98H2qCTIpWwsE0liY4wY7nBGf9aR9SqGRvn/SGor9waeC+s/IDd
A7t06s1J1InA7Im54h62ZSgAKkVh5EIkcU7poeCohS2ZyGO6fZtiacBHY0uOCaMR/HdQxCojILp7
5ooiQIycmzwBon9XfvpFiscMt/pcdCSkaG00gtrgFQ5JHosyly/XzWbIiKoI7pQjmG2yhzDCOzH6
CJ9rnYg+4iZzLkriDC5KhMXIN/rQM7L1eW79Fz/de7aX4n5ITAQc4/LyfYjt29Rsfjk/eMa9iayM
8OqsT4zIhb5rlEnpc80gMGwl+GmV5Oenlwjw/2Dhp3DSOw7aKKJ//d+7vYEm3H5mxEk0GhGv/CJY
g32otHH60lhZoxSHQytC8ubcDfqs2y+ZzeAfuhIghQ0E3Pg2B11ujAA3frri5TywoV2f6vxykXMM
098qLNj6Dvjn+95NjvyYqCduOWL8rJ4yXhin/GMTdpzXKQJ8ZhYAOz9luOLEx5GcIjEMlI/9fVZL
J/qrujUHIQouSMxzOmASghwTqu0OQ0inMMa5wvJidjYhvRSNxgwmB2bgOUGcvqrt9mSDs/x9fVgL
58EgWkMusGmIacdHAEwGXnjaSa0hNtTPWFq8N2RG+Be9PCpRflTZHot3ugRNLsqgIww23x9pA92t
KBCY1ZJ0RaZEV4SdkOE04iL5Y4e8jMIIqg4tDUk8I7PcUIP0lMCpMjXiMnhipDgIjMxldczAnPVH
iUf5vGaPPCn3VOqLMNCpkh8iWmUSKdcGTnhL8w1S+jovV245OPQGMJn2lBppAqa07MGlrfTy4dR3
qinaM4u3IqPB2QRnlbvu4HgWUYBLC4f1Bt7OeqZCpYpNo+IjEYdUWFxYDp1TU1qevAj4WvEA+bK8
Mk7sEiHSSaiilRsT0ovdyegg4e/0TajupZ2uyWKltBed3z8FbV25oIkD7caTRJiSOCRv9oHpwX5G
JAF1/lk0LW/LBGRWyPdGJ70Da1n9tSaiL3+Pc3X4fJSh9jCr3HSAb5vo7rd+tkxuvD1qDM2WMslk
mHCLWbeLmv6ChmyE+xFr5xr5BQS3RftC59Cxa6G3TRQao8M1mOQ05pegJm6Rpz8hei2bs/dtJpG5
RJEI7XZzpZDy3EtET7bMRQq0PlvLgHthS7Tjypzm68NnHR31PrnkRT62phklbriKP4AQ5vAhur28
PtdIvkLApXkczYU7ZZ2UgIvs9MwKOKMKtnqQ3AeHw1N6m5keCOdsM6fAe6oy8orM3fUmC2rVl3Cx
r2yEVZXVG+1A/0CsVX9k1qtxcUaYCYn58UNGoPozvLuxKNnwcPhUyoaIUW8kV/O1ecmnKlben508
ITOEE2RXzB4As14JLUZ3cOxmJQ5ZgnmYvO+wlCkGEBAjDLesC+MaVwou61Odr2qPBLimbLLvBVk2
x/3Zkr/8D1WeWZi9QMrLuq4yDq+yvSCM6XcqNpidu+/O7WeeoYwKVX5i6Zll8W9W+XiYcxFKljkG
xEzPr032QgEwT9kQWUzyUVRdDqGPA0OseovKYwq4zFWsoUG8C5SJJrFalT1BTXzoPPOSSR86Kv+K
QC/deQMoX32iCO2tgOL48zbzHXV0opJrArDJVqk5MnfwFawGhYhcFq9KDp9VnFVljp0xwsDCb/xA
u7eOKWE4CHtKcGd1diTakvKZJvzAtn00hq67dyb+8iVhxZU9ZIznqqBgjgzg/uEohRl9jEFYIdls
XNIaSjunm9NuMnsV4LfYbBljxvTQ4FHL9f7HGtMTuiAOYdQl7Z7d66eM+IsETM/kIEllsoWd7TCo
DUl60O+mcaFYeFgREuOEYrcPoF9jZOrLy5UQubrjOwTRjKbdO7bGULMs1cWo9F8Ko5yZGywWw1+p
nHIoT2h72tDyeXOZ8+PCIDQm/zn+/rgjmCaROvdWh2gGhK+0PAhouKIpn9LXMonBJ34PJbLjtngD
oXv7iHYedkcxolLKBd4cFe1bbSWYC1PmR2qtNCJVNOLGUtgs6ruo12mEGymVtea7ETPj6bFMDDAH
DCV6ECEPZKajIl3QikK/kjCOdU9XVUFkAY8ZLkpWTFv2USl1nVpYQMfI5zUYjAA9bo2W4GgZuIIF
ILcc7Jgc00Y4+9Dtkfd1sqtGOa0FS5W3YgeIaXdbkRef0XBjar6DhSmtzzaEEMxUpIaRFDrSbdu3
icPtbdY6mnoyWuYp/ertUOJHUo9FVzDjXlH5FCEak9mBUH5M8zDoAyM8+vSzF4cv9E0lkdU5JKPC
c9jzmM3WCQkFeqi1If2/xz94JVB9tUD/8eGNRTMxGwYU0jHpcz/06XEI4rYptN0VwT4KR/0BRgXK
2hk8Ng/2xv8eoG5pxWwnJOaWWK3URlv8bLcFpzQrV8ie8P45h6mfGAveVR29hjv4CDc2FuVuOEIg
ZBcv7BQspvylHKRO8Qr/Tb7CwqinLWmrXLP6GMjhKFs6j/LLOAi0jh2G5OKkywcwLc3gLaMltoUn
0i9HUjfsuuMU/Y4Zk82+HzorTOQc5+2FyESwXab7Ch+3lH8nUKOIr9i50fKbPCuKzMS+V1GUEqet
+Fh7CTybjWzqyD91a9uvcolDlh+I67AMeqYsr/C4D1xGzFJ0P/WakD2p2hpgR2F6bomAkZxdIDiW
KNi0aY7fVFpTa/vLMnwmhtrjJNvWJuro/7LJKO1zBo0DAIL1ztEvlaw0dlvWcXM+nxdDq0jRUZhe
NlAY0bZbyfjiv/AVkmySShlvItN8QPGo8X+DSgox0yLkvkRtL+YmxHnZbRhZUVZX2Gb164exyMfg
1Earcj6RCzCXvxQbXNuixcmfByf/+mZ8PqGg7nd9AFynPQRu0hJPw32JsW/uRex3U6KUMw382zy2
xNCB9I/95iZAl71aaL+DO8FKZwoqWTByP++GmIqvB/8rHFiL06y3ebAaS6HgOcfJcPkuTw3k49gO
UOD24o8syH9ODCGeHXwNRQuX2cC1Ha9psJnlEZtg6LOQCRkX1ZmXQUesBI6jT+i3vDrd0Lh2B8tj
dEeSeO6et3cBHkrgrdZAKzi2p+F7hFSEdqyJqJq2xxVfCQCE0BMft7O3N6J3TA4cfAECXf8wxAsk
+pZxe84YIjgOVcKN2xZ6xmdqwR1kMmdMRaDzIuThmpbpdo5aLYCdQynOxt8Ky7QHr/3QuCBIHMsI
iHDLqqzhijuql97yuSGDqKgxUtl3J0pv6e75HhdmQfWxDCM9K6/GQvme2HUVVA5iSR/+oZteRDUS
0EOGGHF1i7Sfp3RlrTBmzlCgr4BdmC7olPWfxg16XGlN7vBVWUpyzwmzdTUiMa+Ft5rjjsMzgyQT
C/CXU/vJ9j+2zPwYTmn8ZwTrC1IgbRxKL22CqAofBP5Gm00trTAwTJXFlIh37EyIbOhaeEutootG
I836myzk9PH9U70mZCBmkD8l9R/Sul2/RpSNHSR5QWN/61lbSLTHf4oNoEUsYluGPsUJSGaBsDfv
9AP5ZNQUaVQJAluRjDGqZ93UIlCnDxnLNCFwPDCMNB5Ji+cf4HqnKniODQXJ9c4Lji5QJirAVtFZ
EmOQ8Pks/pIT+4AmFCTnRLEaNVnj/UU5ANEgeCNyBVLvb66dVJkMIp80ZDyXMhHkfp7usPYrdSX5
X0D8yYVcLh5eYQMhGqrlvS/xcEqJk9xB2vRVwgEusLrQ+VNNOrGkwTuk4np2f3dU/xJYJKSum0nR
hshPVZLPiFAdxo4A/Bpb3Xs5lIfr5BNg2y7YKsyJ+mWusbIMjmvNOlzjdiXY3ACpb2axXZHhh86l
17rR3OPzhqIRjJHGae51t/+++sK3TLtR6eVdV0OwpSnMRQ2Zmucy9Om8fiSMJjOijAsPJJAbT99x
jxj0olHU/4beZBsyxFLjbLzhLqRUHblLj3oYxTLFNlUxLL3SHNrwbJoiIXcUldlV+A2TSGXtXNv9
9qZ9MDdG1vpBY1oPfJvBQctnjGg/mxA127H/ZeDH3BEQG9f9Lu1U3Gikd9HbnJITXrl6ASPJnq/n
Ux7Ty+odBuenZzk7HioMLUJZyPSrIS9SlnH2H5V745wPMSE6RLnVmVgYH81we+NtBuPYBRQfs58f
ggGwS624RSwhqgKxkbiaCm92WcLXHphLAkV4JY1w5H3+BAsz9yCkva7pwUkdWVQX8WjjiIJertUC
S0vwgJ6brnPvA219QgUnk9qxYYztcTuTlYH68J1P0p0kpA8DST4Osd/P0WVsladPEA02rbgjahUv
ON8xRGy4EfD+jcMEIdQHJu17v23B7eosAnqsKzesxarqPsDMVCz0cInviXBvr89R4BTIzQKZCiAX
JYj6UNYZhgcOO8cvXfu2332FhywzPU7fLsWlX/srPJlQyY9H3mk3wFjTmCVE7VDF+hL97NEEGyTe
4XeuLmCLEaZL/zfMhnt6dsc504HhaYThPkgIP9NNIIPiN6PKXbi3jrXbClLgQQkOjGEHalgTNmP9
jPWVsJD5uqQ7ExGgAi1w1aujLVr5rjixHK/MrQaieGd1Ux2d7AQJ/mKXc20TOGrKzf4IkKqC7FRn
fx7r9UI/XXU01lIK4VguCXOuUig789QJPDfLrfQjzR40gRI8UiMx9JGRU0E4RbRQ3JJ6H5D8mnN5
Ibo7BZkne5Wo0FHdsKsR5OwkOzRoxCZBY9E+OFm9CY7TKgEW+RuglflmsNmtNl3WRBPNx9SYwpE8
4uU34JTC1kU8B+sVzAYI5pCF117/gpT4X2HA8xBUynmbloj73peZzF7wAnsCXIOl/wm2S4F8JdRC
c9nP+FZUVMOzXOizzQCBFYysAnp7cA7A/oiIG5oic0kW6inXIM5rQIeSmgiD7B9uKqRUbKpENDrD
9RxJ2lXr3ru86ND/d0G8RCW5fhbcou8FvZQQh/IBiKFDcNogBcpmEHQbI2sdL+QA5n7bXlexBY05
JaejkWxCkA6EN7YKnrcuIofCPyZilLmxzbavoiW7SQmoull2Vr/8hhicF4vzXnq16LNKJUuermtR
fe2dYWk0Ayk/5is+DyOKA16P0bWPxEPFlfyxTcjqz/e4AmOrF/HCcse8Phw8o/LFnQ3GspiQeo7l
rizGSURo233lBRrUOTKEPJwl+ObUl9xZ3aOS2gL8EqzzRYkyjTSjte2/CuUDbbey9+k7LD5/esuh
Fj68EyGMVT/vlCkVgd4sY7MdkzQpl0syvfZCyFJoFntgdAg2gnoRIHSymVcaCzWQw3rcYGIYHAWe
H0JPOO9ewvJEzROL7ZF8ZyzCj8MIgmauo1rbBpQ0ZumbcDJhiLytyTtTqr2P4RN0SJsfSTciPQR/
S5heONF4kUJ5k5d6v+gx/I8etWxov5taS+eHfPP7INQDlKk7RXH3o6/p0q5RMhW882HOgrC+Kkpf
D8LazVUb6N0SYaiJpO0SPtBDuj/C5K8VlQnuivTiyciN0z9Reic3aqu4FYHnS5wBZTkVCQsf0q+I
pg6Yqmd9i60N9U54cxdHIn5Pn36ppWA3qy8qk5VmS7LYO4fzzkwIIq7fZPy1iSU27dFqv2SSGxB/
8gPEyCPbQi80l0Aj4vuL7cRXaUd3n3H7XIc3WoZIFeLtJ54FdHQ+VSTUs1tXJlZOKmBQTjiAEE6t
e3e4IijX+DomSKUPEbxXW4jvu+uhpEhx47ZkCu3k9C9xlOK+AYlxfmQ0Ebb1CmiRknf/2G1TruwW
J5iKmEWxa7UIgwB6D2VdNtDi50wh1EkuO28RFMxp11cb6lXpS6RinglSVfIPm8TgkziiLWExoZP+
vm6d8AJ/J8Pjxkg7NNZVJ/xF+ywvrrUHpRSjtBFtTkl1cf1pe32aP3XwuGD4kfj3WPtrdhkjENtb
i+2BRx/o2k/6lezr3RESVPWvvhHU+vcHeK9gpwYWr3cIj7nT52i+EBTVTFmfqU8gv2d95SKpz64/
Kcc3jstVEVkyT2VJz0HlQBTHHsQiQEd/o9790zQOFDw4x5xCWtgBQgWZ139ZdheD5Cs5/QHNWKau
9x5Sr/DtI8oaRMGUV+LoxA37RiGgL8/WGWoMgqIF60SyU8+R5D+bvXqtxcVTxknyG3/BAazmuC1X
kWT4TLvUdIOw6E7WhTwaCSiGA5NCiXClWp7GAd47oF7L5JGFslMhB+syoFMBOg58Hm3k/5Ly4X9I
o225PEUyVUGHNb2O+QT5YgR7zlknMsSO5Ruv99Tv2PiEFsN0W4ysoWrDaowmHPVHz+Bj+QRsJG9M
69vlcS/TwjC/1JmYgnUnD9sENO0XN0tz5tBeM6xwh5iUpGGsRzDCv+zU9YIfYvnK8KSbC7RKX78L
rdbE/SFka7T0Ns8/Tzxi1ZK1jkvAXuA0uu3YUZMsf187KK8CZ2dDUZumA+L5slVIdN7o/KQEvt4j
keyg1nYsH+TmzatKuVjbW1/F7Pbp0Q6YDUbip4xLHzjTN3HRt6HMe6ItPVyRAR6wl1ukgSKwa4vU
j/51YnsPERBqqyoKxhT3UsZNBUEXXoC8m7+Zq8B9Wglp1nXytbrw19pDPDKeMvSgb2ULAV/oBs4v
yzTyWRhToCFtzmEXQsh6ZvS9SpG4SSP4b+7qFLHCLqqogvS4YEuFUbjSB59wxHPSZip71wSojIzI
UZd0Go6WSqWqkjiBJ8BTGDjfuXVJ8rAr/n537fD0kYnieMxuMEXAAHwoqO6dgO7+xFEcrzwpTBq7
1aYCbphzGrnTHZNgPpttDQah1ZxqIdvUzbzCZyE4TZ3dEqoXIVXFNVjtwWgzoHJ8NYL1bJAxyVZ6
Lt3SzXn15l+3Ep5LWN6cd0XNVzXLxYPEhU8m1eUrSaR1S0dFR6ysG0Xqbw/CMnbDBnqfRaFwAaqN
kmpY2ackNqxEgwTFocY9vCOTS6DfTWCDntCYELh39qg2qcvbTuwGVgUTgYOoKIyXSOWYM9B0ytf/
17/E/rKfsbG976UPXM04BLml4G/CtfIFop9AycP/XBU8n6lpfYQmVMEaywGZi+DlVBUJCRd6RSdG
8FxTcdNZcTNpB7YkWHg99tK9sk8EAE/1CxDbDmng0LFSX1pF7b86OyVSvRADWYT09oloiyLOPFN6
IWkyhG7l6KGriYne9gjdMigD1AE7e43VlBek7v5/Z1HYgkI832FoCaLIkNVcWndvFDdxb56yJUu3
xbGCPyyq75zbGMIsgo0pEUALyP+EUBqkrtASLqHjmXKS7TUizRu7aTQC++Y9/tN2oGa6jsew1wt1
mCH0a1PvS7LVplHBf/25q4K4D2IMySnpE+wajel8ZN+n1NZBspf9srxKKD15pSFP3nQtj8kkHSM6
7Wv4QEC2tkLRDYKU+zFkVVsETQJtDDtLbobhelnYBrAkG/zItkrb7sgsLmEJZtmzD0jRQgfAaK0J
h0R6W3rLsrCzkqDU5Idj4z2XVZW1jDRLhWTR5hV/ZuPlYJx33Mj1x/zXLCHzcBRiPye3vgGtC8js
jTKL0js/zYmCmHCLnHtmEzkifS7Pb8nT0kcMJPKw4HiYLrNJRDPnmK3LJ9/NqOtTRPB6AvNUKtRd
8AszK96VgfRCVOQB8I5tGfWSdt7UBe1KYFEHGTJYfKsvBI+87Qsxc6/a0GaF56p5YfcB0/Fg87hb
T4GwgylbLlc7yUaZTfbBmMhWwUBThJ6RJEFf35M4aKcN4ovEKgwDSf/5BSRLuCRZT1CDHudVOB/0
qIOwVa6rRm/Zomj/5eRdUwSivdBSp0fM19wEbAl2Q7muzSCpeBd0zL8td3VNO1fDfkzrdsqNFavX
sOMVyU+/mJEvuFaAp2X7qkRRd4U1btz+AszvAclRtJA8mzFHAHqCBOHouJh5Bo5NVpCcdxuU7rZi
O3sWrfBwCgrX5wfcd2J3yEN+j1zYlFdeELqlc40j4MTV/qbCPvPlyxU9ONLpyphat7YwFyBNZuob
FFMH2A6rHs+bz17FN9hCIUxOgdBz6Gzle4BNlHfHJX/cpHaNDDcfEIaCYKUbvkXizwMrbmB4Y9Ec
cttxi5KlcBCcXNLJSv2GnCf+AFn1jFaswLzLRqiffjHd25Unle7vvk7Paow/2D9I2zDKcVPkAsXr
240+BIigcMyMZexTKJtO8Dtn0fCZcU/pOKoz4YtNVS5c1IxScEds7Clgrg0540t21vTbRorhQQBk
d/EhR/yxfXtf7XT9ARBSruLnys4vDhsB2mCnVv0ZLqzUuVLPdLkTh4QcEvAGKwRd8BbNdPFEOk1r
YUZFRxtUW4xxIruUnIKXHGoNJxl5F0hHwX7wCY2b5CnaxXRjZy+M/QXqkpTAbRqi0TDNqI0+K6ND
Yoz7oz3VcLWD4+fgM0IGy8OtR0096NWie2M3Og+DZveDHtYfA9nx0LmUpFIeVD8bWd2qTvFwXdyh
ZSrNg9rzV2MgSimXtGmhpWgd3E77+w6YyNWc4P+bSYEFs7NcDr9y1tnvFEXzGHnP0aCzxCxeQRT9
hmHyT9FKAhLMd+uVps1Ly6dJZRk/BwpQjfukeYgK1zhmbzinYm0xozS3Ns92G7Srkl0RhXLHfVSB
qzUlDcPW+ne/FK6gJkBbhOnjhbW5EHc7SvTLWJZvEeYP1XekyZOUpH1Y/kWe+ep+rC3hDHwQpnHK
NzxgzSnP1CvNkUrvqmLvg1n5vjtW4dQUXA/McRd2qM0t2PVYF6KVYC56OBCZ5h12Q4JXtNLIvtpd
p10NPgy31N/ZuDGv1GE0SMli0bn3BJuzmM0KZRVO91JxUtuwvnl661VMqDuCDtdIUrwaZ38xWBsg
MF8852Uo1QZ3Am+3768wIeoMerzf/AIXunFW6vM0Ql866XNMtYONCj9NpH1VANtCPg7Lb7gZfE5w
+tb3OahEa6i3L7nqSXzxoOmSkAG4Y1lVsxkgakwpYqfXnkdbzm5UNFvKYxGIkdJQL1KrwidQqRsr
BbC/WFOKkIyxxmM6CaD4GLQDZlL+bPlxlfYhKlDqwviTrzvstVLQCZnpxldxU/ATlwUm3sqMByp/
qN6Z9kdG3hFzJPAUmVl3njnvpa9/vY3MVNX2awM1uPMDKSlRWOb1m6qUf7879BVYgsUgYdhQ0LAu
EkKJByI7Kt6a+YofKfhZIv0YY8RBeHc2766/dp2FcxmyxB12e+bp+H9lKZcto7FTbalxAn+CmNmd
yaQkSFJg0dGHuXvTRVDq3y+Rk/VjizhWxLM5uS1KtiFxwzyAv0k5Z4p9pPVCzrJhs62qqs9IUM2/
ByCOhs3Mgo4azs4Lp3nyedwx8E50Ay/lwcffrim2+Qe0spr5ZiNmImguZ2ZXJkQLSlxLowy8motg
AHIbY7f686SQM2iG8LfliOCGRIERKulj+VGSvt10OYnMoM0gblIQ+A1KOBIobJ/XAIdwEqSODb3e
ppzYW2pR3tEBua2avWjGUFEFqhQBLsQ8PImbTMikFprfgCpYkgus99lz1fToR6DB/5OE8lTFxoXy
SqlnTZ0Ql8Ogo7UYrIy2r+0xkJIUuHJp1ZVKzsVQHyCAA3UPJZZQ+EhyQ1T3YfZv7m0sKUpRjAIU
Ll7/L1gBLfG88jDLPXu4AF0w85Bd4os5kjKg90PTRGr0qiS0S4ZpS9CwFRnn/NSgNz7QXu4ZVR8S
R6zx2JLvH36RA/rpRPLy8HCHy6Q73MkcTraM1pbrdL+NhkTyJYwh+DClonXn5xRXqf9ZWL5LFRB9
Fsbg49h6qBBhWwmI3F43dIeKPpj65yimb6GPmCHId6c/mHF4p1b9TywiudXvOcn+UeoItBNUHwGP
Sj5b0cwz4LqEqjlXEmwq3gRXxt47lAIB5PGvGa+Xvs6E3W654vAQaa37+qQphsjYlHadyBXaVPcH
7rDNDjPJG5rdTRb+tiXJpNJfu1Q1oXrs7Rr8aDy3Y8nU80V5dv8K7v5WOPpuW2rHbSVYa2ufdsZo
B2ijAaljCArjJv7OvZoslwObN3HtHK1hWgFLd9+RihXFi0sgu6lLQwKnisQNiuJim4lMbsgaC+/Q
snBGMPlzh8mpvuThASnTM5WbrZC8PZk+FCgLHz+4k/xj712iF6Alh21DCTwgd/TINe/jsnKwaEAT
2WsYBm835VuGGB+UCluuHFtefuk3yO5XU9/8IKWG6AiRuPf4Cz3RpIM0g1+c/ggGDkeL5i5wH3YC
9yQNzOSBWdvzUuZ8b417kw2YauBqY1bmiKYcvDpywPbdinwRWq5w+dfYs369hNYy9gQGEMcxKPIB
PpLieKaALPdx9w8cirTmxzKr1AdjxMlxnZalHLi6RWB4vwzJcmwTtbhmXuWBCMiX1wzFbKlt3RCM
TSKOei44KBS1yVUVjYzuATjSsTRPjS6R1T0vb1NOUq8xENXV5J6X4w5pyNBlOB65Xw5onHDD+tLA
PtNDvXh4dY1gSg/ybTyumCgya3nsd3xhAdF2l7JwqkN+iDcKay5kyEX+PeIuAnq3MovTMhzc9akQ
dw+kRPqOb7OrbU6LFCCX4cK49VVuy5TvdlPvCwothxBRuiGeUY4QyN2EDmL7p/ZE48p4uVqXfmz2
pUnzTdX7yYwTreEuWbNd28NiYbwG1O+5/Xp/ZE4SOf0npQQBjpK+kxx9KcifaT4ufaD3w82ws8l0
ekACyI/NCP8piFrKjY1VgzrHfQrqU44ETOeweMHSagkly5hEYUNnKqcYRSERVARhAzhAE+EpP4ro
p/SC3uE2gIPKuCMc/W50u97qeW8wNZX2hWdCEqugxU04FTZocg7ydFGMIp+QkVCR881IL9u3Yi1w
aZxFS29l6zXI7TYIvx1BLETZ9Y3Mg5P3jUlJOVCrrTEoN1biF0E8ZgPhAvOEQ00Go8mjw9Be/n/Q
jmXW13rQSM8oGKLkeXmlOwgxix1upqrAPP7DUm77k3R6guvsOykxwV4hiVXPV5bGJAW5e/kh9GBF
wjo30dDqNxg/YU+NteIqew4bozLapmg0W3kW6IwiHABAaQAvgnjeKlsKCQMVgcnP0hvXp88nRTGU
QpVaqsncOyylc+hlGkTfPNSwC0LK0pXvsPw5f1VZvzrLYi/UsHDm1/oh4HYmA94wqgxMFHWHQUSv
WJBM2Zpl+yc+3edNZjXCUqa06z6AD03EoSbjKBNjqwIHzqzs/l6meH+8OrjyyXuiQvEzwJo1T2nJ
tCsjgiYcC3OKCyAkxLJpwqzra5mRsAGt8qPO7oNhZdDN02PfOPyFx82f+RrhG4HGbRYV5KxUFhGj
tWtKLBMflorZ4tfJRk/AqCx11zQOZfxNGuqSQEXaadf4UqRjAGNwksd8MFCw65qz6yzzBxvXyswX
KmZ2DqasLB++sWoMvwzQ5Ek9Km6RwHU/klNvjnCWUHq+NVtsAGNEdOWPQvnO19YO2moAXH/7gKnW
QBtkD8QdoWalIvv0QCN6D7wChwLA63pE0PqVITRiHOp22V5IH4B0ZT4EsAk3uJcsxYIYGoJ4+E+r
eYGTdD5pGVPflUiF+cn+EL7ubgDmd9JrR8KfEr/KiOeKgq6wo7of6j8n/XRYmaJVm7Nr3aqXZBsn
87xyhxUQHpjGZLwqMp5Q2OOZbt+XEs3tcJyw8VU5cbL9W6ZkqEeVyi0j43bQZ3zdUTSiW48YJfuA
g7HR3Ln9eRmopUS5O6klH0yYlSDgcb6IDC/x6+VtgUPHba7j8pfUrGC09S3wtNueGNMcl1FFvsyc
V6ulnYf1H81df5TVVGn/OL8FnYzXAEqvagdpAjuW5PCgDgHug1HBVfS71ufqkxaFexJAphQO4Cdz
sia/N7xGkjsyLrqhkPZvQd4/FugFb3AdgJCZjrAUnYROZeeDZPpnHuiJWvKZ3tH8wakIPi7mxJiZ
q923zl+ipQQxrt1fy5EwXk/EQSLlRaAHMJxukZRrpJsljE1mPTwfLDA7mSRGb+ncueRcRdP92KAB
3NeDnaEXsVpJqKAwu76JyEgw4te2OzrNxZJTQaciHnZf7FrcF/J/huZKX1g1sdf2pXyb4oKBqQwn
z3L/y5GNEv8ObC+PZiucSMmS2faofliAsJl6D3QygOOL7zoSJywLq2o3rJ6xzT8RyVH4+SZs3W3K
0bVXsuikQfuQ8F3RZTOTbyHiAH7GzsRc/hMpnHuOB0lQ3b5ESe2h3H9ucxn/eMxs0iAZXd7fibQR
5Rau2iN83AgH8owM7i+qNy/km4fZ5whjRY57tPrgpWj9AeN4m9XBvsc97c4yMIOl2Bt0BTTadje5
eXxAKb5XpmlMbkH2z3ucc31aKyY6GbfebttG5KWSU83nzUiP4jdpNB02852gih6Z8vqSJILSUqpW
WLEztosNxTtpbh0UwM6rMpDOQKGFo5QPUTxi355omq8Iur3tdEg8+4AdTLFvO038N8Z8u2ub6pzF
Uc+AvkNJ7SHHNV9Hp13f1QtqWxtWL1qC3yyt+cIPtNTNwLQgn1PwsDXMJ1UvoGInjOQxyG2sYHxm
GyW5wYX/eJa6Nh/V1mOUux4SRZUwM8V21tMqxx0Tmn5CgpgSXwI+cS+B9Eq/mVwjtin1Gnqjj2CF
Cr2T++tP/MLeQhy9jGsDJfcXPhuHSFSWSwdqPtAU6NdnjTOoojEanFOkEYKW2UAfCGJjCgrR6bWL
wsYc8r2EOwL4eVq+zmt5hHJLo0t0MPaEuPKiFOGHoWGwFpb7HHlI7tL+n61+qJlIgbrfkYvraHwf
J7Li2f83hXHk8h/lT01hkdDc8Eo+XLfnMvDx2S+5plOKrZMEFT2mzdYZ/EFpmOypDRIXsLFKGdRl
xddnpBWvNr8+cky+6ZpPUIF4tDkWpMSmAIyxt0kYUXmJ3IOkawZWjz6e5ry8jLYve0BXS2R/UMTv
WT7AeTEpjpbQXdiX1t2zw3DyfaZigBZA4LaPSXfEBs4mReVOLS7e+oPGGLoVerfC+RYRhwTmJL/P
0O3jDA+Sv6LEi2zN0W7h4GBE9BOYQ5BwtUXHfKQVG4nhtTAxnCryRP6uWYXHadZXtsAR+Lc7c+6g
Kt9DUuzM8yH8JxHVZ8PCDyI6/zaDmebnY5nl83DrjXBQELCgjjnvELTrjV4uIdFTjlAne3ukBf0T
tOU4VA0By7OFqLhfAeDMz5Uaj05DrK/2bfdpX0Wsrt0i843mONHXxGpkTel0FZVrZWCVTL4N0L/Q
pt+BiZVPrnrwpY4mldy6EiXTQZHhdpKt658uxyzILgx6ewXUp/T8aBSwVi8r5rmnwsiPJ94U5oC/
pwJV73wE4/agS549ugWZ5fWFDDLHoYn9VETIvaOGA2Wu0vcSWuEFXDJzO08YXqat7L2HNvX90Odx
UcW2jwk3kDmsUJiGqdI4VIUgns4ItCdHkQmi7byDoghD5oGhMwclnRo3eRIUb1fSCaOMQ301Oo91
3uRjoJpTECLadYUyQWIpbLhEYwhjSogi3sc1/V8fhAbSK7+eoN/oo5S0w/90+Bb56M4eMbhnccmx
QY0Vrs0u1e4ftHjnHxRcz1bLGRF88L2EsOYTGiiL+F3/0bGT9E8s3f1N29yhlOrsdfRjlJ+FqfSp
1dPoKxDVH5Lb8POCpRYY5lNcUql5KSSjMzI+TSFCgAW7KKDxSnOmWlSExJH0w5l3QSHsjDt9smDR
inmmPB6asmDd1vdhW5c6qJJ5f0K/Z47IRTFYzz4YX+tt8cp9FMNHAU/YoBXeIYBdLYX82T3aQl5K
39XMRFcVI1wqLiMMYdmep1H+BmU1abpK8l4H2GVrPHsbsXloL7BWh96zbug8k0n+lu88ON+HRuoj
x4qXtijDYWYOcfma0qnM1VqkPpAxmgLaseDclF6Q2obVEVIth/rSeE/xeUPJ5TfjZyGg7wzFUoW1
ZWvs6wx8O7M6WQaIdl2kInjyqydXPn6fATBfHfI/rHIHkorShs7Os2DrFG0Yy1L30npe4dCd/wgm
eLAjvU3RNRKCK26qRrIkzSOdgC9BdKWidNByWJVlxsHBybjPSGH2czDkLhc1whoawP6ELHufhK8t
F2oqbDuF5yjEMhjWkpFr8igWYo7I6/fbIopwNcyhh6cne/IifWNi0hcYsnYBiT3CmNkZL+QjzvCf
dTCqZMDIfAKoEyKeP2mo4eY8GICIhDfuR4ibFAwhirSotU/SXOVG8BRnTLNvei2JMwMfBwPRQLR1
cIaweMbjkuZzpY9lAgIIDfN5N2zx83vLYhXEoOBkOUg+tzT6fIUPSTLL1lEaMWUaTXjqyRa6D27b
ppJj2Olsb5KN8a60fjDqvn5TkaZZdmn6e5a2hgiWkpRoGg6KfFGDsr9QAZ8NtKbFytdqZtlqqkR4
425UH5/vXu7sKQb4snvuOETUXUt5L2go5TjuchEG05CPjW7aDRWn2ebmw1MzMB3NroMrqSZse8U7
x2iZl2Xa6kIyaqTvmnUG0lwFYM8Sk98pog7ti0tM3qaH2fdmeZu/qO4uRgcWOTg66sLRRP6gt/J9
NTHppCeMH9fuC5d0UaUBWppOGpq42IFiJRFrdQ6zGCT1gCi6S7pHhzsvlthf0Ile5YWCWnKWPRg/
YbUs5vI5mnMCgWmHkQiRlvHOeg0lX4HAn5B7B+eBkBNlTcoZwOPpYm3QcY73cPpUidv7uUHjBR+c
1ImBrKnyw5W8r6oEqJYH0YXWNKuE9tlCNR3dHNG2OAkRDH9O9beaDA8lJeCHMpiPnvfkmZev1Ip+
eaBVeq5j1smtIQtFPPCveqJuAMD9Tp3AdEYc3iY6U32dx0lIEQ+GZ1mXmhEn2Zf7ZzmpEyFFtVOJ
cOxbxsh2NAghg7HhsCF3eNcMQMsgecvEJKlMvJFTi/BoVveVmZyl+jCB9rFtgsOz9liEo+55Rtvz
uwEVTY1EC4ZT7QF/C8OiNKAIyTW8H8+guN0AGJXM9/ea09rtBOKOY7TP3gNfupRrr41PMSqgpDjh
L4bQCCvNwROIWXtAeU7xxwJm4CPrLNFXW5TZZiqYyeLfXBlGgbV7z2rgl0d+OcTtWblUO0xnyF4C
61C/jJagGaLXyOSv387j6n7lFR18UcBa3+OEZAoqVvUveO1jYmldd1Ai75xKnE0uhCT51wdrIGRT
xf2hDcKLHCHaFIKe7nYwnK7Rs8pZdJXyVxUIe4FOb/8XWA8Q/sVpIvVDS6XISPRM9Nerxe0Gv78A
HFDHXcTYXu250Rfs0evB/wBeQ2x4y7MPLMb1PInEh6GGcdrb9gsvR+EZywLGcWMcPdvYOF/MgEmb
0qI6WyqG1mmAywyDQ/yneh8kkpB4OW0gyzziT/ExZvV8hW6FEIFRnB+3Q+rakFMrBpc2CkCjVWfd
u4k1Z9fKxdz6fq73lEgfq9lZtYjjTPxSedOs/E+0eP+gbhwbIg6XwjBvWMtJ8p7rVyhHEvjn/ah7
orSmVmM5kuuO+qahg7xVTMMhSRzRB6DlHO6l6XIGC22TPDM2H9/k2uyPWaTs/+bJ1bHXbm6VZ+67
dgHW7fu2eQUBy7sHQH4NaR+sYusJJB+pUNIDIVbjgKvP16pRkn0rpYzjJAbBf65iIGbKBm3gB6hE
J7W2PQFFmJPflAk1S5C4n/Tv+YAQCR6xi//k+Y+EcGuYg1QTxrqNQs1xY+dpY6hofCaV43LUAgSs
MQYWxa9BGWJEzF003RiAG7xHXifXHfnQdby6Gf7ExDFViMWlh7PVTn1G9a+fJ7iE0+a6DkK33kaG
qDlkFWqbZYfn7HrpRGMzoKqUJQ1qzjmd40RR7VApC11Vu7B8YHTOX+ICb7AIU2MMAdJC+ftprL4f
Bu08zx4xL+TBRtOUdi8vwy3W6GhgYP+jsi1QX+u28NQZ9T4+4sGOXDkc+ZgcS1i7Y6YEFtxFdfZV
MwxpJzRyq6nrjEx7JvDU7kaEXzM0OKlIUYc7sH73/jMy37bAz1msn9VKNGg/z0+hQ4ssn31yoRHX
pAlvPyLcomIYUoCkt3V0ov5o+aeYFPRYwaRN+GC3IBmKlgqmelmkqVxaGF+FmByACFpDgrn5+lRM
oKN2xhDiqUj08FYubW9x6rg0Rtypf8P7SdyqMmgfyzngCRbPgYFnmnLxzQDtFRtB33IHQ6hdzSAv
rYYHTzz2/CDWJTavfNu40bulGZck+QD8gxfdsgRpVvDJxgMGuhOxTFalwG+K0FwP/s7L/s/cdznY
x96SbQv11hOJzVFdiL2upQ4kRuLe1m9dZyssDDmwHx8UVs2kiDSert8bs+bvU6HuLd31D1oJWCVd
BweW5WiBGDBpudlP8ceGqev4p4M2tW2KOgyfPcxF5XYUGpg1msl0Rk9RHroncy3n6+kKqBNCcXK7
XSkd7du7rsNsbAGIoyaEP9WPcuKrCHfOzLytm/BdTRhMYdEZ1k84TaMEPqxQoKxmBEKoh+qjiwcC
AGucbXwaIM02b/o7lf9oQnm90gtMo28wv0qf6oQgomusenQtgqXvU3X6BrZKzJkLviEnvlPgWprt
X9lWRg62U2YKJ18cWHQzVIyfEuXS7In1iYJk2nIm00Ib+9/C/NQjH55q9e+snnXNxA/4BR1VnBVR
USFS3X+VX+wEi17Z5+duXZaNHeTk2w+i0Me5utclfC9p88dlTL55V8rCryYZbYX7LI+2rSvZXRvB
kDyjIrFwzzzxeZxTm6EWmP5gSbgpB1lLsp2DTElmaGYl06qiDz2P/w8qPNA7i2BOtpXHk0+anhr8
IVu3/DKV9/E6rZI8QVyW0cXwvZC9HqZVmwPlxnQeMkHQTiyRG8V609kP+X6VfyTWjrAugj9uEenN
H93u+Wp+s7xGli1hjv+LYEcepYdlECH/9MTv93ZdCNTFjgohSaPC0Mtg8m+Nrrr5FfUkk2L0pTa7
8gT6UZSwqluxDBEhIz4+XMjuHZXKNY7PeV+6+0uej2SVO8X9AYGWVCZ4BadQG3SWCW8bMDX6vIzP
A/c4/If68dx69FncVh7hP/elB8Par3YBzcxXLfJfh2gzb+YWXrD8pckG2jQkzwN/YvYFw+UtqX4+
tfVImxsjH3RmAf4EsW43cnUdyuDC9F1DzGllGN4YifYgs49t/uhwvFjpMGeeMVhSEtmtiErBlbwE
UWh78p9Pv8PwA7ZhbmTOVqAgwzmUe5V0/UqD7rnoMY7NWjGBJ3k56HdPrbe+kaJD5D+J5nk2iBBf
Ziu454dzPIv5mudnAhlVABY/rtTnHw62rEyRq0z2fCOQ4uU7D2F9AMS7VvbdgLI3Ew/rKX4fW042
lSugaKowv0W1HPWJPQq0BZLNG9tiCK45eha1kJbL82pBxWD5RQMTVmIuav//+ogJ+8lzd9ZI6XuW
RClZZ3k15MCs29LRdqaS1wadLDl8atCCF5vXU3aSeBjJYqtP72HNcSsg4vNTqoVdw1gzGnOm0LfU
kye3Fk94MpVk/a40dAE08sXpb77hSRjGmubsFgw8VY5HN6V2HuQx1BF4/1rYFDdAOuAMU/vB3mgk
qsYnctEVKCmAPMjxeUjntuOXEKUhW3nX2xmn+x7HBzc1ddFthIKWEhR9b+Q6NxYA3vtDCaD5oaMm
WnPWtRHlJWLwb9spY58Lsfl5SNLhNbl2K5bIGWP3Z/23yXkz+RMeeY/poXjdTtdKWUePTnr2JPYF
+E9eRpSQVkjaZCrNgzVhepPpN2Q/ymaXhAsn2Mx7t9fZ90yI1qvBx7Z8bK6W6VT3/Wkrqlfoqsm1
Gmfc2bzRjb0jSr2Ho5E8QN2lwS2eouYwjErEHwWvFNO3ON6/IuxzYaV2QfsHDBM7v4lORu6bIw/l
LGTVRUm5wNxkSpvJCgxr/wcuSFlfoxde1UdltI/v9K6eohYcUTM2o+xJfe15znhmKkmxWyDpmi2g
82Embdzx2MmKkkH18y28vPMmALBb91jMirAg4QjSRyTcvmg19X0ty2R7UZn7k54XSfiq1m3Rl/WJ
yiTwPifYC8rYswgShQNsUhsfNZ0ZQtbnKE0U1qnqh+p7q/Brd4d8XqNJm8ORxDwy7xj+OfjpIlES
UYRXLBu7/M5TMjvyi91f33CA/0qYKfN5VTIjSu7ubFVebm4oOIa9YKbJIfmehzhCSlOyokuhoiZn
NiHpGGGa96RAl5ocAQ6Q+kJJFgmIdwayvgrmbWeBoY2eAf/kMX5xFKK5A3TcU2I6Qg3blC8lhEZJ
HT8mqKTvyQA3bHVDndLIFad5+gtUEZoxMCBxYLtbbMpFqiSy73QDFxsSFuzWze7cvAtBmohtLuO8
rYFrGQ1VdfXug8tgdWkNv3Ggyt/DlmybsJ3vSIAXFJC56+DjHo7WnbAP/uDtTjKG5PAwxHh9zGzE
jkEZp2+SMcvPncLhZnQssrXamR04FpD0cvfElSlGiMOduYslnlViLcgg0sgdxmCYCfGGyr48ejmu
j2TTfDskiEdox4oqlOdCPxR1xfDQ/dyVwct1qLM9GP2etd414B8pQxscZ9XmJD3tf5J0S+R/Q8GW
OJFOU0wQZVo5QDSkrBJLldgbR8lWm2z9Mg+VFIr04sGYcYMJP55+RrJzw2a0RISD7Z8PDKiA7p5S
xFj1etTUoLooRTBKeSOmuc9X2O1CMnBvJqOnejW9pMWMxwiEdWx0KLOIz5eaeTELguL9fTpvwg9g
BB1Pl0RYl4hc7RhJgiPegfPquPcLoj+jBcD894JHya7R5Fg3Ivisaj4u2T94NjRgim1s3Wl0gEJc
JoanJ2VPfPaqFQ5GN/aG7t66yAjH1hHF2wkNDSzt/Cd2F9NZVVJiLDXAhv+e4si+P1aGOV7y2GKL
H/EjURVUxo94lrCU/DKL4qUqWit1EoKiDvY8eyE6/1G5y4ZpCXcO2NR0Fs1a8VD8rqIq2m9XocgQ
5fop+pLuCEZrgglaey4hny7KO5wc7MZ8DslV/BPhjCHItRHDQYoxUeEXeh3Pjud47pTzE38qFpv3
9T8y9Fqz/ML2NpeGjKltDkQNwEg4sS3IGAT6qkO2HSKm/BwyiqADVsB6nrdbVzcubIMi/hmchQJy
3MspHgFsokfOFECex5DNOqaYTDSa7eL7a/xtAvgZTj/tHzzqRkpx7EeV/bydh7KyZzLn5lKkgmc+
Z9VFc/46ZxcCgDpg4N9iCk0gqnXdgz9VQxbVvq92UULCvqAob0wsEkYL7C0F1sa3HNbm0e40RO/A
f7ITBiJCVsuSm1LfQDlig5+zAc6Uoy0SeBIpii37jy82IWbeA8KjkI9QZAaArccJejXg3GI7Up7c
kEDX03LypYTEB65FJvmHVMIk7UCWj6DMxL7CTx75rf7ie7tsGSiq7rI0UxJoOz2eUELQBrAIrGGq
hQDg41rqQbu8vM6CGcnIU7woy/RV5HCuy076bRYOicbvYOYyQYnw3XoYLUXDJySdTWaEHH9n0RD6
Gyh+eokINvBEGxw2bFZsOyiqDKsydTzMTrDVvL2hOirEfhVwJjACdCoDUqjsho80wsZDF69pyV47
1YftvaD45fj4/tkZLMU+amMD4hztnByO40tWR1+O1nBq6jfdjO/oYyFl93Rf15G37FbPdcN187tt
W/tso3YKeKbOz2tOvXihy0xPB/uy08ElDwD6iu+gr/54C+IFlBhvKOVqAGW5d9zRWIChFxzoJe9S
5n/5AoMGRWrgeAOs2ckVxQJpgrZJiPV1e1L63f7XRwtzDEsYDb11MFzCUVUGsOhOOgk289ZxGz+k
hgSpiG1WHgFcoCfsynhZ4i5BsBVUHauFdku5BViPCiVRCJM8+of7SNOZynKPbMGyDIJZrVtBTWzs
xeS280x22QAgD2jk2O0+H9o00APpVb+9VpFkygvyqr5cZWFLOnJypmUsQiLzbzyUh5nq2NFe0qUp
w0LQibZigybRScYQscRUeERI53s8GoIXexE4SAf6Zx11NGHQ8akA2txgcpgB8l1ZcgRQeLYHzUAa
wAqQmayT4awbQzAWbUFSVwf2b6WOauhjSUiU0iNZvCeMUGzt6yayhmV/PTGkqRjZAZ53edREq4Uc
dcXlykD1RfXUnmG6JSAximyIihcfsN5KYSbI7rDG4T/yjCOQ4LEPKkUGsW9kEET+J6m6v+hfR51q
0ESvEDWdBlB84HaV19FdCy0AJcS5HQA8Lhk7VjcA/61/PkMSdXqZDRH6kaEN6ju4sgfoEOSJ5Vjw
+3EMcQsCa2NZXgqgp3lfwU/Rh4OrnW7iD4Zmfk7xA4TE/dML3TuVDhkM5VXXvXjtaj2l3Jgnc60/
IS5Nr8xDgyJ3JqchIo5MkMws49S1KVoJzJ3CVKBzxe3i+VCYY7zE7b48EVn4lZD3BlQv/ftgIkih
yl0ii0M6JIP6aFa/W7MzZ3rJx7/t8O1vkTZIJrBvwo8yVILegKr5v47JvZCF2AfMGuG9iScLzUNP
BiFOBK9HVCdskilO3zhXJCi9Ovl2jUFxS0vl1sR8Xs9zDf28VmWukJVkXlQfBRAjocL3rEyMcPna
Ts8RKybMj25J/iZUADByhkw/otmLq3z6ODAn1CNtNL9PrzViCRs/TMR3wmeWz4y55NTR+Gw2JAWt
bRPglzpZBt+VXSl1hB0wVSn1BFQcSlCAWXaXR/RZ8ngOIlSCvOhfvdR6xzfZc5I5qpxS8eottoL6
KCcqDtu86CimzWRZ9rdCmkrBNk/6g4CA9u9wCBu3AXlGUoxNqRE7yRTLGyJzSm18dYVDxCxNocec
B/rnWVb1wdnqv7tDO7XWDNuVNtkZr990upj/9VKBE6cQG4IxqtnTcWbTFubIx7cIGntgUBi6hBwH
6SZw4OJHhJK+FnfbgEogf3vHlJoV4FUU33gs74Ajzy0Ts0xS+tjDipnpMzlSnV6My9CzHyQBi88y
W71weBi6t+rHbzvgsYJouRiDdQJ6nAs24K0dvs85L77nrUi743TZXrIUGRn9MXApDfBYMvSc9Sxa
8w7f+LJQm+phwawo90C0SsL0QdIlElIyOCpHwHq7gmVgzZEbbviTZdZfX+ia6CeTqJ5/AYuyg2NW
3nggfGwJdFQncCO3i5h+VlpLhsD/J7NZjHxK6C0S+RzzSrcG8GjM/di8G9upn8RY3T0NnuD6PCP5
lOMozZKECdzSYdZjKR4s+6ACVcY8GTilk4rHiZDNCj6m/JWbvexG4bncEnb2YHGaC+6SGhVI1cXE
y0pVi2t1yMfY+TYOgrErShRCARTpadSEPlEuP4JYb93cz31SZw+O8ImJvNwIoKvhoAN7KGdCBfIT
zF3tgs3J/oEaCvMDtRV5+qqTvZUCrwYlbS27uzghACBc+QuIgRs5o2x49f8SCP8NZYg08V/KfqZ4
osyWfVdwYVN9P2UAJkE/KkSgoV7j8JllOwtyzzX03EjuN0CsnLJDkc30JTURqUIwtEK+0kJhnJOz
GcV0+PVF4TS9cJtuv6kZ6Yu3oewq8cOoZpj/JO112ZnaOg8EcvCaJ/ucFbbASdnLvnnS/A3HWMCe
MwUCGEo8M4rHT3IlrWmf1/P62D6nhluj9GK8n+DrO8h6kntX9ZHOFFps0hrfQsXMxhqaeJLwUHMC
Ekx3ArbTxnGZj0hW5xaiEd4NrklWIeZY5qbrIUF7UAIz7/uPLfZTaCqxTyK3d+daunW/oBa+oT8a
NEti8D9Sfb+XB4j3k68Ppet9DZzqJy0iUdyr5P2hJEWbk/TV0M7xrA8xLTiFT2Ae7yAnsAxCXcL/
7j2p886sXSudZDDzQYu8qbTK7L6jEODzGMPJ51zUA0zbrJGEaUbt/MIwbhHfClBP2tMNYonz4lrf
FdhfCSQ20fJt+RsXKIzr3seNDx9ccM9eTSHt8M/BIdMIXwxRaePQmMaDdo0YJT796VbSIwPQ6eTn
aXSJkZENYZ8acK9q7OhLPe/QZB+YAhPgq//tCzxJV6cVopZOe3bpWK++W109gGRobWKhkEY1g/fu
aPSR1OKflDpUm55Wbzwm+r9d42YiRzKBidX5SXoJH6OcJ41aDQWGel+X9K805KcLA+CfTDhiuM2g
OwNnzyFgBiwKYL2xbGUGvzxTV2TQAXb3FR2sI9yIVZBOhrAue7uXc8yry7USE8gt2opJJPAjeodg
i4L9Upjo4+Ja/7OwzQ3J6O2c3rBTF4m+9KohIsmNlyAaTyYZ1cY28WYkIYVXDgrpmkdht/5EwZi2
4O5U+jOI9EccapITOUpinB3g7guZ9+us6oNgWIRH7ECYV1pmnNg+nZk8rD+tMgrE6I2XZcB6+ATT
pInxRKEdkBzJUBYgmtl3kq3kEA0xC/ZEs+t8ydU++67ssmoLuobp6fBGkIndb34A5nkYpsP9brDY
fazqQ0sCeZbOPxcAADi9vEV8wo16+yn03ri2ipSbbZpSFxWU32nKCvP8glcR8cY2CIeJfwUvK+o1
AeVCLgPtaoqjsgBbWkY/JQsrD6xwEDq6Hxd952D9ceD8Z3ZG96Q/Z7/Wykcy1GcGkIdv60ZMIMmR
gPDX500P6XjthcRJIN2dvAUuP1q3R5w59O6MUYf708VJagZw8XRi/kbQ7FGt3yYWY5tKBUuc7bPY
iN3ZvfVHt71dkcFKqJUxzp61SedU6ocrsdFhYZJYj2U4YhU/1BCmZYkKljHddPpcU/vvU7ivZMb/
almPwcQ7f0wt8f6FkBBG0MKthZXXev76xoZpUPO7FcAGzaPMs8JV3m4slE8ajkX/jR2eTHpOLLUx
6Jfk5SJhZDd/qXe/8Tqnew+YFyguN23BMQFEzfVJllrCuixgyL3bgtOZIJ5DLWYGo7dgmB45YxIL
EdefjIilfLk22Hhjgm4XpuNjWAyzg42ZpnUzBf+FSpLiG85AAbrkmPEY1CHtqO1Gl2RTOVR92554
omD7+NOIdQyULskYDx6fhpOK8AImwhy01bVXlAEWqEjRl0joMuuWG87IpfsQF8se/ce4s4HjLTcq
aPb58kY4dP5uk3lq5gb6FnhSddxSgmis14gX+5KPrRKcuL+TPcjY5lKJbtB2SgvhmaHwCGK7MCTR
xN516VwhnfKxED/T2nLiCpbMlO2WH/NG9wDIPw3VNPbl/n4zROPHNoDvrjJLXiNZcUXclkKHuUNX
3xhk0DxK0jHiWuIGZojfdm3O7a4Ub0s2lZQUDnaSq1VzMY19+br3AoVeQHOtwFfGiC5Kq0VinMrh
GTEuVDzkzXOysF1LM0v9GXBuUdGxexwmqpu6FbtDyfxmuR+tSQzIzWt1YK+zDUh7LJOI8lpNxbsb
z3kXjsrsfgCo38FkEPGEBpprB8NymW7HrF0Of1czES7N5n7I79c21WkjqWg8PGRtfaQ792rFbiyg
OIEYweFQuXgpGTUatgeEOOAiZkeuo7QPB1rjUhlwHebDDOmkSYOZtEMA/AVuaDu0yaN32C8YIgZJ
zhqggN86tJEt8XwqUiWXbDrAQ8ACZobIn3bvpbRkevaSj+qT2c2wK1G/enac+KQkD1AU62nzlOg3
lbC6VSnzDwCfue4GthKwoD6fDf7Rcx+z3EXQ6nKXxFfzLpZ4ffzNSJjwC0YSaqDiJaWyjd0Nt5+R
gml1czVeJFqG3PX5ynxQFLuR+i6kvQ0pKr3862LvSOhPfZUFmL3de3BuppbyPQrwDji15DXy4RNt
dUIHf4Lc/kIyD1bIEOothr2FC5P2l7maDcm2JXpODO3agU6HSJaxgykLFa8VmdXqI7MpPSSGWOLe
/1yF3VzJdM1HoQnvAqwxdhv2PFjkGQpd86briWJhmHTqfQaDjv6c62rWr2CsNkrX41LE171kBzq8
+RTr/X0JyWWvkxrBHwyd6Q01gqG57H59X8QkhcoTO0C75vX8jhuKeQpiTbYYKu2mr4pixTk7/fBH
tZ4+LwLaokTDy1QxocAT3ku61xGcWzNyXYtV74PfLB0V0Uq4m7M27v3Eq4ac8nM0/+uVT9giZytZ
8fcATBHWfOyKt87LzLawr8RM8qA3mr8LnNTufrWkZbpzWm1TSGyCjkXqx5burVkrDZDVeiMf/e8p
c6oT/RzQWFmWzxlG5U6PSU3DVSXtElGZbxDI85fgVi0JjgxrOgat82TEHeX/V0Z/Yr3qM5bUeIzw
2+izWYzG0GV8eyKUdxDJvw8qXSB5cChbx2uBgyyq5PRpoQUbaEPYRgdTmskVh+xS2oCVJp5J+bIZ
oJZKZyDTidCy4ELa70675qoIV/XmSLitgvv2ih/gjx2X7FYaJzdh6fvDo/vESkTfhkmrddQO2ALR
8hRjSXlWCO5+CXt3PvTw6756zUEhSHxnSrIIrm2kpxSNGvVnQLYo6o8IxN6MJFqWixLLufIina4d
hkkMUEPqOlinYUdzHDqnuSsdr+krg6x8ZhCuXi7xFaI9dhOXqvvTfhPApb/pwd0BgQh+37J4N51F
sJHHgjGPTEnds82EVzugXo3R9ljzYspvyJ+xxScFeMfHW8KZ2+JVvhx7UnMekA+DRS+bsZPaqlXF
//U2GLpuprtpB1POGi2TzIuzKJeBjNss4dl+PAC86FdczT8edHoVwIby+t6+gpME4NjH+GVBPrcf
JhjFEPOFWUOgeLSHClUeOgSBlkP3czoGP+bd590nvX9lYFvtNcNoyGK6A+utXHza4d7OAV/aOQ6p
lxASlRK0S/S/QrT8UatnqtvgvlDpH97aWLY2MCSRvhT3ENdw2iNHreW3YK+pXFnsCp7G8nbAZU3N
cSonZq4ZjPFeiTc3ISYjZi751jHaZ7iPZDw+w/CtEsK6khL3IRa/gRoK3lqXSo+n8d1OjVtKC9hT
dW2q+0pn+eOPRwmkBttXrwXgphqTO6BRbZ6rj7rowRZPDGfxJuzx3R1aIoje4sq6LheHcQUClmOb
ePvOnuLaSG9ScX4h/XoKcjZUSDu9i/xnFTzajMaTprIh8AcuUgtX9/99CdeFq5rFvLTK2lofljSM
pYKyyo0TdkfRgws13rhGZeLk9gfMjwj6cS8kDLbO8hMmQHqa1h6Mhg9W7A/oxBYE2LOYy+tx1iGk
QKJuera2h8W3oJjvnjfT2KzzLZrlN/lVITXeL06el1G2ukNLUqt3EbgrI5tweq7I8UpW4XXE91eJ
uDzD4789tMOhJQstS6Z/yVNrnPKf/qyZzfUO1aDAnorfAtPOHlJYFxUEqEVQE8MgjasKNQXPqo01
KkNRQEBvBJsJqEJd7Ou3euXPHdklzBfbBVRMt2JlsaRjcWxZ51mg1BH+kCOJIh3K7urCw+8KhIb/
Iga4vw+l7bKTMNmiqjgbmkoN8OVDs2oMGz1faZgNF0G0au2Md/RsjeSJNOj9tEYWlVAqYWjg9Kv5
Fs7nS2qF5w+NuLtx5HTsv8cMVihB01/Tdl+2gNfQ8qZSDQ4H4M0u0k92I5e49T+1wB8fvNABo28U
UfAGL98sRjEN0DnBDvZkmo2swO3lOI/6vbv6ZyVV7WPhFmGZOHG4G2zp25O0uboTRSI3015t6J04
dCIFKvrCz9OvKqkwWdlXVKdKpyriBwS5dbpfHHsIgW/2xDBdei3E6g1dlzajzaBUJk/vxLBlQnDD
nM3Wn+AOGIcUmLWHryt5feCfLDOGzd0bbQKHT1nGfLRGijVqv8VqAUUVk84/erbNXPsCbz6bGduA
QStwVomloPi0gsIkTJWvYS0ub5eR9wAPLNx4+/WSGGduGTLYhAVE5YTPEEs5WmU3eN6tOFKZTwpT
OQ905JDFd3e+p2JI0rkilCTc09XBlSSa8MdKDVUN/Sd017fvxwJYXAXr9PBL1DIrPLNK+nGq/2q9
W/OsCLDr0jrUknvNtLIFlbsDD9FgW8CJ6/QMvuGzg9QY6jggXOta8eHgHqP77a3SJButTTdL+pSu
2X3iM+M+gad24XcRw3XPOihvSC6Xd8xzGeiWRHAIjmBbJym5xpObGlcmNj2OTG0y2lCwGDpm/2Sx
LBloaj12UjVoX304WCnwuZ0YUH9W36bjiKk31qodpr6wNodD7sRrBtyI2SxRJKv8qr1iCWg/cdNQ
QLrQmbwWSIBR8iirlnyVo71Tn+W4OhWZNDDScGzbiZhj6mHbkGPxiFTUs9ttu/Ea3UrpAlMjhOJk
3O2OvegILZLmL/7aQ+jNeE+pC4LdIGXkiPULaGR9CNN+HxbuxH+bY1wNHWp6Q51W8Rev8LCXupGl
0Rw8uiAhfxYdzP7TuKXSZYKELkv/5vsCMmtFuEKrHsje0j2m2BuBXULQmNLXCdRFxROxTXk3JyoI
eM2YggqebfOuu3+aTmSecnBT9niC73BK7m9p1C15UsHlA3YE5au2kZw2XzmfWGysP+8zS16t7Bsx
HLwXrpE14ljw4eq5uDYtKwYrQDZpwbPfBB3oeb5ErSKaDNWPHtJeahguwb4fs1sqtUxcXhLn2+OA
ovcBPN0W1qNkXt1haBNW1Rr5//uDOl8WuVtcrNfHb+1/e+KdnIE4S4ahdUfSYEWEFaP8p/W74wEh
avPQDOGMUNCSQ5J7rkh2iTwoVQmwE3KIfvanGFPbWNXG7+ceZWnjXvQm1kayXeEB3u73T9KUOqkL
0fGoxViZYQylYjFm62NOZGw4yng8bOzannUGyuk173vIEhRL6qQ9YuUKL1zQ0mkIMCIcQ9ViWNne
LG4Nqb+iy7xGwIaunbgw1uQGn5L/heFXG6yvD2fyT2nrCFVOJ/Y2IRRdS4KTKyjWZYyMthZLDTH8
OoQBwvUEuPpoeFK8Pw2XiJT7zXuzDW7NPh9V0Kcas16fPubUJ2PC0OZxOrARIR4ASGiY5SL1pBks
UDRO6LTH1HI9/rLs4LvEh6sfKvLnA/TSHW4znrQE9g/TyupKXz7MeFFn18lIrjwfjb40tvHn40TG
+ywROpY/jZ3avm6bjye90Dgxafmr6M5NaTRTN4pquuPb7JCvExM07mac2zaUYKOgFQgpe1zirVwT
DbGMLA3jqx/3n+NItPlyvDpx7xPOtAhEq4UPTAUYRYzr00T5HKcUF62Ql8hGUk/gNd4j5ISTkSXL
E16i634ErdGWb3QGkiPmDySEb5XX1SbYTAIYzoKHjrzsWCFRo38gIK2cxJS0S/S69KwnKbf3heIq
7655+mL9+6xcBWuhee+AD/tzhJyjrUPLO1YwL+Ii0jDROLhByEmRGyYuwu11KXcCilQTbmyfkOOQ
q5TEz7G+BmkM2kBVBsL1YYqSWg+Er2CezzlVcJNEwhsgA8UgS4DnmAb5HYZgeqtvC785jwr5B9sa
vSAwfnExBAIGLfBPjJxyw3O5Fe0vG/DaQsRKj8eWbLzYOzZvrCaUuLnavCWGex+5+23kVwYs/c1z
jAgS//l9dU94R5YQIIT3Z8CbOzNlvDhPKNHM2R9OR9pqn/wgnt1tHNHGdhzlcrRow3MfFsZL3x1w
wPU0yL081uyE3owimY07Lp1biPxUhrhEnMOIfXzCTbgflxDnQcOY68OPBNwsL5IFq83iwL7NW/Eb
h8t+1K/iZqgsYmE4HCAds+nkB3LtlI9hrbDiYWe6e1ZZs8YBKnociYDxDUb/O2xfDwM9KUXuYzud
YGWZRf9LvxTLW+Z0FMev7i5UBMbTgzY0N6zOD2G2a0R3k90aa2GIMaEJPwvh2SKghrn/hq4fPtCf
qR+w7yPKsC+YqzDTvwujrRsgrh0u/yJWaUsmJaEoC+Cm10OpHIku1SOX5IDKGB9rpdVV+PDM6ROG
mf7Ha63Ld9ZyHaZRzFVTsFszkkoDP9rdR/yj91n6g/ICRBg9QhEI4cOBhdRkEg/VNUNJQsWQgyVx
v07AM1lfWAPz3M5gi7iiuZRDPkFrsBA6PwNuoY+AGTTD3LH/3BUCo9dkU37CjIGeO3oG0G6g7ZFK
3GoC+vslUjfbi72y/d3kMYZOeyZ2mEOQXnVWpVR0u59K5jhjV7RB8VUQnH5zZRiXiLNy6lCMp/kL
7jYFbbfoXnmOsnoCtcwW6YfrL5UPW4hpD40+huijHewClGTYXVVhRMt0Cd6FKAjUYqgtthDse7WP
AVLD1WT0gsatefSfX1pNBsQlik/FteSgxMdaJbFF3mW+//Mc5RhhuLs23SV+yan9jV+NYZNbk8f+
vv60puQqXC/251NTbvqqqf5QGINDcOXUcdt9flWhN2U1IB1vZ/ASad7DzDnxN1BgiwEse40cQC/u
3wgSFViHGjnAR68znOEa47QcLCXc7lOusLVPJvqNJi9IJ04oRi2W2kL2VixhopFRSlBJUlbHNSE6
f6CEwph25gmla7/vxDK6KEm0on03P/F9oEzW5w8dNcOpVLLcP21rR2boHBo2TcKJdPR6SwMDzFCx
NNTY3eQe2z6EoplwMjLXrIzSHboi2qnKnjZdjL4XH5cj/jLqNXFNtgTOmnG1O1ewLN/FVGHwKsPc
6V8D0WrAXj4lAnH3bJctEbd3rMGPDqY+jxbZdiGVVeLqCj+tqM0pLfLR76WoJfwlODUgGqSkJtdV
mUUTdgIOVA9gCKH9QMqHTjKo0fhejwC/KPpnRhjBx8DYJPnYCdynFaNA30HDcNmrS/+HpP006mOl
7Gbw9V9UZP1FvjopnI8Wmm61xRWxx349IjK0zSKCOKCA9SEvAwopSQvriatSP5uc90iw39YkfzPj
9qWAa8j942yZjW7xuuZtBS5j2+a9bqePksxr1ShjRiSnzMMX1FYJ5fK6qpLOlHTtn2uytlKfEAFO
JWJaMswmzKfdiS1hhA96Wzmr/2viXYEZVS50FgB5fZY8IupShxMH5/rBYTkyLlWReNOjAHCgPMTp
/B6tkovMl3xUztxjttwTF85VHJrW0AMz2urhAsUM5SOtrNkHB05BvFKSpHxSUuUBo/ExYqVt3c/B
XAjnFRW7p+/drgY/kcKgQB3tmgF42ofbN5IKbdgRczNAMt5cWcpMNevnCRSXqDmKcF1GK7eiJ/IO
sqSceNgPMd4L5Y7QIULFowj/N//Bb5IIM9advGl/1PMuDjFkiggAK+EgFQE5I0uvQnA/lFyzlMvB
h7V9cvV6ppYhpo6vlgMjtDm84R5sFQOcjVeqnaO+qkBLdtkqhJUbzGy4y278+4UEmpZnsND+oAym
Jr8w4bUoxr15o2Gv1YQvdRzp3cLwid6tWfsDb8PvKnnADcJZTwlkcI8TnnZu868K87fymNdCkpMU
jKNiNaJVsPG/m8fGkcFiBfEQavT1uVgpUwclwtvk4oEF8a2eOeZ/r8SPw188El/07ovQviuylJsw
MMFUU+imyJTzG09QowWQxivOAFbciC/NkIyHdb4SEQMSbnCr9+xjscj8vR0Nezu/88gdmA+z056f
YccPzAkK8uBcyfiC6121rtJ14TD8LFI9loz6oJBcTro/MWXod8Fi2JvahPGZW51Tor1u8uR/7ySG
7CFgoQXd44pdbqsIP2Sc1RTY8nSEa7YrckoERfELpSd1lppn26XwVCwcUuaqMmXMJeumA17inuXU
eeS9pdM5EPU7QQgvjMQs/DrPRETzzCln7BRA3/H9XBp4Y1lTXWYDTHqalXeImnxNTpOFsUiHe5ku
xyefEYLtO689R3dFTocjblBZyaLT+gZY4fzs09Weslu7nylaKLpT0srzauMTr0P2dVQbs2RTYu0o
iJ5+Da4skIZlRMUbMGrt3WH6T0BwDBkw9jSUgpOpDvLUAHR58F1YWRBbW3lGcoV3vbyjUAvZw2dR
cL2dckk4YUgxzRg4iKIxLl2IEaWTxVwyyRaxhtFn33hBnkyw11RgHQFYJXjNW3joSq738HW9R46q
fJIr/IJ5U/NVSFx0UNobw16IcNFE0Xh4F9upAtx3nuGt76IfBf5cenZ6sx/o3/Kx0YK4uIiAMdRU
V25vM60Vd0bSmD7ZhME5HKjeONTwsXqcb2kSzUHCTpoHu5stOTatVgXowSkT+ZbjEXaA2QiGOpCs
N3NIOs/XKdMjf//vN3J5aYfBWEz/mlkBcsNb1UYgDDBizwXr8Nujs2oR0c6hj7mfqDNeEjwgGVqd
XcZkTU7f1PMVKghJQeReZaoq7NTYuLX4ngbQqoLhw/3/YES2yMSSVlVV7cV/MpYWej/scUtCrDeh
2HxQzfLAYjl+N0hBm/YFd+ZKXXfpknxujYlaW4zsld33ve8O8+hYn/gJUMTmWHnoN4owCgAP+8pn
6lU05qUHwpqsFbiC/XS+SwkTeIqshtQ4kYo59YDNEylM1qzcqd4DZ1oMP0OZI3OyKqwdRbCzJn2d
BuhbvyEy9K+IzUw72ri950yehPdbz91FCmU8ILCgcNE/D854Xaxql0Jm+a51KaOM72EKLRt8Mo8g
gxT7nH8cnHY33zk2SjI8l6P+ZO152snX89rLQEG8e7swadZ1bFF2V4zaEyyMJHsu0XwHSi/96H2N
uvdBCT29aZMv4sKmOHXbdmrbFrhaW5/NN8Ew4/EibPR5FPn8p1jufG5eIkI7dj31hh/uy/A88FSZ
UW8LDZLjxDhz+Ue+oryi2D8UNpwa/HxOaO0H4vYUcw83zksZ/5K8RnbIIKme2YpHFtkw7myn8ldI
0FnUiPRHBUrJAhHqIpRpYrG/u+waItxVA8tBw2cQ+FH8kuMv1POwxYY24a8kxwxZ4CM17j0CygG7
wzB7rr8oATQ3T0h0HwUu1GRBt96qRkU8PW70nPRglbqd5DEF2nY1jT57kbUWZOsJO59TVcb1v10r
ZjBGREoo1Uo/RarajBeCiF6Y7vLwaI3UU4HWsUXktCbg//jFbvuGbO0m4m/D+Vm6dNwYF7F/OX+s
tFxliQMYK18DB2LDuMqDznrIVnuVKYVf02Hgi20JaWQiexOukdMhBF0/Gaj6WUecai/3C5wgFX2Z
HPgsSaUVPJPwPETuqMyXwb1h2aXb3/MB2waMLlKvGWb2PvEiXfBqvk71m5oTUl392RbW50IvVSVq
8FJr2vkyUfMblfRIm16SMnJixF1yrfQdKpo+ciL+WS8RWOP59654hMvI8LSJAu1zukfV/2mY1TW7
lZdcmrYMyXgt7KnzxhZ5/WnNFLeALHd9vDquZDfcShidEDJQl5z+m2xIX6TmuAGfnnx4JRaTjCoW
hp/7bvUwSQr5moPvqvyvQZTYmrq3ChOb6tmLsRcEdwqwAMlUuScqm5EMbhANhJB0SY3pKcRJJYzq
2e7lpT1UR/58/D3o8eiUYMZ4OfyHf017g9uBWGOAZvql2geo1MRXnmlHGytsW3r+HlYiMy0TOnJI
TsuTLx8IGIAzaDpkHUbgEY+0A+8I50W7DdKklYqJleRHa6ebOkx1y8fEpk9jp0b02IXlacGfi4j+
jgWBqc4b6WAg2XrzmeUKihBJlHixNfSBxkYgJ/hFLhdabFz6owQcS0VmoLANqbgSAiFK9c7+tp3t
LnKujPz/DqcDZzEAhg/hgVO9IYTeDBUzSjVvNqPWZG6cNeHJjSqUaxACizF/pYMFCR2xfELWTN8D
KAGw3/3crJm/TZT1ue3N+vd5Hv57py3nroPn1VCjVK37rY5oHqzOnPGNqV012IxZr8H5kMizs/FT
AJr+eu5S7GGEJXJ4Vs7XmqCaxp98cs24c+uDZtxz6X8FxlkymROlEV0VvwQHyWQ14BBPR/qS12wE
rbI6noCpCBgq4pahXdijzuZC5iioe2GZPQVdb5MIlk0Aqks0OEiqQQkKJT7R5SBoZhM602/l06ct
dEcc0OLQCQENhTCzBa0SjYoonuZZp+PUtW512HbM2sl52xBzknNGKPiLIfyIeZrj/SPgJU+rWQEb
QC3c3lRQJ6KEQTrPHdI0EVIZlEpb+HmHuWAhzdU5ZZhjiBdfOSforwrbgByOUx9LBdHgUvw6QHVE
jq8eOVDyrF7pVwLo/U+vtG8hD2+j5E5WjPmzYffMUQVSwrD1oNChc+tbni1qhcX1lG2HciNowjdW
2CTxMnqIVc194b1Cf+YIquGHzjp3YLijBkLuD4KjZlysx99TOWWHzVrixHlp13BJPwhPogFQsY1i
Ntsddepi26Y5AOWQe5Wpes4fM08UeLt1IpDK/tsmyH3t+m+uGbPkmCzP43Fg4WuD3IXNnNqTYNLw
AE8a43V6fySuVfnW6+XnuWmXNaG3XBZO3vISR/7sKMBWfllsv0iq6Kvr0Ur3IXKfwV8YGZg9BaST
Qbe6Ro5g/jv1t4wE0J0wjj6ZmDoqWyfRZhbF39J2EB57g7oKlHx09KBqHCeVEAXBb9AmubaslCey
460y417PoJJrhH/08FoCQwr6eeCcwEXvTKcmubyoRQt/VgQGXetE8Qi15EUre3FiB6iefB1i9C64
1ZBHT6K+Xbn/95e60CLrSHJONkAOaJVoJVW29Ge+jeLl5Hrx40VBHAlyjlwZ1EaGeZFh/hmUXxY/
l0aQKHkH2Nk3uspFLKJjIy0eZbdQHBSMkBNKz41pGFYKCC29pFzW8Yt3nEZB9Ec8wi/EDFr0mgvx
yu1Kwh6oHxA5pMuwenkrc8Tq9xSv6k2gw+m7A5g47WTWpsPrhw/7OUx5OrzD6PUdpJE+ClY/uMLd
0OMDAehZ2PYr1WPDrgKleRs/4Z4UGYLZSxoJdvr0YorfKKWjZeJumlAzSCwF2VZsigvI24wtTy/h
+1dEF+OT8HBppWN8tq3o0QngehDQNLw3teRAV97IV15XJDsKwG/XNgMqI/kDJtxRH2SOpVV8z0P2
g/YUZuyNhG+coYG0g9pymdN0/uO6UJhlRTLHgDYMkCwF4zZfBxHBK/YH47NLDnsJvVjmVpDVakOY
fr+MMu/D47+SowQ4KYuT+4JqcxHWY+JYTrFQqsHMuiD+izDGMdxIHGDRHuJ8vcAOFWZym6Z//iY1
1Pe7gCjvj6fiwEC6Jvoo2IeYQBHQXTlB4VjoS5ZJUPLrGbTKwoCUFArKwD+t28ctlTL/fDGt/jsn
d3kbflI3CezVHa9Xlw0mvsSRd+n8+wYX0fyw8Cpp85LGLVtpRvaTo9t1MxFdWwb1UDmVJvBvODff
1Nuy52mNxKMzNjzxX8XV5ZewXr/t7M7H93SVzK3W3JdrDeqRXk1QuBV/As22N1jmlRF4mr3DhLEi
rc0iBPLfnTZw0JhbyVlpcsS2v9BaRy/4K0uVvSLw3CIcBTml4sE+cmxxU8Ty/SxZhQeqGC+FPVQH
40+5xNlLNZYg+zaBCzCKHCp7XvVX2IxnfqByZJWMTRhg1J9CjOcBwmIARvGKvwBAY2Kt5LDsm6Vf
Wcmea0jWYgmv0+pcU57qx4UnqTAWPWmy1RHYEB8ZSNqYlC0LokMxi+vV/uF96GB1y+cMtE+3+1ID
kz+CQG5rZguAbq8ejxp3/KuGf3SLptOTPa6TtbvmIKt7+OXCtoIW4doZTSNij8d05zkcu5DNT89D
RaEktmAr+HysvuUilV76j/LX9uFQjnDHWPGE/9cgHw7WfFRZjX6FYRLkaqSBmHhWZP/g3lxJAtbI
jjip/Wwf4t4RaNCDgF40oKROjT6jJcTeOQ/1qfAGIgsz+at/Pvmc6u7QBW/eVLHwOyW4D2zxhN8n
0JE0kx0cU/UXJWpKqFTULIWTECohazfOYeffyB2BDzFkCqtBebwzaN8SalxW61ooaXX4qDR9TbC5
uYTRikFTNnlCZj+qB6NH2kax/oYY5yGgNlOmWFw4+Ll+FtPcJW9R3APdhn+e8RgSXEK/v+7QemCl
XkvIMjmeeb9s4Cmjk0FQkdbBD6/1wE5nBV4q1lqYt/B+S8iPp57uXZdCl4BECC4wj3cqgwxo+Vmd
LmINn/4lpNtNtmhlBVgPC8+5UtTjiRY2zWZV51iYeJyUQgzOmPfHga2hcZOsPEdl9gZ+4B3T7y/e
d9hxFVPAT/CZMOZ9x0t+nivMlWE6zGoSkgWvuBuu5RrsPNm4PnRezklNeA9/NciHlU4okbfDvMla
BI5UnDjgM+27V9hOTw+rYTwUNH3ilx6lofKq6VtBBGMX7TfV2eHb6NtWb/Wk+H0/II89BOp6riBH
cn1p0P01zxFO26GR8xsrAxj+yv+Ewou4wfhg/hKeQsWLUcMjrfbQYz4tskOHVQK6AoTA+5fFyOwy
wypgdTPIrKb43xOrwSDQmZQ3LF9vUuZB/HqzOEtNuPkEZEgZjIs0+Aq5YZX8Z8iEIgsT8LcSf+l0
ThgyMlpYdpqm06r0rsp3rK8ujlJlgsw8sM61MtJYsanrsW6LI6/wFrQY2ceyggj+Mrw2zXej2TUk
WJH3lauuF/Pt1znqrktduDP3FukHW3XT8gFiRbOmTpgqrM68sP/0ffmuSXNq6MQl2i3+vxQQkUgk
IKC3E/o1bggqpl4L4Y3NMnSO+T8Rz4K0VLbdniEQzmIG8miEkWsKDNyxCeY1fgmRk43G71+yLqiq
CjXFQlUp60pQj0aYQcX5CgPf617pnt84X6G3Yk2QJW5HyTh5iBopHy9ZZmbkd+iv4DqNwHrLQ74f
PEHPA5xCwtBDgsVJ6p9pENRJtS849dP+IMAlCJKKHYZBHpJGoJKLeRHGNDPflIu5e9OcKBGGnqCH
vWewgbr28C8Z/tth6f22m/6OHoBFsII8TzA+mJW5zp17Huez8XWVGjaUtKWyqlVvUZJdTQoLiRXR
Do6T8dnaL6SEf9StNdz2K0AS6De44444wqUvHLapq+g0ec9x8EXJ2f9VDwCQUGDGPNzBK9kbqbFl
0g9mD1M8XpFxyOqiVuzxe8aiwr37q9jirK8MBUscTmw+Ymn01y9M/j6bwFgzP1V2RE8o+WuSPFpC
+uwNe3D46N92M+4uw6h1L+t4GrO2VshKQgjc3Ja5y+NTxA5fgpx81lehU4NemgsW5EDYANAcJpy/
jpznUIvoO2J0YafX2C+Ozr2Lj8F8sJsy3+zaWSz267yf7VIhH1uWUYar0rJpth6UzQLsJFxhMAbg
xDD8j+sSR3gATRFou5EWrKayWXg4dQBIoOFYIlhYmg67lmiR3g6lBbAwLNpqrqtWhDWnfH1Rdx3h
xg2KBRMwLz9tamc0kEnk922y7mBckivQjYZKe9g6Gcm1ei7ATEUhigAHQWCSiIglHXqMqORbry6c
xpCMSfkfhEOhyTWO8W4Bb17t/CR5zNvwNtwjsrHhHmE0jrC/nc4VB7JRO28jBaI3dkgXaYwS0qKt
ebFfklJJGq/fierp9jIvEaru38HNKDeRSaL1CKKjuJqTUV/of8gLPwLfVZxkZZs+OsKOwTxF/UcY
7jRwOTYsVcpXT9U+vSQbWoIX4MLvG7Q1jAqa36+okpO4Ty66Kn+u30qYsp9oz/u2E6tO5zyZzQaJ
JeficxDqA1s6alngxlXRkHldayK1C9bQj9AjYv4xrJ9meFUO/YiqNfrybkwIrqKxb3XH8YSTFifn
ZZ6PmQFXwuC9YQODFCx2aJj/yOPUA+THO+f7ZWms8paHg7p+ICETS2w9mcWxjB4k7TAyWMq4pjX/
2+n2IrbxrUHZ0cGLf5Obb9iZ2hCKSEk9xAknamVAdeo/QIfroCs5d+81QJh+Z5nLH2Ric0zYzbiG
KPVSpfMhMRhjoGUMjnHOKz6/6bOj/vRcpRznjIE86ndydMwWctwSLKM4OyACZ11a3gOOFfXuZBpR
u3QX0BlBO+J8VyxsT36XTL4Uy3BWhiZXbYLmxkAnQrj4IZCLhYdgRq3reErADvSu3c8DrMlfTdpQ
ax64SqJNTuodVH9TIrA6HEYvAJ0Kt+r8M0bgCdfNtBoxM2+ra68crN+wqrk4EgflfpURWDrODNyC
58Rh6Je9CHKryUnpjqTBuVQPQUKRZYIRj5BgqMMvCs5N59Fy79YXuUkHF2mYkwdbuPWFoEY0fh7M
pgakp1iRDPYRN1m18E7PI5pJ7Jx1GsMW+4B/eMnxb8K+r5T9ESPbKEBoITedPEw36cA3YK44paVa
vpH4IfKy79rCdmDHlh7bRBXBoeEqdxG7FKcKkLZz59nMkiz5PQ+Pe7Oo1vojrnOctbSVPLDrpn0Z
IzIfDJ+2EOqs5WEq1UtviFmxQ5k3eCh38Nry7hy3po9gMv9woMdiLlIvxVEENuEw1dQ9snS9FhHX
4SMPsdTuQXEVFqon0uHBIYHC+SrlAdg+OY6PNtWHwsnVWUZXmcVW+sLhdvVEVYLrvzbOO9xFhxgp
S28lX4zExMLF6aM9LVJdUOek4RLWqifLnjMeRL7qazs5fMo7g0B6nicH+gv60yfJAPeGis6Jv06H
wRZFQjRmyh578TpC+MMCgUseZW0IqA/YnlJbRsAc5URjXiNll1nt/4RVTVdroR5qnKtQc37147zn
UY3tFWZ7YLG+xhymy0hps6Ne5v47jJdvPQbpZfio9UmslHGbK9Jus+cuzDKaa2yxq2u27EZBgVhs
5apwRRgP+nZEmknDKW2/gucvs9HwjY+6VIq/pSHboZl4jLUSxvpdrQ9OULjPVRuhgdHV70JW+8Yc
U2FfuZd/wfIgeRrQESGkRCdkJkRS6Mph6KduLACdVxShujMf3H+7L1vIjqrwkPCfyJJMDW7UhQYz
Rtf+x1DCe3Dv777PTgB4sb6VKA40y5ZGWB2yipjCZ9nKv29Qna6XbCT4KZmzrY2YBij/GtENwn6/
yVjfvJkyPIi8eEwp3s9qGZbi5fwHSqoHPe/B4ZrjfKym9peDTjVZ0e1kY9Wr0NsERsH0644lFnnw
ir2VSHn5lU3SI2mAQiW86uEGlQWUpdfL5frjQW7UqLvtW3tAL3uywuslVWSYEGIf2A22NYgYjJxt
Wsu4ksD9i3Thy1qUNiV/X8lX6uZ3i9xuHj+L3FBH/ldD72wjm6TWk7wBm0zv1pXdIkUVeLiPY6hH
ihNihVw/5kZQBeKLZWz73A7+XUD7B86igBlwOcEPXRWzcvVWvznYjETQLaPIjU7qHNKErVLI/URL
eOCutk+7TxjCb7TnRxmaVlDTloBOG/q3jh6pE2Hb0MuKy7LXc0Xaf1WowaQL6L9XND8LrGFgbqC5
9GPhDaqx6eDd7f+q6BBivClU79dfAVgl34Dwr63NuPA/FqXzalHnkfzN2l34rrfJJ+vGF1Usny2r
ow71JzDW7FFvjPdE9IQKLINQpkJj0BUU+6p0BC+9EaK5LuIjTSZ2YcFik/ZeaJblzIk3oMcTqogI
ip51sNoRjBTjD0QzHRPz5DaBuP49PUwcESbjXvf9XtLSoQeTRcP6xXdh1DFtYDUfTsUUcwO0SPDl
lVjd4RfXNXwpsJErJvZ0WTBryeQdF0t0ETXDlehrFLj/B1T4CO6W/ANhoBxXw8xp0OpugdbMCwjI
21Q6XJVU+/uLiEzReaoQWb9x8OGKVv4l4VyIrrREAFPG2FgZ3lbIvWo5cITGVOxRExV0fgnrA08u
lPktQJQ1BNCWCKryU5Ckwr/2kNHpHXIJQXVV17oBSA9QyrpWsLZPuRIG2ukeYvy2qPAJEaJPckKr
Zm3SXAzSTTFLwJE/BC6vVEebo9WkQVvsuBrkK5BG7pAi9Ydi4Wob+92/4FyNy+de4b+wy4k3kqe/
Ld0ReP1xNxqm8WLrfkblBJhqlKZyhzwpbIXjw5u7acu6yl027zKr6mTqFu7RVsPouSSzs/s9/ke8
4MNBNUpD378vy3Ji0yjRbr/esoRQHaoqsVhC/8c2NCpuxMtPwVGM2zzuXHsv08bcJVekCXo/G99Q
GbxFbodK1absgKv04teQaotK8kOCCihfxTZsoMd9LukHtOcpNfyn8/Gwi3G3YOYrvfyXS712AE0M
mRt0ajaQUqv6t5t+QL3qH48cDlYu4Lx5odEyT5hzHjLRlZtTlAPjPHKEK7wDmNu4DqCVo7wZluOy
iOCs5z1XgtygPydjAUstdBQZvVHNDj2e8a16pg2X5NKyK9OkOCIwsTJ1LENRURBTCc1vDR076KyC
LHcfJwpIclR2Ej9UglDINpOqT66//WDNQ/DVuSp6fIiGFm56OOYElYB6RIavDuDQb9T8Vcw21dLY
Q2O1+onP1ycZB1MM+cvyBhVZdXKH4hb5Wa0oHYkUiVLCM7fX4VVjTz3XVQtTvvR7wyqJqUGaSzIB
FArlDgcxju3IAtVhGfQj4dI+WCSrg44Y+sOrVaDymqDUn2OPt+3ROcZAkE+SdA/Bwh2iGELIzEr/
58jme23oqcPsjuqfvIbgjmmh7YJn4V+JYRtkRTnsdOqnAuBPiHeeSFeDOked+AGTGr1/wCqgXDts
CIb38OZy0kTMlRJ+z6AulaBEu33aPY3J0BqMA/hAsFl6Xq/OOBhhImLXJTyeR/Of9Noe6z/XP9EX
OJ/55ZS7RxCaU7imqh0GPURfIMYLubiymKWTb+O2saRjx/UoB0Aod3nB2BMYjhTEVssyK3EK7Hwq
yeRMuCcLSI+gBhqeqBXBge4qvJA/Mm/q2hijDQSuZN5aS8O4JQGdrmYtq3e9lqPoCmSzil7kMfWt
z+TVk+/PTYmU3lUW5HzlmPwuTAGLiGMy18x5+zIxY3hOV84DbhP7xcKl5UkME1SLtpXzVbFB82kt
q+PWfmItxwJKk0rvhh7sye3hx96AbbPdeGcot9yvsRZTozf+Rv1TlpEGokdUAsB2W5USQMDN9ie8
cUP1r3S7aGJjo4LkSTueMfudWeKKSSxl3ib94JvCk9yL/KI+IvP8FBkQt1ygCYGEusBqCYLuxSE1
sF9i0sqM/FAbIg7LvWh67xYgfDy/B/64VpXTeh+LOTp062hrdBcm/JFY/Gnk7ZLJe6spiVEnTPR6
hedBeh3RolUp92t8yLDt+MHiGKWtT076jnRxPMRHbV6C2qqOz3VtKBcDMqfNSdx6AKYcP5bwg813
VGaxlkbdjDBTtpN76iYC6bCrcgLvmiVRvd4e0yn2IE8I+TapaRnA1fJkHi3Ex5NjLfRn7LBTyJ0r
othnCU4GcA2BsTk3Q0M+vNY958v+Jg+daQCUrtEMlHFLgm9ETcYvSJTONR9eVJC+DZQzBuG7FZYP
JKSmKYkxkoZgxRC2R171bWr0kTyOWOvVoWE4oSbest5LuwEB8k5mys8jb6Cy9XQoVcKBMK1RDZxX
NVcamCjlbRVoXN+7/HBGSYTOYVxxSN+ZDCIzSguU60Mwm9YTqoTYfWDsNjuFomAMTGCne703ZmJQ
jwxSNlMeMRxyAFOSlbP9yRRFKa4qRBv0o8XJZh7NkYL3pFyVDvS2VdAW/k+1JmfZ+pkZAugikFDO
1uHGgigudok5r374FGWbRLPoxTjlKoGbgRg2hbcbs/xB+06G7d1h3c7POTkDdozrpNc+77rIGj0q
TYHMAsaX7Wuzu6LBIgKP0bQg3pbfbNa08MukbYukyF24b82pivGWBqm8msauyykP/je2zBI2+YFO
zr6ekkkXxFJszghyURA7BAzEnHfvMnHSe+4/PqSvkNwIk4Qd8JBIx9+yXLAtXZMaXTb4ZyVtEO5q
7jUY9GycANodgsZnld5jhxCqZ2RMA3KOHhHbLIkT7ahjIiBC1KaH6SmEfZqbeHtdvLWAfG4Nc38V
2mmsbg6A0cqY/0yWOeuryzKxw4widOxwHzYOrsbiXPmMHBHZXVvB54x2PXpbjGVAeq2h4Ye/hLtt
RVTDzu6OeATT+f5p0zKDIJRgpkTCa2UAIO28kfUNnlMhJ8S+mClStiyzYCbc6Ua+O1ZGQr42UMQ1
xcsMKfeusQGNYYFlwZy3D9ZY6W8HNaO+5R3GQ5kYQVTlDMMT0+FMsxOVjC+NTGxRdIQ453zMa8FV
TxO4wD2HNhi/QNsSTvGCC2zHYX76xt7Q/vfxyolWWxErMTD/zJM2MNHnrkmGCACHN5jnkYUImDZR
UZKh+QZGbvoZmofAjIiyjAND0C2q0G4LyjbfDQCnZTDKC1+VZ6FL0dYrxVskAhv+IL/hcoi4aIxH
XuzgZqOmZfui5Bl/Ci0L5T0uySYWXEcSDs86OTuqomwUZKN5yGfnUw/gCEwreJvVQad2puLQInpm
z98/KWlmWV3qDRwvgV1gauUWg58Kd26AVHUdwAZge0UtRyuxQbatT9OyWRHMuZUhMXyvBK5ySKgc
NujhKQiDhTauFKZdBCA1y9bHqtYZPG3S0BWJcmbrmtZ6P3eJ2XQbMHSyq5sh3phHvwi4wBluY0Zw
cH2BkG2ZbTm6FWtHr+UukJHIABMZIjrauOU9B67VxCw/VwBbN19fGdZ+CW/7vh1D+j9zKRTPykPN
+CPp9adAXHMGNDVlgzCDfgUMwsSUagHsVbxY7JtgTlRwq6Mwahze10rWL/4exZFF+4VpHE8QQFMT
P+VEH9916F4h8O6gdqJhKBn0+FYa4xEB2+MUJXhLOnvyns2mNkk9J8kZ/QEwoJlZGLuMOTa/FzDk
dSvbZ7b61IRzKD33jE346dZJ3tWXX+YFHVKcV4tKHKaNfBF4zPphrmpYggN5LkBVVtZ53DO2SJjC
2fmvhOGDAGH2Crz7xp8XgqOM3HoNkYh5/T3R9jdPwngd7bsjsE/bgWgrCHiZ3FIH7Zhz9Y2LkJYH
3I2RGqVm+ROUM6KZQvnBZ9+M9kjRp6VaIjD0pL2jGi/eCsAaQFUGvolq/07dT2WYk6+TATP2BAts
fhsQJ0cbsDQ9HEJAwWdCk2zNXN4NVEmzVlBbRLAA/y0Dkxb/Xb6yIdquFRzRwtvOhC9M4GmYV/hU
cBRz80PhY/QbvD1a5NbH07cGdWuV6TtDphoNf9Uof+ScVGhcfsdTszJFqB2Ne98+N3lc8K4uC5sI
9vvGbibI5nql7gSNNT+OwfcZ4htv8kYzVRLDpcC57D38meJBwtIanhXuhWB7ysHlXoTPHLP1SmIP
gkvNJq8DDxgZbPc4Y6bKtVSZFn1eNU13yeqzuTz8TjX1QTL8N5mpSto6nuuxzmhvuQO2CcmsnaS0
LrK2xDX5hBssOnEODHAN0TxjMv8i6NgmuWXVh1ypzSZMCRcAIoq3eaq9xRn6TabGxyUOAigRnqIT
JIfB9fO86nrh7/95vnaBBRQLl13QL5SaOHNjsnE6mn9ELSl+i5XCFYkliPMayAEdlCe7KRJASI0M
BNJObhP55RfC4xgtZ97VnYvkUgpJ6P9zq9KGf3NRBDeqGvGvR1JW4DHel2ehEGUU02hkavyJljrX
r8f1iG2zDXRpa7kzcraYunEYOEtCxEuqFuh2A9on6uuBf7nkndf4vupBN9POgiG1XpNNXQ2QV3mg
SjkE7fIw1EwD46LdPlvv5JDZcov5O2DS4x941HD2uv/mJLO+oxJ9MgsE1eK4qT/sgdHMZiEbfGk1
KNy8i9/8waJfa4aYZs1lcN7gPws1E8YTteJ4tjrxnWu1JTJZ2Mh8rZ7OzO0CYBxSvxzvoBYRwvai
DtfrpB8Bqj6EwzehrBeiAourpos+xQC73uSAqorO/GOVKLE67XVZQGoowch0IkcCfmIJIc+jEzAb
k5TT3IiK7xAGU8El6VNRVBz6z+uyKSmOVRhQkFQEDOo6+R4jHg0io4y9k13Y7JGHgVsiqA7Ccsaf
YRDT8O1hNJ0w82ZSZyBkB5gmzgXAKwqDDwbVhTlmk3PefvEXZuj6Ng7eRpgVaP7zMb83UCJk8X8e
VL+Z3Wjv5f9sphgRWirAGnbc2RfVpYJHA8XaQUs4go0K2HcWOdquTEPO0d7FvlGFQNarUgc6VxU1
v59kI7LR0YuPCgqrKBjkiNYuKvLAnCSKg54gmGkVbg1csbTFSvZmE/N6nNV+niRnhy421bx7Dmxb
rjQfstDOHYxB/1lGAXnXs7xTBDLvUPT3mcCR3/Sn9JBsonXE9CYCMhs7LW4ZK10+SSntsldwSd4u
3+xeNl3LgI0dkL0Kq6Bb0Iz0JGAS04jplw2FPljrqxBVjQIKLvZbo+wfGfVRo+loWwtmyfgQrJ6y
hybj4RFPVgcgtpYdGzWTnpjuroFKy1NwveNGmSK9KaVSiSWdBdwoJmBvyEu1sUPMxOpW+Vnwsv6f
AIS5iw13dtmk+fqgeXevjBFa90QufZXnv2KMYIUjj/YWrypo8wsC9FVcin8tg5ivceILLWSRdiqX
NLWeX6Rn30wCrmFHgsM4mmbqcMz3qUY2evQVbU/FQWf+fpsVnVnKZk/F0vZwU4D7/FucoA0qb+cu
qfMhPPiVrHhzOr/2riLUkck13W1Y8h4r7PkapG+51IZw/uX+M6HfL1kJIbYslzifFgSVX9OHhdeD
ZKmz2liQQvhnUdYx8+LoZ/7MDIBRaJD0c9By1VgcV00dgkSD7ybhg27VKt8v49y3kuQjxZ/t3gLN
vpwpoABm/u2YmSPYV7iuUaZkN+s3aFH4MnuMHZkkB3zwcxcRkOSbBAq2qFD3nKIpOsAwuctcmKSZ
k2eiIVpaApSEMiWFz/5IxbIBzWLhhb4Ic1HKyF0/8XRUxd97wZiMNkocIZNaLh0Kum4VdQBnEWQY
S5xvlA7JGPhsIzQKbmEs3Rc+98bl63gtxhutPsbZqD2lgm1x/2jJeafaYCNJY2I47z+gFHpYKFAC
hMKfRfxkcHEqMNntgD/ViLsYEgIU6uSuvqUpAe6Hu3qErdAU59fIPcBfdUGRdQQIsDTXnY3SiLux
nKtgxi3Nmgw8mCP6Q34StK2KJ8q1wZELIcmA3DQDmh8BtfsrFBWLtaIthcXeTEh7gqDrt/xfYzTp
d+JbyKbxLOIwCC99Hc/4RLDsfTLm6xGAiQPicM1Bbtj0jnZBdW0DhGgEEYDMt/7kZzcoNKnWI3Ch
6u1hW2O1xQUNEUte2JE3nmlHYCWjN8Qv2yjnnccfvPJ9TVO2iTFoZPl2Dqnh483T+Pgyq5uWtBV/
HSIx9k4Pl7qbsYyBOCFU+VinrA3cY0rqUbNqx5jQxSCxiHVeU1MqZfeNHtn/fPPxBk40mdSXGhti
Agyh1EKSC6bPZ0PF3qYt2BHJmzKIM2R9xrAurem42/zEBzhCTEYkR9T0Lwkdif6Ym2YAVprD1ZMV
pctcaLIzmDyGuTzhKJHB1qQXrVY1Djz6vYWrkZVzdJbnAgFXbqE1MJPgpZW6I1YIiD5WdoDkt6Ly
kRXcuTVOJLdMKKGsOModyJw/0xgsqoc7W34XoU4tuXrfJwnCfKgt80Saoc+/r4FsP2pcF12uGWlF
sEh/4ognrsZ8B7h6wLgest9O2ATWvaZ4eDp+wu+aFsiANJgJq54ofIf9hl56K9YOuRhhJLht4LOz
M8Ie67XG5WdH38EWbRfjOlc5oy4l8SksN2ePM9ZchtKeJcS8DrC7b9/PyjWF1mzggG9B6EPDZT+r
rUQQSNsJI9i3KBWz6NMaidrrkoi645WQfWS+bfcEMfufZfsTFHG7jzMy8M93k/2p4G4T2T99Cug/
PEpFOB0RybN8AHkM9JX7AyB7sWGE7Qw5qcDd25BfjNeVuqAyU8efbX4QnapNhF6PMN/Yb9CtCt5e
ouwB8hzE0NVoH/xvG3oBo4aWE5qY5u+iIFMqfyC+6+/f1iA5APSruqJdFFANq+oSVDn4RFYYipL+
5sBldk0NEfat0mM6zzmpQ/PsqPmAEDnhh9vbu6qaYlzqEo8aRxngYAvSuYGbBm6t5j+n0YaoXUhB
o93O4hCVxLRq/M7XlJe5FovJE/lxmbzPKInbb7f6fH2jzpVX89ZgdIqxj2HVGqB6GqTeMsX3rRmU
pBgoyCSNwhIFV8F6oC0ABTgG/LC0tkSH0KiZdIQbLP70e9+TRzRTqet+TeOst5zPt8imAK1D/0lU
rpF+tr5SCwHGRs0cWh/JM7E9jj1y900YX1WJVAyF5z6nLuB6YuD1h5Opick68WAFQd0xR0KXFDDW
DdEZjfTz9SW6ihHflfV4EPx9GRcO6GaXGrLNS0caO66xWJknXQcVGSbeoMZYweVnFsjpCY9Sftak
FQ2X9MpBhdUmnJf7k0dX8Ue6gygRas/DirOgUPcnwfQ++wDNFbPoAFuDm7/7tJb4K0nhSDmrdSph
Y/zeSWL56dS2Uy33iAv5pFNi7kFiSHo4rCFlpfU1/6B1TJo5VUh19FlRXu1Mtks8wq42Bx037Dru
bmk9NAzZPWKY0vHFTfU3tBQ5Lkkr/PMpHs7CfOFqA3mb5QBxe6dYFTc2e+RDC8EQDRKTLO+++azn
BR9HkKbmIpkmc2AuUa5IWwbGrU93b+oYwh7H1GicWafj8ZttTCnaCR9ftfWEysxJUyWGyrMPbRiP
qWOVsy+YaNAVsteE2SUDhSQbMppkkcKkT3y1sHyd8IL2T8g94aBVNMh7D/vwoVfbdCdXAm40Zdld
0ftwc2jR5OdgHBXSVOKX6FzXZOWAbmKzFVnBwD2DwoO1nNHKw5OygRBPb/l5PXMwp+Gfpwd8Xnzg
07eTrA5PCVsvBmrY+PqTs7Hs88tCt5Ceu1XWX7tMZqSbVngCEt6wI6toj6jH1r/DdBu5tNXKZm52
WQS9CCHlqHtXUVPrbJguwyIKz9cOGjH+RXXw4iBLovV9iLLI5OcTeep47YgFJQSS3rBhljdXZRGs
W7ujJooviUqHr9cx7jc29gLLTlguC4Ynfln17zPGb25F26IQqn9yyerrZ47k2/BFN9W5bFytLdSO
ko5BFAtAQaX5mbEvgvNEhojyo/V0oNYjBKdUpb0SLrGWRazoRtWanytaERrhSSHM8gk8+l21OLJh
Pq/tyVpHpANJ2cWZPs1flDN9Mzfk0GAt/aEoXJOzySLvAfdzxT7V/oz2kVjdIlsYAJ1Z3aZP574N
9mTEAAWPhsbwmNtx5Knn+NJ/AhPQS+Wq/elLRh2TwoLfQGkbI7nueGYkkP+X+QhrCowNpMqYSFQa
Ib4ljDpkMiPto6Ep7TQXr5qbhKgoGi3LlwTPFoOe5uzBxhGY3htkLjs65E4k5C/eFndpaeG8Z36d
lT5dcGw/XNKKHl6ArP0YqzJ/ZqpYW0F0KCgj4ZXcufcbHwbz7J9IoUi1RXBkUAozYQ7o3QLAQdnn
x59mPNLPMZVor1xRU5pe60x/s4icxC9aqwTluBYE1OACazJiT0kGvRTn9x9nAPl6Fyf3d0j0QMZ+
RxF8vsdepM+pFuKwG2f9NN3PJmrqBMEOTlrQtJSIwte+XPNLcmiHWvt1g/Qov3zpdZZssTMjxPNs
FFecieWx3Z8qDeniDezc1ms5AeJJg3LU0VLPCa2aYxYfGnfsm5zacjKiyiZlnWfb2stiZq0c6aoU
hDxB/21gMfnfqbrMH0yy0WA8m3oO6P/cctpt3DdT6OiZfYo3TDkk+WHEutRzhsgm9UxO8sGxknVR
BM1pSW6tQm1/bf55QuRbbM+DQ7J0khottmLzeGDZ+M54Sc8I+4+SDiTJePRt7WWu+iXjpw08jEOw
vLJ8/z9uA+SZ4rpp62RerU57kDe4lfLiOjfKTcGXpGRE6zB1EMF0086XsT/P7u7Y6UZGy+alvQuB
JTKpB0XrVXbytx3xcA2fhqEUSYvp97zRJMneB/t0poiUneCHsb+qFuSXf8zdrmn99N9spT7pP3A/
LNoVbDndLfZfWEXwAisrBDYoAS28vOwgzrbaP85+DxRb0YmqvFw6NO0NcolYDh1Dj2IQ2/NG1TX2
JhtjqCx0XI1b5t37kfAupBax8dj380mjL3Of5Qg1LpIiQtI69pv1eILzutW+CD6fZ68p7R/oeCVO
AJs27nT4sqhOefbJ4cLmdjNhGZY43L/F7cjMNR4xeP/NClcRD2SzdGeRKlOpjswPiX2SvieADKtI
kvt8B9q8uBjY+lwfBagfUYqhzeb3WSB8NEPAwpbqTmamljcLEDIVYb87lGND2+Ksep3xnKzpl1As
ckYz2wdCRqBktQmayhy2UBnvVFrMAP9Dt7/Beq9OTU0ueK/pz4JRygZHv2L1h6SxCqUSjSC2L3jI
fDbdGrZhIDJZK+E0Dss7YSptBWPt+dw2cyNEPpVMrNujOhdNjOfOIpPaPNh2XNsA6vukCQthrfaY
ACCwLVODZDL6YeOfjUXulqNiR9s1AskL0ovRHR8lOCAj+YPs7B+gyq96UJ89krlkBAPdSco/UadI
9DydYwf1EO45RU+mQ/xUpaH1R+74dzG8+pZyskUjJ/3cYYyY2O6ipydBYj++gpriRHgkRQLQ9k+n
VDZd0ckQlCyQa4x24ZuJbQf0ezYThoA4R4Be4MqWQtq++M/1mdq3Ffd65HdYCix764B7SO78fuZM
ndKNxxaivGDDRf8i9ld1selPgVqU5TBNS94Fh120U9W6nsU5aXNMFk5jGCzsWfcqfDYtHyoOoodm
MGQGa5B1XNPP9if9KncxEt6GW2hjj2/SzQ6pD1JIyeLBm7pyQDuL0J+O+ihooJ6NTx4SN8dMIBOR
srQ/zYBvxyMWXY2tPkiVR+ozgOTOXoYYjnFY+FUjrYcRNm2BXMKqzUKIC/VcHjZ1Nqj8HvO7A0IL
LIvOfJ2uejAeWqIaVYpY5ZP/vPIKJRq3sJGAPDeF8WDFhJDXpOOj8l+AHByJK+RusmgwVFJ/8flU
tdhVWx9gQ5PhuNJ547OO57O52nr+uVbBwuoWtLTMeR308cV/35z9KClp2wGt/8ag8k7zKMo1Rqce
IKY8Pr1BnVmCO77K9YEj0dzqbJMqZDP+pqOTB2qci8CHJgOowjTF2AdDH2+Impyrnek/Vj+DUaQw
VwrEsQf5OAlj+SBspVGlXKVjUtkbEaN95HicOB4OqqieyvzmHy6bx0DdRBauuvpbg3K/9HM6oFwG
qO1ys2zIeYkAhLiVWwY1Ky/c+/WGqydu50Y7dWGC7oLJW2bTxVGMM3GOB1fnXmBKtonM5SzAMuqZ
umjvc9KnVGNSvO/P5JSay0k9vVwOB51AoadpsiRRHKovc9brcIrBW8V5KOOuVV3HPl5VGtIFqExr
ZAL4d0UrRaAEq2kKjiEkmvbhzQhavSsG7lxwbL5jXYasGlpcTsWj05vL68CAGGD+N1k+tLe5Fsqq
QthGCS4XMJFHMPTg/LfyLd0ypSl+cz82WmJMhH0X2w3H2bc71nDvBa0BUI2GMRshVthvON9nWWXy
EgiKfQSnOnPXZ/HhxHOXTOVGGwGuAf1PVltEplSFH6lsGFYPwoq9DibxS3/zsOJXlZX9CB0bdAue
iXRE5Zw7K3C/IWbs5D3EF74JRjCeOA96Q1U5nC8zUYR7AZ0q83xzTIc1bmEEuYcxNdg3ecwVGsUG
6VkrNGz+oqZnsutm0bVtIXOcFDQvEwLLxpdSZPM4NAY6wphqOiAE8fNAI1Zia9Y00lFLN/N9Jgsm
+xtlS65FmvrD/vro2cny0HMbmE0G0CD7Kk0QP4a/GwDj6vkennRp503xS27A5Xp+/ubZhQYe5AmK
MYOv95TqYHoir9joUKWcrpE00Fume2uzJETKfmNwvaA96R3JJeUZlDlLQxwv3fEsWe3uRkU0Dz9t
re+pxqJdv6SUgS1sydFN61XS0KE04mklLN/xferywQoo0aZfnCcLz41+UIdPVc7ez462GZ0DBjDQ
F+EJw0eOgQhZwoG/4xb5yh8V3AzBJvVT6D2uSRMLnPrh/ak9VNMcMlzhe5KQL9MplG2DRJCfqrzh
Th8VLAIHx7cY8IDVLtMrOEyyLzgaa4VQKyhHdOx/84Yalc0i+fQ0285IwqapsJAadJIjeNcvZQbM
bcc65I/7TCdN/YLG4/uEFh6SCbEtYU3gaSxDiI9kjy2GEWM6EREuyng95RvcciKH7CYfQZTSy2qp
9GIvBCGVAF3ZB2FuEJ1Otz+B5gegSCibcdCbW9i/DoY1ZZXQ5R67x5ixQwUcrUXv3BzlmJDXJ4Vt
cIlVEKcZF6jvZm35ZrvP4OF6M2tuDgk4iJHewltsFw3ESFOWfF042aWGXo2GmKAJL2FDCR+lC+u3
eU7vwMc5p5ZSJAoeu6TEtFh5yEcuXrbU+ZkNvANLc0UBf1RyWueAw04aXHYYZd7SLk3Are61+8tC
nAaKMip88CJ38CgQTMSkA9QYcNKBpALUw1gCkZJrNaxCucPDyALQxaP+qoTrons8svZ9Ys6JK33w
MKy5Q9cdgxk4DIfg3HluPEd2wQ6S9CLCyqY6Nkeq40GaiQiAzN23LPXz6z/7msVJrSChVo8wrirB
xYxPMb+GB+6nNoivFCzpTwtFLSp3hq0Y9osQFydoHGS7rT4ydCQcffl8fc3QTVWpd5/J53BbA7Bf
9w0cph+fX+ZuYTGhe7Qb228G9W0sJx8ZOdbx7dtZOIKHK5sjqisKaUfMPuk47oVmCibEBH0oEvup
f29MVj9aDwIDwiZwOGyp6FfGRLDol9j+zs9L52lkafQ4hxBsi31DUA1zzsGUg8w7oxOwxvwJLCNZ
XWWkVqgeSEKIGrvqNC3i7B1blpwFX9jNAo3AZdamHeDcGM1/kK1ZrnQ3uPJtsYEaHVBnJMEdtFii
EtPpC1IIqnM9r8w8kOLGw0hKbBlF5/MdyjmQUfrNTkRqiLvxyn250XC6mp4GKycdwPlG58foKyPu
FZaAwJH+DE5qFkExFmNgrlfnOuzHVGiL5MXDe3DCCR2lLYxpA6+2v3MbN/4+UihpJZEcmVWJM8ey
Z/1m7meNogteFafSiUjyfPj4j6AstxWdq156E4C0+i9gsB5LptCA7qpbWlY36g4zWyyzpo63pZ7N
M57KROSQSSAWG3Em+VEizNbgepu53gvqr3dFWpCCdCq/XHPaB/4krY53lCJO4cXfL3AOnyLYEvbE
9NuUN5byB82ZxpuiBsO5tFA9ULKtZtDrbiLQ0ZdSJy94twEJX0hRtCx06EXr9kVy5IrT3j2rltgO
xnrxL0bt3WGFrQSpG2kzPokGaqAP18QIpLDeEwKoghgz4aRIe6mdhDLXC+olw2QOcP+srzAYVDzG
HYeg9Kn327d0wuj9zDaehsHtFeTeSpkowwNjtWdD9m+GJsEE6PqEWXGM5mq87CFKy5uluOMLzGNK
1WmMGY+P3GlczJfVwrC9Ndyw6Yqt3fjfJF690mcfABk3ZtoLzUy2MUivK3bYx1N08d/mvuG9i3Mo
vnbCeBHiye45siuSnD3nD4UjjPAbAuOM68WWc4adfV013MwPO8SPt6q4WaeMxv3jT3mptqkbs55t
5BS16ML8iuShw9hPZ1f9V1qU/PcQIadgzcBzWIPBrT9jqYge+X17UHMm9Fwgotz/TpcDiKlF0BW3
DVMLl+LedhFaWJsdCzvRw5FBM51lOp4+giN3iL+dE2WFHs5NG7QoVzaGbHRy3eIdzOLXLoJQuBia
raFBROF9R81rORBAYcgKkhm+2pRxF5ivzYVEDQ+8s5y5OEYFmBR1u9cG4UyfaBWpQ5co0Rx08Vxr
bIPjSVAd9PDWcaZWFMajs5EthZay7iEqVDnX5oGtMQnvmnOHtgpdkhRpAoVpcaB70vv9bRVz/udV
G9xGb2E+vO+ojv1cDMEGA7UwcH/XY2LZeZLOyE7/gBe6Bsth5WshmAHZQ+XPtXoPt2IicxzHc/Ep
VWFnIDHa9J4wVmYvYuaX6f8XpJtyJEwrgzaA6qaMyxemN9eXVI0kiIttWFcHUXkCwg7cWIgW+fHI
lmpVKURxDhB9MITiJmwBcrlult1lJk6hWbzxGaX/wElAvd/UtfJkNcZ2PFc/DKMAmQi7thPdIIh9
LVW3h1UKRPWou3UTeK6Qvs9dFjzmCUSsH8R4wSD3DpvGdQPlmDtHH3/3xkPHO3o92C4Pu8jIFQ81
8+AT0QcTKkRfYdaiZJKNagIOdOAt/jDxPnxUaBHqLEv0GY3OAmwvskxKnCu4UcSw+ODb6VhQ0gUa
tS6D42waVQ8lm5FXB5k1kTy6nxTICvDFE6j6tGNnuPZ8oKRryHbCc3k/J3nOg/vAusRc2JSnkeeE
jDly3w1J7vXx19Ab+7GxkLPmio1K6KfWS1Qz3Ed/4apKXWRBmigTHUZ1Ij71OJmdri/YPVJQ4+PJ
Mzm29LsLrJZ7scak103IKI8aGPnhuo3m/4Qg7MI4pB+seFJE2qcu4fwvAzVHj0+JIZSDI9hhdhIT
TQJAymts7Z0k/2xut1Rc/+aioXhOIuGEumH4lSS5g1nC3215SmimptpLXvZqAOX9Kg0S3XM4rgAM
/32ooSLsGOYQycTaSThT/zPs0hwj4J/xJxg1Oblg0xzJ6Jq2ow/+8///btRx0CXXKYaCp+QCRDzh
Wqlzakjlho+eGfJ1MbjHZE91FyBT15G9r4VJwggtRALa2aT9LGPOp8F5Ai4ReZ2lPM46d6Waclbv
P8M/dyKyW/gvWkaPvhr2AosFcbEjoirQH+exn+5gS0vHrRfYfHSS4rrzLzHlwv6wt1GAEViJawaa
LiJOt8LaKN7c8rs7lUT4fVASHdjcSshPywa9wbfGmHl5ysamKuHNeTKYf8qf+t02L933y/O8EOpI
akGLBUNVSsDLDWwxnHQDkVL4M+p5LfnUGffjB57Dz3MsLYMxPuCB3SaL6hydVHHbmcXRBCL+X8QC
XKEgYAi/EE23REqodVdJa+6mpjllf+BYPwriDrc6Fh6xjdLRMiSkA9VB9ZBuoNcXrrrERdhvQBWW
lrkJ7broMi13HE4hAsjnBHDiq5AkGcG0ssVAKQvSzFvUFnLYVJGVX5AxkTBDum/eM8nZjHrY5uPn
WEhm+kMCePmwqh0rer50NBNN5eqxIlPcvMUtWmzx6W9WKErNvY8Y5GtleULyzOsp/xuAKwjGcRD3
AyltdJorgtdLF6Rmua3h8pZnhO6vb9hGeyrgssn/twjTn26e3OdZTsQAegTbQUByqjP3sLSYuQ9N
WHbtihkfgYVn8izibKqWZrbEA7CPjBeWL9l44j7S1QZZ6pEtd5TPHb5Gg1+uo09pIoE5lNERV2Uq
V/rh+8sGw1n/9VeG+qYuV/z5U7izM1IVoXLP1LJvfyR/5t+rncXetCUvzgDMxRtStH6AGeE8GbVg
2IGoEmlSBwnqVg0AFrcsk4i7eFgr5bo3y33yfq4hPsTNWb6d7gjZea0Bk7i+VGcyFXvfZ0NjRqKv
YWH4XHzv1tSU9mguK1DwalW2GVvWToK7mdJNloILFOASxh5rnn72ZJYoosTnMu2DOiXTytGFvQqt
Um7VHRU1IDG0njmYuTM5caOSAyxjxWuQilk/XGxUzbaDQJ9G3BxR8AeZQvhzJo+qjodqTAdDTIMq
HVTdf7SvB8UpAVc5YLP73MHKIGL89zSNExKauifunaOji8tQOWHhlyiDkGG40KLlmlgrimCOwoNK
/qSw4PI0/21UZKNW7ngj9OgkbIpgAFaofoE1GGQOWtQzFSaVad5uD85xr7rHogq6D0wseoDDtuuw
9/SacIA/Qv3bbsS+MfxIkq0CHNIypcMTTW50l8QDvinvF0GgE3Q0kgvVLdYbHxl6Gj1iGQPmahLw
Tauzjjf4kaaItpuyNe7LEpHuTAI+oUs5B3fGe8yFjLVDt0+s9oIWImUS6YHjglAeQXZnsKFUJ88t
sTQsG2mmwQMVGYx/JwV9i5A7yniaMHfzmSb1r6Dal4OZnKmGN0eui/mul4haaAefOKiCB7ZottMi
6jA7JUiXZDCVf4S6GUb9obzuD3XNkWPjZlcK97ap4bxIJ4+jV9HtbERJ6aaRAJ6DjMaQOlNOtnU0
jPexgTZa4jJjJtHBh9ieKg5OO8opVEIDmyjPcdFB+82bzT9BzqzH2hrqgN73gSTTX+2KUcMcueVc
pyKIW9N1/BAGK+MdZbFG9DaOM5cldpy5DkabIHRBdFwCIybfJDYU4MgEsdluGaSbRQhWlIKvK/sx
SSRSCEfM4kNYfffcTL6YLQjNbN3TQYTG/ekwyufEpfVmv8EamhRqwRRJ8yoO3udKUr8CbPPwlGBf
EX0sRcTONr7efMBJYjpc1O7qtWTjGHneMEZ23VBS8J/jYoFDiGyjocLG6/hVJqmUk4z+FgJizdNF
Ybqag/d1XK/DDUf074x8dYcGrYUFzjhAGFAnzXTyB7EZTBRwHtJn7eNYXuZ+6uP5831PAfCXNECd
8SO2EP3oXA8uUDDdXAl2owrEW64p5X1bK6I23OtOtrfZ1xMxh/J52lcTsOfnh30k3df2xAVc9MVy
RjlgWiyQNoroBJfRkPBrQO0WTNwbMrZ//OTurVcVn41867SDEY95udQA8TiPRfLI3Q85AUnEYK8+
6ojiDbzYVIzk9VlpHdtOL1GDfaOue4faRhiFRDm6oMvY43Ykp3YIpqYqbZ3qNT8gqgCOIyAJUURi
yOMLwsJRPZNXtXxQn1XMbJIBQeJi3RwUZbTR1itUhYLieKZZyuoE+15fB/Ob8ZxHbU9QgHxPX/PR
6516q854x76XLZkKK05DOZoDI74BWmGczNwOxWeqn5V6RcO79TrMmd/JVQE7ViaipyDvI1Jtt9JZ
b3N+R0zyTfMzRXioZQ/7OKuK/w5x5VPAnVRdQtr6CqrEi+F8Lqi2LKwv5HuSWEmitk0I4ogWpDPR
FNWbRnZzujtnp/fHpVL6eg2hxq5rHwGiveaqBQ8MZI4XZh75kskN3XfcG7m+cHbojKO0uuSxCgZC
wbqYu7bbFn+7+yOic+HXb6Z9R3xVYXg+Pn2LBBV+FrZZScxZ++WZey+JWDJ1l6muuKf0RVVPfuge
4vC1B6bHNL2bsIUHnGIzF5UD6MZbB31W6pUSnGMif5mIxjR4mtoXdnwFmNdlVuDxB0GlqlhY94xq
+FRk38kx4UatZcpxGnjQnYAUz4+NzIO0ZO24i3vzEOW/YLjRcBB3YRWN8XB365iYiTjcE36gtyFH
ZBszlw5J+JWneDQ8cF3apLB8aKrnc6Iv/Fund1gIuEFrMdlzHF3ixa4mGqHwFP/pswAQNxzeiZPG
fivULrZm10uOCynT2s/cJt0JE0/QgRV79Qd25NBuhPbP+nEFVRqw+lSvFElQ1dEkC8icNPQtmuHY
pMOZvN3EbdKVnL5j3FHX9MOANrlxLJfNEUJbaAsyY8oZ0CJvZnf9466K1fMpZMOTIAboe7miQkpR
QRT5VFd6EZWwTSR/M70CcKPeuTTENaVZesFXbCjO2OrqDyPxmR44I9cgOwnykMg3a+S90KNHTAVo
ow032kf/dxM1B7ram5IR4RtKxA40n6xDWk4UhNRsOBzB0QBYZ+/D+w4kxSbGhqKLu67cAP22j4Yp
+kICLsWpoLURKrIXKckdn3d1FARl4B+I1MmOYm7winfKntqJiOyA0TRQE7v6eoNPzZ7tSJNZsBL7
DDqGCEpn3Zvzp4iHjkkYzrtmM43DKfU47+z3SuoJpwNk+D6j70yf4kI+rs7dDXx5FjHYioeDavk6
Y78nmLXPP37eR39qIhQ0hQahIMn5+H2TWzDib/SFivsl/1bvbQjyVrCv5wSYSnIdxixK871xSPlk
a82SWF3y7TOOBRHpkFaYUIW1mA28ow+uMbFFF77N5xPtdK70Sz7+yjopYnSiIv2+9t4vMTUGsOjl
ktjuZmlrAB1Qs/QtOMRZDJrQKAnunp2aRzKw/VEQT3pLIxu/YCHwwoICpDyynTJ/oUYRsyS/ew2e
+FfX0hzpB/3ROurNbJoQ/f51QcpE7BuDAeW/NmDLh7v39JY8u1BC7ym+2hxzv/rj8XfLwqOvhnE8
RwKRi/Rtq9jrz19RY1+XTZyWpbBF8S09nOW37eAJ9ijP5gJg+3Bkf2dMw7hCPxJ8KXwMa4oc9Avv
jNcI+24wXVKod2b1KhgEZFl5iNYJTU310v69mB/U2o7WXIDO/N8NNPLtE8sC9IESNL3pB+2Wes1d
9dTIFN7z1+MBXDDwOXZN5k2DZfLVJvPd9sPmVoft+0XBYqlAIFGcRKnfTt+B86Ipqt9AxlKerQ22
KnzX8ySWEfuyEaHCExxhzsLWZEB8nPf1PeZY3aekY1ASuYPNWux6jDcDX3pEQT6GpExeZwrMaZzU
BsSPSFUE/L9374Su+tMYeJKXYO3cU3zJcHcVUORcpsgg7cHsb7bYivatR2hbu2rM56Aprr9fh7UF
WJF3VC3k/Bw4kSqjTB3Styt8/A2+XM5GKMChnYzr4DEAJMmI2hrobDMxV8Ps4jkpuNAoqe4m4NtQ
Hjkr8SPdysC1tO8mp39Gu5D0qfiwUUzuBlEboUSQMRJOy8HCHesRbbCD8OqniKCgmbqc2HvttcCy
WdyO47hUJoitcI7gLw8qz5CIlM0+iegNooVViikXX6iDmKBr7ZMQrP1oNF0+nSduZdIR6wpIYRNE
EnRf/zafQGkG4FGqkL2hcwUhJjYB/mljFqsUO0kYJv2cC25WRxE0e6uWbjdzFvF2goAqhCSWMt86
SPBeFpS1C294cPS26tRVzPPStqH2Z0TdOUx7PrgiwFoOgKTslse+ogaSIBk1gngJOolL3bxw/H6h
QYcQGnyMk/Vm4mv/0WY6dXs99+9PXHHhjakRK4NyiOrQ4+c/hz/Ta0prY18jS7Qt/HrbVmCWbwC2
NpZOegq35QVXl425jR9lG346Ja8C9ezX8nZ3n32ORbxP7mkpdv1AQ0TppBYXgo4ca52HdLXSAeK/
nGgzQkTnVo+4LuwJEriUQpfaiC8NzHsGYh0REYORaO6SzjE6t1vBvJFyxHMSpAOCPFK/omQzeqGV
rjVw1KQX7QgGQVDNx/qHT3X1LO94IrWEl9en/IA4OqlyKD5X4F375TONIB0WGCSSnhIIP9FYgzWr
cfADSLEZ9TTiAhGQX38w01FRZl8qQJntdoJ5+QLvNYVxQDdYmotslSACeEFI30D4y/FY96/96lvS
U1iLc8BK6mIP60GfAGQqfLx6M65+9whLyL13gotwNR9vjhMvtaBnjshjfs4+ybvAocj23f2B9GIa
QI93DBOhIdGk5Czt12I8Vc1x98ZwaLAA20p6T8h26MkKLUD/LmZMHc6jBvMfxfCNxBaHvriK4+A5
qVdyNxGmVHzbbsfalYxy9FcWPpADnpW4VK6Iq+CDw1Pp+RtlbwxvoL+0qVdQSN92DGsa8s+QtLIo
PnEqeq6fUsy38fq6ZK9LPWrMRgRGrXC20WBNGuKFIPJacmHaXU2pFJtg0nDiO4PWQOJG1szOtlLX
gp3mjn6kiIYzrGrpwHn2QxocTiqpyuCbBtedk/gYFV06DkvoK9+8xZZefK9Tvgl5ao+nLW81ATil
U3vWI0qWR+SHEq78ytNYn+FsIegM7+7RTuSlshgGv1XPSfpvYZiuTK8UrGQjP2TecwywA0PuE+xi
KUjeU9Syx5t+0aMvHG0HIFA7QjmC31jyWVTtk3dgJbmLnPG+scDgvgcjQbzQPhMy85PxwcKo9zEP
v7B4+YZww62KH0rsVm/GrELsV/I+L/qSJaDmsWEwruG4drKoYtz+FozXQ4DJE+UxHnReMw9BrUQ4
VrHCEvWlateruB4hAKltkpoX5MZra9LU8fqDqpFZRWLDlQTF1nDoZ03riPMlw8+m2L8HjkjZCnvh
0Ka3RmQ9CsgwYCr+RRMOM276Q1BU8+6s/DHywqC/Xr+LucwWPVPM+K/283a1ZQP/Pjqzd5Qde5W6
wVpfvAbUJcAu3KjwTKypGJ4M3Kmrbj/K3QRO/NK2YFwv0tCTsESEcjyTbxagII6FZb8vV9+Wxcrc
xsFmX+bDiM6l7IFOc9AiyMqwQIdWiuiM8PcZ7Vq3Iq4v8+TvJ2j8NYuXJIvTEQyjEvmtUnN++fGJ
pxoJ/hdXRhL4gOVbDTjWvdONiq5PLR4r6D8av27CcP9RRyrsFrVR1tEJxERiMonwePQ7C4SUxWlg
guqkgWCTWPljfoYmA+8qpEjP1hMWwdUfOlwYuLcKudq9wbcd2nMuh1zSlvcSu7ZmoloG1JCjHry4
ur5swQmvNWZXkE3m2NpSzyO5yfAziGYMrP9wyBIKmCRx/4t4t/xn+G/FHFVeXAxHTNzXOLl7Ayzc
qei9UXy9N1EtiasIj0BgJ/rPzJi+mZQeN/X28xDfrlxWtIyOqXf3i/Ee2peHXdRmJ00kxcKXR3TQ
g1x9s4pjYWgjfVSbkq/ZTPq5ApjTt6Pxbak2FuD8AvFl5s04MM6ex+SXGQ+qEdNPEGchHSiWJdyS
b+YMCloiGW2Ry03rMtZjzN/OeKqlCBj9NusfjzEg731q2sT+/Q+6UjmBX3cfvh6qw6nGozE07sHe
ac4dsEn1Qlx4uJqeWEsb7LfXkra5PBb630cOn5KLaH5blSECtHKA4aIXvX3mZRtRPX5B2CySgUpt
9JpPhncs4NYipV3BgnPNheOqFSUlGegu77LFd7EwjmIB8EZtvcGM+fRUL57Uz6Ib+8V0L+AMOFVc
RZ6CJgoBjoiiCIpRJXk/gp4ZuUKDJ59UJESpYh8JEXUAjo+SJBSIx/iiTh3si6gtwLClbFQ5AF4s
GapdC1tA27dmhDLSmYcAe+vnllkjdcWkcNF1251CP11AwOAYcIsp/BA5FcNzktcB47aHgSLdv1b3
COd3MBSqP7bW4fF7zcmhAlZ4wlqUin2sMg4ufoeQo6iN45WJZw5rCDTyk0xNADCdHQ2j+KrOhrio
X9LByMAKHfktGxXVRFChhHPcMy7AS+3o24d76qndtChQYoiVzaKx3eDnUilYZM/8Yo0CWUHOlGwO
+AWJ1ZrYKBYZlaaWY4iZ5swWsOHsKklePi2r/TveqPUgQm8erLH6bD2XvdUKvVECImDiCVM4Fqcu
t3m+7FJ+toFPSJkrHR/HwSzD+pREb4Os+IJ06S9zFO7vfOISUcRAGwfcQGMqaqd9V8bPTtn7cZAu
T5lWpTKezU8vxJ/QW377Lfz+TRh+U3YtGETzt8+bCXXXofTQeSd0lHBhL3WgPvhq77BP+5o0eTB5
Juba30dmcSB7PYb8CYVwk5bNCRSLg7ejgFACdYRhTswn2TCZYXUVTcDaUKAMJFe7ONdnEalScMSR
c5YTyP20MdLOJPzJyQkrcUAdUT2CbMoBWV6Vocoxr9pCvSpkl6FgWOBBsiHPTUz6/+Wm1p3ioLbL
+E4vatAtHoiTsKlyZxgq7cQYqMwWAEVAJ5JwRptiI87uMMYjdTRpCcDLwE9OD6jPsjFodYJhq0os
cfplKHAXkbx7dlmrsEdLLrUxsb/LlzI8E5VqtMgp5pG0paxpgp/sEblR0pRNsadjGLg9xMm/5Zdw
4zjGHqg7Hqg7bOL3FJ808UIGecYbagQuSAiIhJg78UF6xqYjAIWD6XK6CVml21jCoIooJw6Ad9Na
ta3i8xJnHhzF2cuPdpqzajymzcAqZpUp/sfi4wREL9KkYR3+5UrkowkxtArNWKVoC+zz1jn4ov6r
WYq23bK3BAz4frrjnFdnj/IJ7gdTkrJLkuKYgF2vL/SM5MCjCYjLpUNeG0CTFoSbnYC6P++5eZ+q
W6YAkMT1Fau9gHVrHCiR+DuSm0KP6l/XHXSbHOj5N1Cbpra3kEUMcQ/Cqpe+M5FK7ErmUBFO+g+2
EI3+XIsNq6Tn5zLK+ya6BTy0KuDUc7O8H6rSj2JSNBXyrcm/5Knf4ahaG49FChlbu39wM21IyFc0
RZX5k/kmBJPQ6mYMuQGAJSkhDP/ONRI+t0RuofQsnEzWriBulwWn6AVPBZzpUMaAOB8RneNQvM5t
1QRKVD1mx5zHqoxVaXqHh3sJZLqbVNsOhhmOTzcNVFTNAzwCdZIILbKtIcCn+4pPWHHBAuG99dem
u/w3reSPAJr+MPhVOPa60b6nZFl6HDlJ5wnCzwIWFDKylhjTFNPGJJMm83Edyev6/obriwBW74M2
BL2FLNRluLwpjnnd+2JK5Ra6bG2mgqSum/A8yKk9QjEC7qzf6a1gp0m+vqGiCKvIise8/Jr90wuQ
aBEzWDz4so2PG7tqc3cR4Tw+iAmaBUvJ0QiXBk1ZiTyejlgk9+C2DYRQalChAza/LIe6HA886VB4
MNpUHhODaSsqgWtZZ38zhb2iPVkXJiYeXZiWSvPKotJ2C85bDNSXKK+TzcoJrZbHW4gxNr8CtvIK
rhmggHXxOPMGNVaJup3m7SXDaJ9mCFUi6V2VYFrcNDmHAv7imeaTQWbBWi/NTfqL3E4f4Wpo4whP
Cu8i4gRdGtRRWuwrz/Tfk1UXLBHzbARtlzBx7VV6+LrmfmZK97vjejUIqOmL+VO2HgIkD0vUUpnX
sjYjvI6AuIw1el6AmdfWEdU1g1kxaZTsd60yofubPPXoZquNLfByC5ekYZ4kW9vmSUQS+xQDfkRC
E5FuBdjbVOSpgKcimpcl//o+q+FtZQfEskprqM2c630xx738I6bkp0hEg7eMP+wvtAYdjsIKyn66
a9+fJR74iS5koEs1AIlRj+567M/xH0fDZZxmvjFJdqYRP7GTP3LI93h3V3ko/1J9WapWC/DhIGUe
/R/oKkTqqewAbstsqzpW7jd6czzdB1PkfPy8TrWequD9OIk5lD0qfUYZsuXFxSkfj5ncd96N6n3v
0WSwd8IffLdrSU5WdGec5zmTfIF3lHh1GkoYK5qiOcIFjqGHtwF8xlQKvB9rLOWdMdirP5srDT/A
4acRDSahM1XfLnovZ6Us0lLEf2mGRv9PuNA52OWmeZwqey+b7zSSt/ZXEBe9T6Mwk8DTNqK23bmj
opULw2D7XOAZOo41WJJ3Bals9dsOmvUKFVHTesR3VC/7mNM3TrkdxsDVGqwoikDAZ9FKYtaXm890
jlzXYUb7bUSHONXiQ6DeiN5892bx9JND3NeYWzqPj/JLU+FWw7xUwMcvZ+WVTnaNtx0VP8Pw6JOn
8/zqbRR76OmBYXSXTiA0wiMJivHGYCWw6iQlEXIUK4v6Kcg1xMkfKu0kRcDAi43UxerqSB62n0VA
6LRODevjp/2o/N4ZEoQGJA9Ic3tIOepOaHheioQNMDlneYNxV41plCgwwrC6TchxGOEyN43k6S4x
ZZ0Uiya+8Dx/F5+nMPwBlZD673RgL0A4DS16dvYZjjUWp/8po+VDkDdMBZmcs+2+luM/RcOTUzyW
ouYJPre59Yzuxs24yFwM2oZpcsOeTJV6lg0ixPze1aheClsY4KMm+occU7DBMPqdts6s85TR4eCb
nw4softbFSdpBs0mpIeusKvxHC2VvRJc39WXSFWBh6BAAVGqlj8CFMtjnfGYGfQP5CkWwGEsHqsW
XTWmm5A6pt2w+lsQdE7uyCMexDSodE85UXAVQ+tUinaiYAs5deoErfHUfBGd20yhlTAL4t3/fMKi
3A3rbKR7bzNX2QAyf0h+dKC4FKcnXlXDRJYNsyK8y1ilkHWk9Fwkpfkl2vmAMUD+Vx2Lda6iVZ97
31/OeITujc737xR4yQzOdjjPJ6x534dEOluTCGFqTNDpaSNeiRIT8B6VQ/vD1cKjBR/RBg5SdEO4
xn6k6VwkWWFktOBCbJPYYqQ3SSZZJgROgdn0IeTc/UR8b5+jgJlQV2wqtcecpnb8DKrRHGJPZbY5
r7kU+ZbeMOUwv4i2nx19AgBRJnZkxEhvelBzEmZIAW0hiUKy6Iz2RAgXeH1k7k9+Gunoj5U5OVw+
sgmvpa6LhQAXyP+3BTLlw5gSxma2qxSvnBV7Unca0KxFQe3/LkjwE/oQg6cwYXAQIaWljeQNBNuf
ttAIicrxQQshZWlLGHu4leh2VVTa4whHrk3Hefff/8IWGHah++bzlLSQS23Bhe4MYkGDbmz+wOjT
zsnDmn4UVxZ5vmxK2y9+bYusiW0/9VflXYs5NP+Jv45ZX9z1Cw35uUD67b/Yq+sfe/yVMUvj/opM
xJTR+kXvn02F4u995EU18Fd9+jH1E8ezYRcMjMzbwOwWR4dR3u0ubvv0eEsha1r1o143gMD3oxDj
M5Py/GI8MAmKi5Lj7vjBEocSZIIDCPNvag4Xw0qc+N5sL6ajP3O5DY57I2+PwieU4UggYwMJhqSr
tGjL8M7q9VdX4G+2JOCh5vMdNhfo2oMFF6VA4sKD7tqQcj3v9Vf2SDwRwiCquSiLp5BWhsv7EOaG
zkUYiaLlg5X+jNShNHFmKySV+FOUMNxwbmglj/yc+ncYO726O3uJL6tq3e6xr0uEhmHFjo74pSuv
Uwll4H+XCQ4OZ0UX7yFjbv6wEIl2DFWkRa56euPZ6jKnM5lSx1OvnXmh1WF6GuLkGe8hvYu99EK/
NFYB89KssVPhSALuWcU3Tv5mgTJk/cdL6VWc0K5SkzoWaAAw511CKSp/8SanICjbC+eW1AH0tzhX
ptqOhQdXyIfhfjT1iMdkJ0LaLVLyFgW2XAif+fNVCs/+/2sQZpG5sjge2OSvCf00XaeU4eFntVYG
N52MBhmSTXQhbCeRtm24Hy/g57ESREgOVCL0zrFSTkB/DyRAjrmpTx7uYVurHWbR+zr6jUmzUhTC
VCTidGxvJubrbQUw6PhhMwfKEVet4n8GmRdxIGWEumGsuM9D89ZJ5UFcqi9VPF6pmoqVQ99YcwbI
6AayZMKDwAOv41wa8lX5AY53eCkU9Dbv0DBFLgXmbN3ly0oucxR1Ia3AlDLA6HbWVGxdHmKZDokA
d9DxDQfpnz2sRU4NHwvcRJnhkD29p9E2eLGOwBYJE0yeq1TWO5ILgvSt636ysaoTf+jTRB5uYApL
acgTSN7RCnLHUcPNWAuEDKgUuhn5DFsag8OX7NI64E4NLgPkTdfC8S2X3IyXh+tkWMWmnn0/9Aib
VDChsPNQWGZy6ro/n0ngneODOC8VJ1Sp5FZxParsuOyeGB33rcicRJa+rXmzkTcO/R6d16z8jLrb
YqR4rn3eHeLc2MimnH4E2KR49KINRe2WMMzCdCEDnQdLtP+aU8m8agWQzTfY4VP8hB0B1r7cSS99
+qAUrG5cv4aI6wnQqkyuxm47o6QW8oCAR3ctACdNsSgzFNhdbLNn7hlXxPWJI7xcV3ixe40e3m55
gXfNpsk09odWxsjrXjgF3qCiEyT8x+KypPucj8fZdwvmlr7lnBbofqwIgSwUN2e+Ocj/9HZxbwj8
xN0QLkdVHMJbG+1vYbNBa+LF9IGlyEEO4GXZP286I5LsVMoXTUC/hi6eh2E3ESLnBphdC3HoKXoC
9Kd27ORW3Wt/SzPwrdQpLTcdDnfC8ykuqYwjhKL8vagOjYLk1uk2j6NmmSnK8zjsnZwFG+U2Ydje
QlCNv4NpXwvHg23ZRGFI6hw6lCNyESrcs56Sz5DtRkLFUWbhXAEJ0LYl/e5zGdlZ38auvEtHxQUJ
433eY9OR+edONtp6M0htph3d5moFHGrb3pevG8+52U7b3A1EQFLT+UP0fQtKGLblLwBnrHhGecEy
JFrZ2dFLTNFf+L8uTyq7q55d/Y2q3IW6POmNCGQhjrrWgNoXz1DGKiLpEzzbIKRuxA9zuCJbGUXl
g8yWuRH49vOVo1U9gqoW1CcHjDOeuKaWloIiyDskd5bnWJN/8LHaBsXA9N8Z2blzc8eojbIhE3if
2Qq2WXZ/zNcO+4FWldmH2zPGhbYloencloWh30fnUBu9EivymjhljA2UpVlSKE/Zjw2Eb58TUpRz
wCtlbiPHfJrQttXmcTNG7vgI5m0uv46+vymQLQij/7WH7rjKiY+Ctv/fV+Xy0B6M7NHghwuJcJ6e
MCEp1+o3sAvp4HjgQMM9aFUfEyaPHBYm3AElWwHyScllaA60JLIip08YszkSa5/4ByKx8ecA+nST
0kNnTAbM8xP4xj2jz77ZBGePigTSyKU0d4F/oxehtVUCZ/tpWNPXMSiy4Y/1N1pinWzBfCLuP7s2
qTFEiKT6ysjVQAj5WF1IC7Fg8jddO45Mz2/WgwUBuqV5/XGYWkkJRusRa0LVYG0URkFZxi7EXTBk
DG09Vwr/8JXzSNGN+wcwz62uk2M+RTAaYjF2+uuEvNRHu12FV0IT7nKsM9vojlLUjaavA9AgoHYg
GUrExkqpjXKeTVTW5bk6ZF6e6fvZ44k2AEPxa0q8KyCQIJs+xLR/yBP8IVTEetrHaIym8w5CLn/q
sNiKU7OGhrPVsg1r3+/LBYhhdn5ytCGq1tvX8mNIYjl7XoyTJvkUSCi8+GGtEfi8jZQR8JYEkIwZ
SkQPxfe08SUyktHvtNYbRQkCIK2xOkLQ2n92MuaQT8PYp0XJiswLGJZdpxIjfiYxtZykreAzblX1
H28jTnyfZ+C8oOc6Rmv8CG8f7f4e6IpVQiLUXUr/lllo7j9L3UXQdtnpTmGwAxFO7kRTg7M2JLJ3
pTD5H1CMaupUSQ7EFsXaN23QsaKCX5qYuqDFFYzfXAkIqj7h+ikG3Qvqh9gjoaIucd5GboVBrby2
MqrCKxuLHy8Fo1NS3Bb8OOgkf3El+087vmpZQu0qtAChEWvf4aKrviwzm5UsCyrUxJd3NpJhhcfY
oYpSPchUjH/9ti6vIJoJ9My0Z9051hBZBjqLXWGUZHtCsDx3oOeHbJwV5BHODVSgbNCOgFxJeXOi
eGqjsRflEtklq42voVt1rbiAm8Uj4hKJsl0nGmsd/JMOQoOuVQ591jQASQkhtj4O3r5Aw+5ae3fb
8jUcv36RzS77PorWXzZh3je9XccJmuNUh8o3i44YXkP0lWaWhi50RmcRer+x8vywwN70Yo6mDSWh
79XHGPhL5HgSwKbG4JS4/xAcw8YTzVKAfHwWinDgCElwveBi5v8VmxBKLyWKjwJHOeLsMCYcpU+O
UBRo7xdsrapzpsd3vVl0If3HosDkMxcxynkp5qo6h9slZYsjxwvp4s/N5Wdl5I7nSb+LDLBZUoZW
Zg13f1hTlwvMg4vvycVJSGJHSz9+emwO9hli5GsOZHlxQ0CtQujSzqSZihwupSZoTmKq0IZdpwlz
bHzyHdGYeyb+zvpMhvTcz0ijCYie2DHTqZPDw49Hq5MzGU5mSTWoMQ+itHZeaoAZ9iL75dk+50/e
cbU7Bgf2fFhCknJ2/TzxJnY8YkBJYF8noA4DtW8ySQbfI4UEruBek4XKnE/XIDDy+NvBr1kdVkaU
8xSApcMU5yCkbuiggRQY2ggsh58ey23/9QU3omXu/JxQTStgri0UhLrqz/U+SgdKJGMEqYex+nZh
uJ430oQdpHGWaxDBRWcQXuIu3krWT95ZpUIoOn2vVeR01MQCpefNxdVTmptY3E7U8WRQzpXyINUq
7Piptq0dIR9QVIjZp3dDsGR9PHMuWF5Okpvy2enlrikkVl7k0rVD4oaQL+qAfZXUJCyS2N6GtJQW
ENFH6bCFcrC+4lLDxUjhloSJIFqJaQGdMipD+ho18IaBxcUqsFSUUvsSfH/v6HK5ZDRLctbyKfcb
+BGUp2D/Zh1TYLzag/7KZu9nPx0nCf3neVALlOO1qqp1yWujc+OrYTP+AbpLbkQ2SiKSg6dEGrGD
Rlmbt56QwQsDl33/VQMQMtZ8PbLDNyVVw9zyfN56xKVIJ7WHEg6DNsigtIA8N9fyPrzo61v3AQxi
jJYOIkyJyXQToxQPD7YeezslnKVtde2JrLCW6GRYn8XKucUFT9bt3wthmdAoOGNZmACFV3lhZ8Nw
KckzkeDeuPap6vKnLb2HVhV89ASYvTSEAU6qgEK2N3gM05ZywVYbclIg6qNRtN8ld7fgBK9vi28Y
7G0X37hsQ0vkoICkuUN2ZjxvjhtZGuelDBMbZgOk53U/dlaGMPxWLL4/LsNfOwp7LzLuq4pOIp3d
lboYNEMrp2aPNslwxEV+y4pbuAzp9jS1iQ4rlayqI4w+ltQOnN+1fzVgGY7SYWePSUjvhkohUmbe
h5CetOXgBPdeL7Aj03zD1mhWPGdulw0pkEouflQ0pDlHhj6u3VN+mMsGfldc5a00UTDl3BeBGHLl
qBqAY7EjwDRBgxMhEed6cZSkSeShruHnsKZ1haeQnZHlqr4s/oQ7ikFbfDTLjC+yWwBdq6EjXE8O
E/f9nmAStdw+3fP82JDWYQe5UgwY3iAkK0PojygO3K40sGBhhZF2ZVYD3nt2O+YBUSbWP0uM9Wvg
Jr76LogWygD+V/Tqc3JsdzOg9z2Xvf+pnPT8/QHDcNfKmNktFdQAzc1cT53pCTAm7pxgEzvsGfkP
LfYOpo1yNJENRNgKNr3mpAmozt5HJ0BZvd63dByarlhNmhR5vwON1PyP9gqtr2zAJFSKyK2JQ3s4
O9jUkGGQEzBL52mfPnJNplUt7NvOEIG8Dz8gKN1vQZ81vNsyLTZbE9ut3N0Oq998Znp+NIHxB+pm
F/9Ur4jlX6sMBtulMAI4hX55A75xC8iw250VQE04+LF8rn6K12In34KFVYLAzkjL/eLZkpOXN0e6
bBUoAQW5gRcfoYlzw0rpzoMw2Id76OpFEhXAVR5JqViZRNpmhEV0NlqlGq56o/U6J62lhwtR5FR4
kzdB0Mx9SnP9DyhtIjgicvppwoilNDrEjYfkP0EQ5+AlIqfVRguMcRUd9NXOl0wbt1V37Amn1QGb
O0NcU/bqNR8SiPbvlPd9HC8nR6Ku/zQcpJlUZDETHzfpeiwdhgUqNY5FpxORin5xfykoOh1KvXr5
mLBj6y4F/ABO2g849manL7UimmGSQkE1mupBIrN8xZz8ywrc+gb6riuT5ttD9KadmImvRzhWew7I
TWbLKCIRWkhfrMdG3wq6TolwE/fi9W9zkLpgmFMlVOpK/BPWIWr3zUJTXOMBaAPqIRDywgeERdE5
DGyiWm7cRU0PRDWf6HQ0T/nyIOkx20F4nLgbIQMUdv7RerAsVzr+TjZ2TZ8r9vzYYZ0zitTGu3sn
QxShPXIflL4FDsQNfdNOQo+kvYp9/qFx/xv6lrdyiMYej10vu8xDORxFgM2whGbeJZLYlXoLZTVq
2MjWJ87rKtedQwewRSB3L0cTBv7cwK6p+Y8GhNo8fCX+NniPunI0ZIJBm459bkjFJUnVaNwHx43j
BgQDVdtcpLICnSxvPPGsN06TVAU4+vidHfMdJ4lGVpP5RHaIjEBb4Dy+1rsYAnIojcZw5nz0Mg6O
MPbn+1lt55aR8/MD7HXslNmoITM6NjjwvD9C+dQAu2tZWQICMZEklQnak16k44JPFkkbC/ayR2Zm
xnLKE+EWLINcB1/Uk1wPr7/Zd4Yj4fkKc1hdYihdsPkmChENn/3Gc3mDwP3gq+FWq5AkxOIjbbXG
U3pOf8+6pNVr1odUUvBvG9GlokPsp2oNNpAih0k7TaezCxJv92dRKz2Wc56v7iqJUSL43pe3otNW
m/70eWh3JHPeL4j4drlyyFVeyeBB8vqADSQ4Fl3EQajRQxGWGAN2a7SvSzmUrk9gj4843bv9HCzQ
SaTXMIWbvzyIXQaF9+14q13/5g/PW4fdd0AWoN3V29ASm6wOAD3V8VjOxG8ay2DafXJ89BVvj8t3
rY+NSNYv4FOnmE+F4KV0yLadB8O2DvyC6jcATYBwbSgLG8NQ37LcmrthlUPUL6PJL3vjMJARBbjp
1dP6RlBenjUpkKmlTv1d1ldvUfMXPIzP1CDC9ug97K7U7/iItffimhoyV9QUOHQhuHiKfHUMW4Vh
UFHslUffn2oCq27D03WGzx+hiCcJLLCEX28983RZ3defqnOdCqMnMkV49gE6iaU8qlD1skXhIjl+
A5uQGlNJgV8wfFaeLlwUeH7l6+02wXnk/bV22SHunnE9ujkVazSXjVXKoI+1uIPZP7IVrE4TLHlc
V1CsqGbw7DDoN0bSP0lCBDpHWsn3gHa9pipoXq6to7U/5wJ7gtjooAz/eBkgcDIrErue1yjBxCjN
z09kH8npLic/sGFM6RXnOkf+HeNidFkLmHNBATYm6I8B9mSejCv3arT5pKlDEQojvmaJzZX8t/5F
rleVPD/gCpELDYkpv6VHXXXT6KlN0uVV3qfaP+977SIhUI5c3VWPoLk6jOwKr5kLzj4+DC5f5MCb
SPEOw6eI3hxF0zmc08oo97BkjIGUZG59sxORPHw1Q2Ce2k4mIhPaZJHMXTgylKOSh2u9NfA+1+Ce
ZxaujTzWBjSd9gphaHWHTNkvBMtnSEdIiPzqISFyB2Ymdx5y18wBf/3PEOY0dCKJYPK6Xx77vCp2
Xtj7ulRn2HKEkbHbay9y7D2jRfSVO/ztjejMIcskonYBoH6TNC/7AeZUBmCQgeOqbGMNBY2FKyQo
loqgIUYJ9vsw+2joS8Gj6ERqtDG7hGlusBUWdgYzD8nQIIxrrAH/TG+esUwpPMN6lqTdVI03Jwk4
Ifeicr4yrwEOeFcS+/1TNr80rGPoH7Lmk/NaDeDerYJj/9ChSdWBl39NImFCV5ZdATA1BZcSJTN4
hAIh4cu+0BMIPsp4ZsDHR20g/V+vxPQ6bDtEq5qU5KbrjMblhRfqpIGCbPHmMmvVrkgguvl/dR32
U9uw/yrsOk09CTx6dvb3ACth60NjttDoyW5k3Ix10ayC5SehXqi6DC5zFnrQ84FSOWkPnWgeT8uD
P+n1rbfwYc/qga3mLNTPe4qR/JO283Ymd6r8q+KI1t6yejBrT80PTEXaNq/lOWz/GdqcIKlLdVRZ
iNGcK+nzS4j4c34x1um4EMis6iTHspKVv3EKLpw9+jg6SUpJ1/TVV7olLXQowxNx7kJDT5876vdj
/GhGBIn+9u+2q/SCvIRhxxxkHTY7iiPuwI/mCTigarovpxYpIBHu3Cm/s0Fe5B/SY7D6E82hwg3C
uQjtE0a9YvgVUyuNs60ITXDIf25qQwyRRc5nNfo4JgIiqa/cFd8xR0gg9+8pXQxJ1hUwAusgIHUl
CiqETh/NCKfcr8UXB0SfVZn1TzVLZ2YeAjwfCCKF4jPbk1eR5VL94bSVN3P5NbtQ/339ZaWjag+8
LnhqKupWVArcDsQNgWMQph08W5CbKwg4/We3VMF8O86B5I+myKw5deM9Kz7KrZkm0QbAHTojUW40
wHUgD1AZJ+HEoHj/tWvw9JZZxtGtsN6P4/X7qxS8rZvlCZDKN9nK4ARAWE4rXY0F+bw0ZOBUfD8J
OhqEL3LNK4wIK/MieCQ1JroAgT/sYF458Lu4/CccoduL+SWkXcVe8/YamvmgxhfTOZFBYPn9OLrQ
PhVYr4RuUmZ3aSq7NpSE9npjnt6+Ze5C8WB7krJi4bq1Zw8onbQPF2bfcJMSdlHk9cL4v86vUNj1
SR1zRWs86aKL24Y9+ay19jeLtwFZPHooVMD0ta4By6WCoSia8hLo2w2Uqpbn1vOCq6mbM6qTPDwh
U46wprV25O0vZJT2pDrR3NiyUR5jgJ7PqDlZX5LED4q8ztXV1zYysbATwpQvA/DH+QcjHXUtTMwy
XJqGtekzp9Gp/NxzlPJvbipJmZXtCmvjWWumIeTnt9lMWOIfC3km3OdEb1opFHXL8VuWnMBjXgth
vLX+pK/p2uvt80jrfdCi/zNOSCWxynL5RoxzPXBlg10jbIn72bm7LL+77+63ejhlEXL4ZtWDySoF
FfodUz8Dlr9U6FNueKgvopZzFefLgwWYOnUJW9zEdaTDI2qGzBrXi6e2/DGozPgHaT9RYlManCzp
Cwc+srHN3Qm8/F88K4ASQdiye/2MBzoGLgOAklNhnyDgpCWRa/DhN4MjDAp+vV+EI8XionNWfXYh
fFebApl54F1rJA7jqr7bQyOSPKTyQc9MKNwkEw6qLT7TyS4ma/FVuYA9k11ydJoJHrLivDZio5My
8lvFKwJ3wi9QEKnlYM96TZtMEqfJ3mT4S9UDVY8+DZJsoMpry7Ge44zQHdPw23d+sFh20nESSfya
x15GeZxaLYZMJaSl0+SIulZ/sdSKGzOMAOlAIMIftlk1lAdTVtgKnrCtCIOU0TYJVe2uyV49/X3Z
teWtrd1amsOddchHOBDWicMLTz7QdwofjZutGv3LiC2GgVKqbT5bKjCU60kOrgQ4gBCNPhW+w6U5
e3RZjTfmuB9tKC1B/+gLRZYRQ4ouWjoV1rsTENSamQa7HI4XOvE9uEqECeeLuk4ZnMB4IgTMgSnn
dE4WEo/Lk9Mi9g8JGFCPV7gC0QbtbHrf9fXQgpUfJwV7Htw/vzZSXoOi22EGzNGZ5mv7V/UCi8Nw
jg3TQgThkPJFnFrhorhLyZ1nt7ySoBZksBH7+gMRuv3jfwsghsmcCWkDOHD+PJGgX3In1pz8oSPw
Jk/Q5r23Wpta8MsiAMQCbGZlwOKp+KggvvOd4VR6T49Nlq6alf6YbUCbdel5Zkh2xFUIrjLgnUdn
GeL9NvoFTQjPtCWHETPxtOVNt3lS9teL0GrXVc19m+NLOgbyzZdmEhLxIOCTZx4JH5TcPFWZRQrA
ZyU5RPkolzz9/LEARpZS5JFKJ8Z4AASkuu8iGyAaqdn97S3RaMM8+1TO8JVa0yHyCd9WGV3VTNsr
RoBTKtkWrBn+9J/mVfw3+vIOL8fPSIPths37TNAhGQLiu8gNXd8Kt13tKCLgvPs+8I8czWBk/zFj
nVeQ5dBbZRLvm913eQX48Nj4Luuv4FMMGVVcmAopBUjLH7aU1U+r8V4sOVYF5gQT2xSussP6fFPF
nKB9+05Avam7MabD6iicvCER/7Vi3yotAyiddQ+MUapIKx8QDLTaQjmPO7bqPxOk/iox5u5KaOM2
gQVV86JqCCVmZzmfMkrucz5Cn6tHe+0oOfvrAfVZKHw1VastEvKJjEFLuBPYi2RBVPnl8s/M5mIp
Z3ejDoF5782bVwmvv/ZwSdZTpSX9e3+ZTVzKpjupAwP5iuVmIKv/vc4a+CogQ3bq0WZSxc9Xk6WH
OLP7Vi8TJLdZp2LFso+w86WTxv/a2pfgpYN3E3QY2gPEgouhfcrGqZknvwPblbq57inibHsF6eTR
T2C1+7VmchWXGCpzOBYpu2XA2/I7k7iFlnxcix5Tsba/8BIj6JcL9VB9867SXJITfwx+zt8twos/
trlxGr9Om0Q1oK0p2nEvfJn3lZhfAzx2KkJcoRUM1AE56Y1uMlD89kmNjiQGZJYBefIv75E1u2Ss
6HQrj8bjtve3hZeRIw+zwf7vo4nwHpU8E40amrQ+JWIFEqZ12Hw5G43O+imsR5y9hljYq43vxE4n
NAS3g48zedHkWffWQl6Nf+Fte5lb0JZXweLkLMnSR05Ulbs+NGyjw9YdNkpDPYJv0M1fiyvN120e
aBTn2gXYI0ohlwXUh6PVivDFYna9kZZM0FYIqgbXKx12fAs6TQEyJfpUF3HIW8xVvIz5Y75+oBnv
LjsnT9l8xrRyHjimves2AI3Rmpn7mPumqw5dJJ3UyBVzJ98FpRss+s65HPALMYCQbzybeE3Yinba
ZHIlH7n6S1MvEqSMLukOJDnUsE7KsJL5QSrg6lss124bj0wn4Y21y8My6nIuO/4HWYWXVf8RJxzZ
UQUxg8Ozafk65vsW8bzzGQWHAUp7B53yIkw5fLPnmZ1EDHkcpFTGW2r9uCVZq/GxJDA4u9RWEQmO
X6rv7oc6veAnkip7NbtQh2uHpqqzg7ZxDsirM5z0sEhd+Gum/bYpjdzL5qzSQi0Q5L+r21mqRTE0
DB4/qTmO62SfM/bH6CEjvfmUq6DqqJikkRZsQUUPib1UbTcA3hksVbXgGPRr/oFsf4FTHRXirShC
lhSG34fUWPhDyItOkhbtdgviLhEQ4M1kDs3YxewoYB4cQYE7wWQo7ml++lnsS/28XKj5HOjF3ris
urVptuwP6yRPiZCN8fQGyLsXujtUStEVCMN27nvsfr2IR2UNHDJ2Mjh/nk8dY76lXl9bPgNwnocS
3SCPByU+X/25Huk8TN71R54SYzq6oF4JNYdSvYmoG866mUvK6yqGJXvMN/bhB7aQ3fsUU/bP4a8l
1dtOaTcW8ADhcFZHZSYiFZm+49POom304kqxTPWhczA6wYIuqCHxB4rSOruV/pHToW42U4WOnVuB
V1mG/wQmckFrHiwtyNDLmsrBXWyirhEviPAJvYn0HHfOkKE6BsRjHnSG3hhpq3lCxSyT1BsMBd+H
VHKKLniH/A8X8Qvt6QkHgMX8Jeu8aFYb8glnp9JnbG8UhEZnAvMREN4Va0f2IbjkTWV5AzmRC42m
jPFyCwRs/+hw89OV7ukq7klG1f2Pc53wIfw0uBfeKLCJq88njdb6K0DMl8k/ZhzO7TwUNbiCqLFA
RzfbpU51yjYxcqePq5eRlQxfpVYPAbgj6+dxnJG1g2wv0oYaj21c8qts67jd+VHPALL+pYDledvm
Wp7hWK/6CGkq97p7LUke07atDZTnx2LTzwNZM6EsM6uPJILnAttXWVwn5oUGtyIuVWBZd205EsYn
HntB4dNTq60lsrNHFX2lzSeo/PKEs9JoNHnrBenVQkTqguP3WhJ+ok6yI9xqEirbKDcXkqHjhOa9
JeEOnGlbyog2l753VplOdzEoKeIJut4F/z38kEl1kU1i+2N/TaLNQNr/+WDlK43PZRmtlurQDsmx
BROIJiZSb7CjFCAtaCcYe45ToSQpLW8gfzZuXGHt4Z/jEj3eTbk+AABS14/aRrDYXryyiygv/28r
hygpyOC+odf9l/qglKPcp55nHgHWtNx3vGCcum5zenOUA/dp2tjjDeIw0nZGj1wok2bj98xPyiCq
bWDoqI2GjUnQhZjMYYWbQ7J9bWuAA+fsiiq9RXXSoVlKxHUoY5fuCStXNbxnhOTMLtHPhUfN/jel
0pLNNVrinC5N09mrmy6KOl65JdQpnz6vZsch3cNp7E8pSsxn2kWYiajj+MYa7lSPxGk4I71NFPM9
J5QXGV89btwzuCuU9VwfriWWKm43RlEtn1S/72jgk7GdTKVOmywhXqMQxRoMUTCll7fR903xUfEA
V1vEfLRCXu7vf8p2/W+ddY6WdgOQ4PtfsAOU5jxFupz5c9KwLoWEN3iP8phi3vfWmH5UV4I7KRbR
C+LG6n4DtzXpHdwZg+IZMl+BUuHWmj3B817FomoUrU0MpZs7yKmZWnT1zHjThPuYCaMyWJONx8YC
DoLDuGFQXnuKwabRznTD+ti03uDu3oqjRhw8e0UXxOkDhGLRyI6A8CCnGTrbP5uxwJf+j6uwy784
EQVPl2vRkmNizKi3LEnmmsCsQkIuWSHeICmMjSEDuYM90REnlg5M7YJYxabHXoGvtwYQ4Gg9BO7P
vJpxcoZsridfVzZCe4pFVC0J+c4j+9NwbZgHQiF98K+Qi5wN2MBFcs7TERJLWuiwho0pVFsEiVX6
2tlAzx7WWFR08wJvCC3m+r3Qrwlmeq8E++UVf3FIi1qYMDSuLkv+mprqlBrc7OpW486tsgcJyW/p
iK2pd7Lbgd0SiwXl+DsfciuCrcOfiyfc4lenRuze59nwEFTwQ5i1xzIgHy1fc5wO1KMRd+JDUf+I
Ms2ZOCCT6qd8m+/XpQFKxU/sYP/JgKv2zu+InfB7yJ7x2/QsIYyzZ5MUeah1bILDlspPXHjgn/ak
2ApAyua3oTw+bhg3dq+iSPU17x9GchCe5ityTgc3hieIvMmW/b246QSipM6ZzB23nUbueMhWkyVQ
99eLP/6Gn9LZy3oyqDuV8ch3ZJf5O4C5cAaavQflSA0jBbC7pW27acDQfJfhDXoK6kRHDzWOnHsO
7BYACHCfDnOKlENe/wp20y0a/x9yRtj8VfSgGfKmSJJgbVKHz7M2FiQbjhtp5tHRppT/p613+s3i
QqxKLjy/adI9S+KEH+lbZApepAROonlVFMOhsAAyXtkitqLmhxoPg5bdr8ENJ7B62EW7aVP2prVT
hmgnOIVV1ycm6PXpVFsdd0/upR6nd1ShohjkbeRFGtcgy7sGRSRpuU/vLsxSfB8dvTpZ30Jae4cL
0sG1Ki57jqisMWbIp+mUGTj5H2dS/8eNvSf0O9Ym01xIFSz1MyF3/U7MJftuSte+Y+uNEixhWXx8
e6STCdch2Xf0tTDbq6tACdAWxtRq+YFNHDDJC6exyPElbHzqtfJrOGVzvEt6wKJ/Uu4ZnkwhBWr6
zL0rNZoqSS/jdoDdd5BCKOJQifK58yuzjFA0Lk3sZKicEKYFSA9HCBzsUiNGmJBsw3fg0YgMrdcf
Fg0hWUnEa56kWhdSApyVHj8I65lBg8btv60V6PeIWoHEmNfczOf/Ckoqlx1YLqMZAIAfVFDjgGfa
Q31IDDmzh7e/vwL80ZDAn29JR87SfRkBVsmD2XNlARCXl3ABVWFGVFs5h+A3RgWMdAF0BTH0XHFB
aCD4vn95IjZHyAba7Gs99yOvQ0gTHW9MfmLwxiEG5iZztq5ker0DwiydpN1xai9UXn7AIgbGUe7q
i+h4MNv1Te0SUTyaRDLYjJbsBJ+iCFcBcwsS/qARJ1zMgbZtq/j/oUBN/CkepRTzXnxRXWoNDOrV
DKrLFi5UKXjiLDC24ibo54VTT7x9WkUhow2SaH1MNtipEnaeBV0Qdzb2RUm89HE9PBovkDx7lNTr
0vXEkM8CJsz3wTuTZmsXb2HWNcH41Thc2HTfhdQ9CM4ifm+zt3gle446FOBjYqpRusoI36EiLPZl
o+/vlKQDC/U3gviTkHNl2sRSXSnm6qeOllkqwRqtcxQMCrGj3aIG63AP4zIQLJt7Y5FMoLnrk1zg
zicHJCh9WojqK1VYj/f6EOVZNBib8isCKc6FitGT7Kk/JJwF2hQYQnQ4eEl1yeax8bm+HViokO84
3x+w2r9xS6VRr0TBz04Y4wGWA6zYR4tC2mMmCqoBo6wMy1a48DWUxLvuZ32T+rYQXnTX4VgVEuos
eAFg0auUZOzYMcIbRNdHGNNOZv9dhZNrRJJd4Eth0up7cGAXvTNYuscdQ5heo9eKboT2o07h+//j
wjDLwt1JtgLY70oDvbaKgy1WCqTS25+P+QiQH8dz5vDCoWgGavm9nd8/CbaWTzCSOQsGCu/jPJ/C
E1E2zvssfMkjLAT+avtK8JvMqqUKBnwHZ1dONsbnUyAkKAw89wzZEAQtfGvq0CxxFspnb71U9//e
dxrvbs05VcKR+nqm7D+PkjMSydQUoPR3FtkXcogQzA3jNAG+ItWaubNjGQqhCVylDhiT/8bZFro/
I/zsutzxGeIX3Sz7SMrof/XDRF7zRnHVTePEqmJbygDLhXkj2Do4vsSMsIyQpXD4zbPSH148vVw/
SVjO7YOPad5phsQeft65mq6s86N/6YhpK0DGXQCBx+YZOjJ3/ysvbWDDifQxFRG77XC+McVPlHOj
/xeZo7RBcCngron2rFbRPxhtieAQC9DFW4YqdlF9GP0v97iDGZx2u78XFflgzgfY4MIy2AqyfsX8
G6pitp59B7VZbMyYvS+LIHZb2o5hX8yjyp4bePOO86HKfmBKnKNDjw+D2QjxcaEztOGO75e+iBRn
a1XuTvO4zFbJMKzCNnhH+I0t0ruZzOIG5Em3pZEFB5pHPe7g1dK+PVNoUD++spYRpuf4N2sCFjuS
htrNGsqOjGC1gMjLOxGCkc0QFwwJlOyfF+KNIX7IPLWOFZ3V6qErYpMq2rXxrp47aHpcsBSJtjf+
Iuu+mPSfu9JphwJaAWx+rPQF5GSHAjCVJcg5LUxXs/T1awyeXwFDvpWYEfZTF7qFiztQxHOfVYIR
l+mi5caAvbya9i2sAdzQN9PK8woY7AJS51Zk81XnqxOeP/yAtv50DWKnJvkwnRLemG0SJ9AIcDyJ
Kvg2tX7EecW2AYMc6akOsrA+cladjl/pPopTHu0ii2zoiaZFkx2ae7/CG5U2EQ5+LVYRm2zEC4Qg
GdllpeHOJVEmB8rYInLYz9hK+zkfWAPEIMG0C84iLFMC2ON9hJmdjFRqL8MQdOjK7iVz93iHgWP+
s7W+Pr2glh13C1xCDv/cGPGOMq7cqF2x4bX7jXotnPTVEADogEzsxjyC0ZHKiswyV1/XRJaiR930
6zRWvhd9sao6OGcMuryCmsIfZ7BKKBDxbjjy2pywrEqfBPJVm+fFciZtGiqygRRW6tWquw43Gp1E
5KPgS66wz6AuYKjWFBt9sCUjqOlRijOtR3xBM9xQr77gIGmMWS8xooDKq2tVWJTPVgOxeg/8xy2T
yxDm9mzm7kX6MY/hQjBtHAXHYHMvF0+o5CGDwD5EPfmUZIxOJhiDxTFUCrWYc+qbNi1zG/a8ewzi
2GQfWbYzyoKcVl741zYxm37BQsl1McavlAevoJSvdZ0NjU1wP2tM5L+mUdsU0qSW3LTac2XHHBGA
Yi0v4ootSetPQ4eMhe2nuvhs1sU47PZbH/QRTpE7BkoemPW/E8M9vOyRGXNHk6O1uIN5UrWM/Mnb
bsrYrBhTFuuiODO8A3YBcPdJBvEYbgSpypbOhFn8bZ1X+A2L/LfuU0vvlcg0/4cb37+KM+Qz2vMi
YTSSD/e7+2DFT2nH9iFjc7Qnw0mOUeeUVFeyJpW2bLbRBC1nxC2jlHOJp8CVq/S7QV45SadHLYIE
GcnObf6naXbZodZFhhT2uVBKU4hB7F/GbReOACO07YrJhiAP9j1PW7ND/tprzsKzAAMCtp7HkEl3
FQHiZC8/dUM48wxHXgGF6vj1ktJFTpUsNVHs07MYC9M9pDQx2JpTuYudpBxaxA8DzJIvzETCPLQv
dzQ1jNCqtYHRF0LKlAn7wvID3apwwO2A0dA2JzyfmJAWxUHlpg9s82fGOn66WsB14Bfwc5aJDqAi
WdaqajSHX1McWMVy2hF3UlwAH+XTgQtEIL3PfjtO5ONL+DveFs2UWthwO8H+2d8XjBxDMYdOfoQp
HsnKZGA4aMt27cM+cpTPbMLZArPUBIekxILCslhgubCihIauCl1cJXBnmWR0DQrmqU/DR8IO/JIp
cWAkAtAQdhJYeHxRfLoI4w8dIQEG0uqzZhRo8PznMlS0cFme9gtSqF3cHxSJaFiddca5a61twhrC
lIFcS7u6miZz0ymeKRYANauNuZLS3lkU4ip9B4M3Dy1Iz7OEm8U5FjoOMRhtuTU8kNeV4V0ivmFa
OMrBPGRT8c+KGUTCLnNrEDZIdaUURflkurLcb7kfeLfLSfO8HyuqGcny4GOZhZI+lEOlSRZwWoga
fDsMci9x5woEabTcqYPGIyGk4lZUT7Jk7bflWxbY1K1cw4W43uAstagReQSV7UOfCAV8ByOCJgM8
QgjKhM1kxmElhqN73woGLVns1HsFo3DfmzJms+PSO/haIAYWRkV56dNGz2Zd+A4c5v/GYGP23Cpk
nRpWBa4FdNlVWDoPMMdr6u/JYx+8OhPor6tKWXOTLVvgWoE1XBiUUeMSQbEn8o29L82jTGI0xh5R
5SjJqpEfo9rJGuXEncxOYT+KlPe7cK+FkpymWZsICNi/i36z8CC//LUiU0yNSZ7xu08vbdL0Pax7
uLDnG7r2j1Kx5wbB7olpDHg88056FeOViyD0ZySwy5NRQadlArc3mdq0ICyvziKLEm2POAU9GavS
NRZkvXkV2WdeqEjJGYFTnhkjw3SIsCJw3lMW266aXbyIrSCUHjjaqmhcE43Jny7hwFemBd3/nXmM
epwd2i/BaYtQPUhTCgBRAk/KB1id4bs3ulksSWuxeeizWegQ6N7f7O0oLN8MCA3T8R6KDAie26+f
ZMUu8GAO6Es5R7/cGa0sdGKp3iZoBGPQj+nMR4ElqpxMxi15d2/XawGTl8nTSMNfnTn1l7PKXfUc
mEgM/SgvHYxmVT72tUUzvKuUPQYgZLzqpPbTvtNEekWTFoZCRK9nnL2Tba23impAEyCUOdZSc/Pa
AUAv0dq37GC13BQOO9wGHOXnGqDowtT3I4ABat9uf0B9AV2a4BONhgaENZknxhTuuEaYrGh1HVK+
0JOYHCitkm+i1ogl4cHeY2cPfyStl7JtLzPQjmKrLuSWI+4LmFazO7fhBZ3xGR4blLRpSX66B3K2
NW/2RYW2LXH6DVNSF0FKfmPv4pU40GZhXamMk87/oR4K4mQ095Hf7JjS6kEY5hwi4PIKk0rUfh96
/6mLQwS+m8Ah0TaMjncmNgiP52Oz98gHibwngfrrpqX66sO0dHiHSppdttTJtfSidrP7cwSLpzjb
v5Te6X1G5fMHNUTutd8M9YsKqpmb5j9krhE62yiC5s5mn43rzIJVjH4hATmO38GqW6cIsSzfdRAw
Vld9BU934AHNpT/9IRxv1h5uA1RYUWgDkC9RAY5tiACD/64ZupzKGadgKf+GJoqD/1k0rA8Dqg1i
xkbAPOl8+YR75cA7REUV6JqKa9feZvDIn0TRB6fw2R0UkAD2UDe8XGksRMwPYGAfsj9Mjjg0mvzt
L5WYN766mf4TL9w+fHiSv4qsbHWJ3AUiKtT+TWq6d6VQVVtz2TZ01q46S+jfqUW9z50sc3FSze/l
72dtZl9ediqzN3Kz51XJRvbOlzZl0LA8adNWTz+kJqMWQCNlTMCRMfPvPiyx067loyrFpQV6haYy
uEbW6bXffigH4sHcYzlODfiaNVbZpNnEHmVXE48xAEyot45WBumlvTawpegct3J7g8EPXZo5fJbP
PpHl4u+BERUwhMV+He1wcNtDp/uXqNVSVVwNE9q/mTgOfDtG5xzltAT/ZgxroXeX8UdVewIgNrwv
FVYpyM7j1SF7lEEhe3pphtjErLCf/kKlxURyPV4b8MxDVa2fnq798m/fWMLW7axD6f2U65WQCP8n
BlBp3tXEGBjjN7UbGtir2f4SmFDbV3OTXhJabTcrgoMyEF8luwhaUxQaAl5H0x3T7/pJozW5hhAD
wHHexO9UvEc66UYanS8miD6zzYDTo4OOJsxnK25kzNcP9B7WN27LT3yP52qoxNWBuT4Xz7vwXEI2
pXBRHBt4/y8d0RcPWe7oDwZSrqIugDL7GqFtFArmWj6nDzufkheN+tKeWuAb3XCCRSCmS1D7oR81
DBNH878rqaN+XY0cJth5WIjXb+3GjCyKG+3ewPva9COL9YvDZ9mRKY7Ewdmzg5G3PTXCBsLIClb+
brlA3MOQCS8s+k8o5TaLQ7IsdclJapB5u3z2FSFkbPb/B3LPgPZu15cHoRgLfDEmt7m+pLUUtcx1
Ud0hS4s2k6WEtEThhdtaUMxtovznJ9ZWiIf8FXRHQh1EC/OXHHI7Xw7C1eT6zB4Kr4BqEyyhcBVR
Uvv81x+nuOVD46dpTpZlLD1ZGgUkLNo9XmWcVhKF4GZVmFUF9YU9cUOEONWBLzrjq9LUNiw1fMhU
uopWTsuBc1+aYB4PZQNCTL8flzUK5u75awuemB+Y43h16kB2JWFy4r53GTDSglzu1ZjIQ7xyBD+C
U7j+F+jLCPNcg822DivoqpCO7a+f7CTnWNJPzQaxz7fwGKmYRHLRbvmKBE4Ln1HXnwye1GcT1PEO
X1ExMsb+PgYDJsjwK5z48LbvYNZ0uY/TZz+H7vVUKdNQVW2+QCUmNKwgflpkgZ4J883wZiGLCjEg
taBsM5Ea1S6u8APxmCMhcFVW+yOUpcRmHqBoDSMbqbp8qxIW82R9AkW0tST3BGKRuT7KdeD0mgQF
QoiqLb72BgEFQG+Jnp6HaRSELIIgGnmaBi8lchuPagcqXTRTe91QBkiXhCxLVJ68HXgcD4/w7eTI
ECIMtRfHp1irQ6Y7DVgTlrlSeIFvH5mazSQUZNUVPWUHRzk8u/4vDt2zcQnoMOdV3oLzpryFafrd
4FDTiHWWwXVf2ib47IpVaJLPfQBxldBAC1L/pRtzth5KHjXSaaboWkWMG2r/IoQAwjjmH2IwMIy2
XZK4IjId8hjXMh0muFx4UkBGdsfLnGm/grwps8c94Y+fS+Qm2lJwhfOaMICvGR99FFP8huSX4nYH
IfJuwOAfSEUTYkV46idjxw26bCfRIH3PDZkacm7F5VJbte9t0moLuBIulvp6TIbBzjWPgtf3V4kZ
sBylr6F58qXwnaQWKvbmUVpxvQnvWJ5DZ0M/M3U8lOeyw02QHYv8uV5CaOOgX6EyJ8zHhfqwpTWS
J5aX4vQcmm2lnp5oan7ORlpaAu5iMZFchGzKGQHmtITOgBJikacT7GI658N7GmX87vmwvA1iNPsQ
kGvjNPWM2UoQ4dgSh+0Z5IDqCfVmw3fbxk1Wd1lQw0lNBnmIhK4c54jIvc3dM5lU9LtyS1/3EQ9R
RKbWZE4FfKV4wL9gTfbsCl9p2tWST087gTgokgepNsJA44V4a3bbMdvY6RboK3dKhkWKkmsasA7t
V7xw7SQr7c2yHfo9o9NvcHN9OhpOiPZTyNLM3MXUzw4CS1ynbmeD56Z6wzDGv+y8cLOCrPQRriGf
1UgbvWwaMX3WP36+iz2JKvMOyPPmUW0EqMfeNiYqC9r1sUYas34aG6ldqvldqntntO6vg2U6SkGP
O1a12JZv3WflVylLsoOrS6R5BD5rWyB25MaZA4b8vDwEOcqXUOsgcPfkwfnZ5QROBzz70AhP/xnn
/wEQPeXPWdhwSgReDC0a95f387k7TZWUo1BkpaIgZoZGNRk6W5o3oirzLymLApBGZ5oaeT55TRGK
m2amZsPjPfuIavVRoHr2WfUqCZhgDK4iDWGAHNfmRh71gUJUZbXyB1JaLcdJ4j5WU6caMezQxaaP
29obv6AsY09/bs9RM4iyfhDkq09xQCT99eAZyVYSUrNUxc7/UYovue+6tE/oewK6lGrYcfTyYjxS
FnBRH59EBjD8h4mXVyKrrslnYkgF4C68S4eFlM23OBACWl2L5eXeIuOfaMQJ6Zzg3bQ4iXrngyxs
kcxVewkNPUeDPSvQNE6LoHPQqmohruhIH4+3WyhXtPejFjk5aVNxgwPMQAT7Ahn0FvStivm84V5A
v9j60VOjfl+DXQ6vMJ0PQVoSCLCHChA0E12w48V+CExc+LsKhtJ7yCniH8iHrL9Hl8VysfHk6W/C
5OizXiBOlf6DzM4uOypDp1FgJ0+tgwDKaUBnD7RxDRrOiCA8NkMlNl6hmhrfZ9nhOryQ+zevgX4V
PHIxDwrRiz1d8AgW/vG9jXcIDQHwOUin4a9QnehIyle5OS3JIkMSfRB0zV1c9jFRS7DpLYDZzIVD
wgVR9T4ZZ1OIPyAAQzuwKaWPZqdoOXDLSByLkN+Q0fG4j2CL3CZWfzwmJJ7Fog4lfy/df96fFtyS
RqVLA1Lw6d1rs+F8QLbeWaUjSsAT3tyxo8tcJWjunoRe7lLJxLpXNmsQIIySOITymdQ1q4FyyCCs
hjM9qrBZKk9QhnWtIKvDVDNLGnPxm/lK4ygvtwOkTh0mUF9htbcMs5wJ2eLOkfLQXPTj3VzJCIrD
dYCvPFv/TJi/ZoYP49KV1mxkejSxrj+AlGyfRMzPvkfbscRv7TE/wx8bxavw5CNe+1ll9jMRZqhO
WSBqHDHQZi+jSyKyrIxbCSD6JxkD4kthLOdpht5m3xnyI3+UXnEjTPicQgdjcN7IoKTgXmf+IXbl
UOteKxSElF+1szB4S8lP+F3Tn7iIPwp6yaBUM2alunGsCasj9jPELJ/sAQOC0diwnMDyfMUwa1WM
Zqe0XK+Coqu9/YOpE+IN7eHyUYDGXVE0YrRvTwZpYaWaV3VCHSx4VSLcqlFs/sX7WqKDgr7K0w/j
9uqNypMHVBZSTHlaft7Wk+IEX5Pn9PVW37YjQbuSdqcvhqq8SezWLUuk2piVOtj82r5vBl0UUIIc
YPH3+AqmyiLUmqgHF+ofW79RRansehTo/U96u2qXTu6G/E9D8SvX6mvpRB3LZzKLf1KRqeJ3jmFK
NuIE+3eJ2kK5TC55OLU0pUPn03ulZKlzVKRqHy5jBYjJ/hXzWZdhR1Nxk2YA1MsFv39bc/eHQhJ0
QjUZ+pcrF2fEYmQF/iWccRDkbRAmx2Ry/M2l2cy9K5feB5VWyFICHXBEsMt464vvvCs9GEUIkBHn
7lbRcnkr/Xc/Cyh+9qo/cXsVzi8wKKquBa96ISKDuHd0v/iSRLqozoUMDCxPN/uZFCeFqfV0PDmz
/F4kASd1fon69mDc0/nEsr9rNRO+1jVyvz0Afkt6fWFSPnmGEHV60e7/JPi2XwTRMOEIbsPf1oVh
sxyQzA49Ays6hmnngwkyVr52OYjpBL1VNLPARleMuArXj5iI10h5sj9IV6/rpa4vr28TAyFTahBP
zgKol/RhRcaQBdrr0Si2TlB1nDUfyACGNtak4d2w6m5M9E3cqyEpmt80WTvmaonXbm3LZ2BJvN8t
5tmcIT2XJBa/pQxPplFyW8njOBkl8sBZzMFGYxkylEpaFM8R3/uhdOAKFvyLHH+F8ILxMWYOAzHQ
Hk1v3Bf/GAU6l8rVZG8oyZxrnWJobGib4LUoEUTeY7ChoDuOXYralp+IdYdvXnkhawFd7PdQFLez
NUJcJYCDZD9hrQgC0Khip1uHfAKc0JJU0kX7aDdJpLiXPwt9pUKZdst7QsnA2p/S344JAFxoT+p9
k0GIwxZqNL7yMlY6jJbCkTMQ0F5Lk3zE/VoKwVD7Se7yHzDuVEe7rW3kNLmAe5YPoKrgxNoqdrM5
lhUrRfszY/L0XIoWmwLnFhZVVS6MOQDKWQw3CfZyKkcwrH369fLzrXb22SP+VKa9vL1oXIC40JRM
U7mjeMquxm/tZ/cyFFXTOhAYxnTGEl+1O0D0dDSrqK7sJ2wFo3ZyXZrPOz3EZ2bLFtnjNVbiYKvu
mxbjBoJIjSbIf1YoZnP6kC9RzDSbJsMOq78ZyOBgFzHlbutzFfUp9UjndCQJaEGO/YWPTanPtTNm
7/0c+K//T1kvs8qsLxxYsDNb6lF7rSRrHj/CFvrKy1ZfvWnpi1RuhWrNJU2qahQVojvdevT4vxIT
OQRCKSrJklhBFH53mDIhdWC4R7A8QsUyUkd7JWw3w5JDMZtsaGOmDpHbmD3d6mYvS3eJmU0wSf5g
nJElTs9nS/aLpqEKGicB62v8g0uN4oANtTPm83a+lafR33FuvgZh72V1yMSpyhlXQWJGd3dKDtND
RJWEwvBZBTdBgdbX5dBjuqlnoYqOkxcYcciGembC5Lzfhx8h8u90+ZxEe+LESNKjAc/3lrQNvM77
jmFqYzxGhjZoFmbJN+GBgOvwZr9wegZd2W3ibaI0HXQwGqchBzpx8qulwg/irXtvgFCP/nMNu3+H
u40hps7G3n2o1oV6ejWejWpBIlasYCOqLFPMh4OfVnLnoPeHjnaKTC+hzJzChjnVMyw2iQqaUjBT
hJJ7yZ368Zz80aal3yjVhftVm7gtbUJoKu8sU5tf3BBpo4kOmqQ3HM/1ggXGw0ICakQyuF5E8gMK
hN7+Gq2SCmTJq9itR4psBw2Bo04veZCIM6300qEpNKyr5Jo6LAlI9VcWN/9InLBnvhXBYQpC6wdF
yZc/6SAzLVZ9cJrQe/wP4JvSIixHYnz1oerS9CTwbNiAs264kMVNb6hmr0UUVpThdRW5zaCanVny
W8yvgqZwU3R5HPs1wzsgSbMWi52Qnb3f4YHmccWV4SDkWRY7dnPN+A/YZZv5QJvxC6DDxQfwa6E0
eqoWOszaHPOsGItAIwgNyWpIwZ4C6MfHb6Y+PswnIL/kpNSjw6V86lb44LHoc3QwzyDCqOLCMR9p
WjvzbUCHx3BT/j/o9geDE4KTGV1YFEYUh6h6He9+phylNf3jGJvPt1YOlq2XvlGut5KVgvXL9jcR
ZDT8175Su6IAK5bMHtm79pMfM85cEhIbKL8I/f7VT8NPx86F8JprmJu7LcPlp09mdbTpr9x50Xdr
20MLS9yLiEIhUdl5ygL6PAp/GzAlgPd/ZvJFs6BrGlTYpPcFoh+fe11TCKNZL8x9x/kFEXzLHH3G
Cx0PcoR2mHtALnhOvexWnJ4/HE5bESXYI0DBQEGuhWqjQx3XQYEhKDK6RDhrWvgeTVITnnla5ruB
DPNlYYXD/psZEqYHsuB6c1Mpc1a14eN9cAygp8udbDxuGk2+c+GVM7Hs/5t9Z+kZckcpX0i+cEoz
yscYHZlpYmZJLRd5cwtYCHV9XHAkIfYmmSiF7YDPzofBAr1naQ9MDMCmTI2hvGBoER39KzurJ5NQ
Vui78V3E8p7TfR3e8oSZCWo2TsewfNYlVmTnpJLmFZ1AnjbGmtsSnAylEvQOY68zsR/WsEiYNHWR
T9xdr6cWzzc5eEitiAQ2GOT1VFyEXAFTiydLwe5sg+QAvpFkU2TnrgD+GxMIUELoHBp7OaUW2omT
+I6PS+N8tA1xZsgMBye274RXUE8ldie/5Acrz2ygolOB/wQYQIzFkBRIwepwvLf4qfBmL6NKfk/d
0t/+y/aU4BINQ7yPK6bIl3k5OUQkDvCNFJSU4RD26avrk+pKw9IKZAod+elg0h47oCZB3PH7qkvd
+UQebIk6BPjI0j670YhiNo4QSuLZp/5ZcXNLJs31vKidyyziry1Pppbryjs97Q91L1MCHyxmQFKc
d9KoOODhP58gV9gSJx+GqOiOUMfBJNUXBhQSZn093dMlmVkhKSg3HrMlpRcQ1baVHYITCW8u948k
cPuh5Y0/UaEqqCGv2J1s7dsFGR4G3Ipwa1Net6kTV4LGgypZKN2tFLGZo/S/NB5Bi/8N3ZHhxqI6
5QWrnjj4OFQyjKYPJPgZR9KCZF3sCiWQJ1QzIGHa8tKA1XLPh6a1ufEBQxsO2txdk2EmQ5lk82qO
bTwDs1xcM5NVkKUoRoYc3S1X7ks9Pcc6DxSEkG3m/rmsdJmiZE//LQFCBRYJxdRVjDYnmwpPyJOO
xrYTYvyYRwgfXiujke1GQz+STSwnZ8dr3ZUoV0rNGDGIlfEHqYuCS2z+w2iHsy8HB04TJOmGnoIV
NYbUo0h7d3ofYJR9YlzvfNnnjeq/oaBqVpUNGogrymyB+wIvURJzhGt9D3EvJn59TeKPjqxEvLGH
ZP1QybIpECfnToNJtxEut0wehsOL6Uz7gip8rRXCYDsrQFZwlwW6MT4FWK4oKU5FaLIk+9da6jPA
OTLfnFjIjeCCL6FWzEDzY1FOdPsF4uTchczsQ6KQ6zOzpGS9a9WnRi+gp1FGtLLVg5W75X5YSpaQ
ck/Q+okNF6Jbl0UARTJeDwlGwaC9H8U0hjfiYsNK08Hyaz8+gOUV7vXYYc4a8bSgiVhzhRYem5EK
RViOvanu3sMvr8EOsZWBqeio4wlBIurru1rfKC4ge5L7DIv2yi1ldOspaMYVob+K0WbK7va++2dJ
6uVeHvZkcl1xK0GmajaQz7NmHIgPNt5QLMEhekcMBx7EGp6klniy0SQOMbl/SradhxVOm9x7knWO
co4B7g3K38/u9TsDepLDrhdKhcayudO5hrkNfHDdRL5C9o6nUMI6kDqO1WGOCFiJuzn6jQfPRE3h
gdHeWcHKbcDMyGFR/fnudLZkX/8gfEfqgoihoXln0PtK4bQCl6yqXJNpGBgD9sAW2Ehh2qfOq01X
LlO+H4Bfeies5St0E9yruPZR9tUZ668RAKCHVPzhnueeQfuy6UDZNQRuRPTVKvaM4MD0T144wACM
O0r0Wk0kLrso4CgJ+o5Vzw77sPvRkftXccYoMzVb9NdSRY3AzB9YBpKmkwGZWOzbILRkM5o+A3w+
zuSKUFouwq4jwWgSN9O6sI4AoOkIqNOCNgECsrpsXEIyIH7adTeLCLDynM1rOTya3Qe3kuaRKsZR
ObXPT8sU6FYA0sKoL5Kc8vfBcZW58OTcQ/WOAkxcvrVavobpCm+OAY0SfCdo3s1WjX72RIKvzcKH
6G/gLqgDy7DQvy1uNnUKIngKg1u3xuNmZdhoNl7Uu8l36SQ5rkrWjOt63cwVFRmvwsTDk/Aav4+f
nayuSwya6xh0GDWXZkSzh+pyn21vj7YMK8ooyaLGXjX+pY0tL5r3x+RqrT3zWtc3McG8W+ldg+xu
Koh2zIYln4J68i+eyt+ZfrngDZTd8KnV3D3hWo+RlfKtr9ewmOFQ0ShUWIjlRaym8N4q6fytW3tg
B0NszPEZS7M/t3Km/zFc56AhVuouCBE27EqV3T5CD+EjYEwxNusWHKGZ1suKP2VmqOS3SsVolYIG
VtgHtyKGBh/EDgxG5VMWPddgN56QjMSSYWX1Urg4Rrgjf0CQkHyh6hNZOW5DaITevnz0O664Yh0d
c+KiZNq3lMGpkijhgU2wEQJywWo55bPz+EUH6Ki4l2A/DaJlsz1LBgjItff2TFJSnZGVYxDEhSFm
McDNJWGrTsGxZ6pSRyEMes4x3RDDj3qHr3hmq8f0NHXYBCqCI7Ht/YisBqNx9WR7YCRV448egq5E
tE6CNehAx+L1RK8GDQ+T681Dfg5L8JH0GLk/oWx0KlRbm/6ykYVEA/ePZ1rxotY8iEN9v7afwJ9D
bVDslNSMiMzT0lfm/J2Ju87owfvu4rDw07Z9UBPYoVDNp9vAeZtPWAo3V5RrATPTwIfoBw+TGbre
ordy6YAuxnPtG0mIAnDnv6mbyTOgsIgqv2YyUmauo4V4wehqHqWT2vk1tOUnTbhkD0PXQVssgj3P
MiBv07wBbJs3FG2bJWNAtA/Sv2ur497T2vhOcnlnX/xL65ORNG/P7vAyhJuWKhKiJbYWoRTPAvOi
jdJ+PQE3kSHNgxYOLQVNYmYvx82v7gczo4u86U9HsGmjzlUsPxdFhjDVPF96w878ZrxOkzEI07yx
wIMfRQcBKoVdIntaPltRzMptclX8RtTv9Xz2sXUy8/C6jXFflLSzuVFOnUsKBVuWDWqjwPsIgd73
bKBQdydzm8T2UnJZWsygkSVavWHDNWDHf7gO9YmU4R3zVZHvJ5+yCHApqf10zLxQE4vkXt99AaQA
PozbTaLPoId2g75SqybdJiGpmAeE+r8I5Ku5On9qMOtlFEF9ERqJK2bXN3svZTcosmVn39hPxOO0
T3o3IcaZOGJl5YZfGCPw7fuPi8Uwhmphqkn9UR5lNcpIobD7TgWFlnTA/XaacxO0XUR6hNVnvcp6
a5hIFFU1YxKMr2B4fiI6oOh4imXjG/6v8RnhKTlboxAiCOVtf2Eo4nqY3Ji48DuqY5aJd1kwlF3A
qdIbnHKmj4cRs5l1DlWHv3IHeuJqGk3z8vTyhZd3ox7C0SJORekOB6U1aCiaCh7urw6nGi2UZrt3
jnU/PYGoUu7H/AAhcJYV80+zwyJt+noE/oArdwfu33ecb+IVwJSAd6Y3ZMuhESZLJrpRmTvv4USA
wT6PmOfl0Fh3kqZn+NikNNpfGoKIO/1fS4ORjdgdfoBhRpot8dpz6NLZJ+goNX6Isqwb/byip6ye
T37afc8rXs8PdXv+xAIoO39dOecbrcUwLjpoWJZ1KBxXtpC7I4K9+S7Dr1KkQsDFmx1Mi+wqMkHI
6QEyz0l9C1zs1n6mLfex2I8m2snnyr9l+WVckHMybYSK8FrnruGQZmPjNRQKtGQvXG2ytjNG0R4T
SK4PHzW0hm3+QTuGs4dPXwPtFab5Hz4DxlAXC3dFw5dRROGSZcgC88hdMdnGUAZvpIApY/CsRQis
bUv7thE0p0lQH+zz4eLR11kenLvla1HG82a08+WoombGfgiRMzHgjz8PE7B39MY1qgxuq0a/yeTd
TW6Qikjn5CL2PYiJn8QbSKrkVHX9LfP6odrPx9tcpOh+VUj7IqKKN3G2fW4va7ro+jyogXu0onx6
BNjfxjHl25ePlvkgRD+wlfBxSCiJFOJXEDHCXtipX4xYFbyByaClW1UfyQL2sTOw9J2zA/Qi/VU4
qgSJ4RuJo4rRT7E4fCi3TgAQFc/Gsksh3Sd00lC6mc8d37hxDzFJTtAQbqiDSk7egGlCBsiV9KV3
0hhlRYILpaOnGKIcLY8SerR4JRJdXxUkF3qIH2FGlUCexi8FWCKY3MSjdChtGG+JM7hjaiWtVLk6
hqqqmn+3cz3zVyRveK9g+cSDVKxxMuyryUwYbqAnfxrdbXAZ+s/MJDYXTphVln6sMrNSEoShcEgP
OpZgYUe/y7KsAygpFJ5riAEnjq1UEuNfeNeRtflzLluThxkclgaEHTTtoAudRYE3WrZAhjkcs5AT
ZaAskZMk+iNXU0mNsW68zdno7yyQqsJVFC5ZhF4ab7/4wFKQd7z9q+RKJLreov0COJkW3yNq/GwN
XhRFKfhXcZqLZKb4yIPjJySS2GkKeIu07hnzD/omp94JBLpilyoyJyFhwQ+h/y3+A5IlkClT8Dyz
+NW4k4VYsEdBtcQVGatXu4YfIH//nkpE43ZsR6ZKQaLKPl/q+8O+1OAGzybQINuNteNhj8X47lMP
G7lyEpBXDUvf5/68loczWRlxCdvs23VFejlylybU9L8Yy1QfebtgQ8s2VXQfSrHCKbNuidIGDdO6
MqnmuDCgWsLDNXLMcfNV+mWr6nrWcfCVmfBVysnbdHsvGq00SaK1nmrw9gUgr8sRXHYOCNn91yz8
18SyKP8AxIpbEhfwm0mR56QywOwvAzNvgDfoyTfiOqkkLljqrpZrc8kKns9TDrrxsmFZPdoi8kj+
GwdTc9EoUZVbaeEYdog10WnL3VH4KLgzxyQ077toYuTpiLMDZDSH3DKfIXM197Hp08aEg1mv9Xo0
HrcItCljObFtYWVaDHV0dwPVM1H6BRFxTif2rwdPdFl9jm02q5HMLUNDYOR4s3dK9MNUpyfx5vZE
0nfixZI7QTWlAewfINj6GfGCK2WBljt0kLvhXLsXBaB501wVRM3YZh43/NV37e02G+VqHefzC8bZ
NpsRDaxXHL7x2Cu2YM9RJSg9mNlI23i433wGn8lIngfJtJu0qX2gUa94+WSlKdIa+EzwEFcaImqb
Bvw38oDfDv8JPCM0B/8JRlUT0HTpdSn1WwmfgbCHrREZ5FbLJDIpy3O5KfegDSeeUcE+Sd4Gho9H
Gf9PosXA2tsA6yfweBNHZNLwF2OPheq4b5k2AXcg+H7BWDXZoMRAq/1vnekYrXPJ3up3dKfapoiR
kN53B8j3K+caX2A05wuF5PGLga7Au+nXpYmSorFAp1WjkWBAdwIm5u3mVIORnKZkvaGZiqVRk8/s
XwJ1bHhWI7fYRbceA2hRkOhwOCvZ1A5acT7e9cldkZBpw9zsq36OFW8l3HsEnrhWfEClB23npMgX
Pl7mrDuxTqAssP0AddYP/iKgEH7emzmpGv3X2ehnGa8mgq+sfWh0ICLg5zD71r8hCWrQN780vQxH
tkmuahGaRn/y615rD5dmq8+rK/k6yh0e2hcbM/XLkwBPUGfQQujvQuwou646vQdNV/DqdVF4LW5G
8Fi4Xar3DmdmMv+S5Q/n5OmwPJetFO2TdrVXISGGfE4EDsw6xjVqBDBPQ577NJ9LpvsUzJgegLHj
qsSm5cSOCdD5pBidfGAhRu/rlwWRvnupf2zN9uV55PUDs6ufsZoUqqiL0EaQXOi9am9UDPytGvWa
lNk0PJV5eJWzx7e/CDDyqCOWX9+uCyE+t0d5U2ADSCDoVQ/H/jFlqvk1aUq3532yIDBry1xDCcmz
slBMBbeNdHne8gSe8y348f+OvhO20LhCK/gxxcHnXsn4Cp8lUnCgfF3VDRxMv3xYlTzSqwkpybI5
5LxVHHs7bxox/kLqSRkrx2yMnuFANej3uirbD30Oc/gNhkdAxVObUbhrdfELpGDF3NQ9phvg3r4D
+lGSevPv2FlpKh/yYp4nXIThhF6YV7+qrsPZwqG4kEToBioF3mMpqgQ94iSfLi1C4akeLx9crb7/
PQ/MKpx1BCglrjNAeIAwkq2/4vMLkq19Kbzoj5VLfAbx8MRsKh+Hu/tUPvWr7Wk9xammbJc2x4fV
eoD/4pS9g21NZeeZhdCwDn/BQ+H5HWHw34zbcLPmqIGYnZmTRgMj0mUsvzX2yLK1yucVyx4jl0v5
9Tvy8N8xNWo1nnz6gWJb577ECtXJJxOllHh0SPvVWwX+2sQ+2GgfexSjsnkhoap55VO56yM+wGk5
CywPFBilKAmzXU4qTWkXy8fGjHq+qBLbzXn8OZ5lpgd/3VZ8uYDx4RPCxHr+C0jxD37O8wHNllpV
6e8hjFjW1457utdN2A+ryzMS8J93Njo0m7Af4wkFDYNS2z9vQm2OGyZoT7y0ryzRoe5wQrPcNSMm
9Xw0YNxSJNJ+VUiLzI2eBsbmY552HUiCqWJ1Gq3Z8JQQw4Di/3ChYEkzgpZbaDbQKw7a7dsIYTkq
CvvvsDogQA3xPjdEhM7l+2/k/Ff5UfIZrxB3EQMtM6CdFNwO+m60jSdhLaSIkf8mT2byTcYAf/yl
JTxZJbosgU5btMPzW34elBsJ940zjt6ayBYacE9+SXqEuFVbVAaAfr5OQESzCZTZWiTl6DIUUQKH
+siZbudZSZxipDqt2hxkhS9D4W/MTqlGE4m/ax7O6a3qAkg4CWhKsAK5FsVTdEqufVZvHFAOd69n
b7SMhRxGiLzQhaDEqcRcyQ3WwrgijTgYss1H8Njy2rLW3IIGgtFFOg5EojDrkE76DM/9GxaUrC/Y
fCUkLuXK9KkR2m+8osYfBjcZ4oLnZChMkOT5SpJwMtKWAHc1WimfW48dkgMVo8+JZahVpDlU3D4A
130bL9VyqzbCW3lwXP7eg3VlhuBBxqW73KewKmUI0Wp+pzyPqnnhx4PLcaW0Atle7RnEQqnEf7fa
Z+mk/dgK3D6wrFGVRpABiNr2MtmauzYCIDFh7A/kCEMP3AZho7agLKDBVDf1YsUokOhWM4nj1Ek2
73d+T64fW2Xr/33F1fTGTDC4rsW6B3SwfAERoH+gM03hlDFdnrFvFSbMrbLq7hfakV2MnGQ93+lA
gDkdN446XrgNMwCZ81xof50kl/FXPeUNPM11Hz8Bsp5VCnvHW/7Y6cRRpbZHiVI+GVAF2qVJQhgu
Bcker8kQdNXmF/QdU8acWnoUYDqaz/tYArYu0e3y6XTme5sv64jmD5XF3j+Q4Qw5V6l1YuYAj65z
443PeujI0Ig1co9RnREat5WbpgOkl4DpApuBRa2VidkKBYKLt0AbEom9VSvefwUkt5rTHvJtKItI
ycDYZ9aW+uL3ztAMtqLNjKqRiqU45gfdK6ElMaLEgAgb00rHXTKhYVKILDSN815UVHNsRZPKozdS
quJuV/w+VOMQyeLbSH6AVPakD8grU2/IoLYC+0nqj7wtO+EGoSW80v/Pu41aQyXArQAlz8MtQ3qq
RaIqnD97TDKloj4vAz7dsWZ9BqL1QHUy1bkEbbCRJoVXCafTmXXsrr974YE3VkDRiyYv+bcF/gW+
Lh52l8PZUYTQ+4yY3irLkAxTVQEMTYpR9sf1bpn9fC/Js5WI/XKlPEixBFWrvGO5O6sLD/zsasJZ
x3erDqaj2ABti6Hg0sCveVI0Njrdk1P9tgw4D+dQv+40GEaU+B7hHhUkQTyDW/jY4E5xLa189NNN
ex3CI016OlzGb0tBWn8V2x3Q9M4jeIPBPD4JNMS6L3TXURrTeubaT/QWE4QoxtTp189J4BpsxUAq
yxwpbdgsohnrlwn+mt2+cCLX2N5gYw6qFzBrlgic8E1qHIYDMUdtohAvDlFgOt29ZpzvJZxg4Pz6
jKSYuziOetgTPSetYWP/CU9s2aBbFAI1/lxIXp5WXAr3OnZWi5q/iTLfQbZY8Qe3/aCaOvdkyvzc
EbnHS1GYP/TAJfl70+fZtVqQjV1KRbScQVEWveCGednjMAj1GHViW4Dq99GY8GNVdN5yBqcOK+hR
xaIqTkCXQ4+dpqap97Mhkgt8n7S7PRla/Oo0FgkfMQkiqSeWpnQhZGSUtZj4ZQdWO3Nzvhw8TluE
lHOP5Ho3f8wfiR5L8yjufw0iRrGlqgsgMu1kfFamDEnj5XDuvmX7B46aNfIL7ShreusUxKRZ70M2
g3jI1PQi9cH/cDaHvs0jK0LJzQ09hwxKJ4lrQGOPOjYPPt2702Zib/V7qb7axHBoIGv24D7lNhJZ
8yzICOQefW7XlF3rjL9IVaxvlxpfF+o/MZiO1Lwte/uoBwoHz1hpNjTaP0SpfcQYguRMiSBAI9kW
eb1nnDYTzj0w3DI8hkb1EYkbRk5vn2GXShm8BYGfcITr2I4wy71M0YxMsm3vzg8kWA/P1w8qFfCI
KHy4hsYiOgZm7Oier5uGObAw2XGzsI09RhXldttM06hrAbA1quifGjsC3JGh9YVc5fFjAen+RWFO
tNLnnqM7m8xzLjdiR5mqP8Q+j6Ml4kE+8bRYRnlnz8q2wqOQvV6V/IQvg82Hod6Y9pnz2VQQ+G/4
YS+JomycxsLjdWPveNGyumQoo7OWe4ocnsN/L7X24gUocHPA/mL+ks6JKuxHO0Qp9/7QT3YjOkM6
qQoM2EBdUUXeYLgwvsqyDjMQlq4ZKtVWsIqvqYYkoxZQZk2PrWKzOXTuLKbFDETtr9c1Dp6aP449
XCib/aAWJFDNKdXTnGPfzc2CbjUOfkQE7Ew7pikhEidf7OQk/3oU6iUuR/LYYxYlMWSrfbqr6ECN
hO2WMNFj0X2czp/7VrC7ntlGnDaDujq9UxWEv4nUEfhrKcxID3UO6ls+apcULtCjhAnXBazStlpC
Od+eHeMJZ2BwTKw2+jeLjacSgOFdW6iRg364INVzzWuDTV55GILaqh9fNPriFTf9Tms+0wV53Z4H
4ptNwor/n+hkaFndlSowSykuO42W0Nd2eAB7MliuzB1dAsIU4vZfLnTA/h9VwDWllKUdpyfKBARQ
eFkGxf++OxAx9VzqnIjPnCknfIh99oPo9tz2y4j/o5nS8DhQwGZ1DFs0NUyp8Kmd7a1K2tLBwZtX
ODjSb0QSb9Q+1ByLZdKP17ool5owlat+eSvx5m8yU2JVwmbmF7YCXSfeWWyGlAk0yQyQDawrhpcw
8IG3tpkfXflVJ6K/bTOboNbeRJOwPdAA78xP+F5UVF/uZ2zVYMRU4stx5EmNK7L6uliUmsR9J8SC
CDGDnDJmE3K3i8j+2LtBi7y+Wl71IpvrrArxUhYcRAzHlaDqSrspqlVlfSWTUpbDJp1I2v0fWvOM
Zg7edfrmlAT4Ag0G6o9WcNS+fFAXU1uuNQv4VDVJ2MZrWNn2vD60DQs+SorjVRQx7md11Vv+Wepj
StOmzYB4KmwmRy3nGbd3ZNbH2yunjKrumdUkwVUrfQ+kSfZSSZapXZCjJrXiVPBXmMFIvMrqn7NA
r3HVnKWPbeEOglzSt9y4TfP294W/C2PHGH92eQUtJ1t1rd8ThgYXXQdd6Eh2wQmSIp1A6ir4XOH9
+kuw0OlD/eASfhTBszAqh1fWVI7GtyuTxC/RcURSiUeuIOBVb78pd9N3xhcSYmK+3etw6Vm4obIs
CNtrkWMFXkYYid5DlkYsb8SNOGJVJ555Kp9I/+QPwA7KG6i/MjpIUUELd92mWX4tBuC6M/u5xgup
oLiWx8DO3A+dxUUsOej1qo6uVHf/4o4w1XuuSW2NrAhS/XzWVJg17mT7vVcMs61f6pjs5tcFD33m
RdUnpurWQLGPGGWBoZ+ZMM6D4zNZMuhRoHpbyKL2a88mez+TW1BWxXu548Kac0HcEwFjT7vgcz1I
QYisb2yQNIbmsp9GQzgQKGhF5WGUurAcBAdjAOZ5MeT0ASMNfPsTBLR0OygdBDKh3aJorqVhvCfp
8y3N2Kpg/K4uImL+vJXq2BXMaPd623QSwPXBkCJqD/5vGyKi2Pat7lSViO7/UFV7VwuYLlDVccqA
7V7ZNhEB5n7AnPzVYhXcDWOtC6j5BCH19mmouTSz+TXnmxyHz9+H9JQov5OraEFnt1wiZFPjBVJ5
kn3vU11/kbMTCkviuUp3I/BeCUHtP95iVYCR/Dr0NpVvAumII2kEx8XIXhUfuPWvF27sRvTvK4rN
SXZcju6SqJ51dQGWFhWgL2Ao6wq+T4bTLY2WPB4u3uF+i0eMNddb9yz8MSFKmvG6tkb7B7uFQQR6
93fg4ALGR6Vp+p/2YHIBHy9jBIa3zWPwCo0euvp3tjxIUXTiboRqZGejN0r8VtlgDRYKNNsOdLn3
r1g6+j0jJfbAAoWNPedpwfKiw82b/FPAyqcTnzPYxOfC4AD09pdH9rK0/hkdX1GQA4HHWbvp/gQH
VAx2iRZJdTBjhKF8Hlf8j/wV6AjbiqpzncIIqZ0iqRQjhBIKp5XsTJubFTb7IkngDpNiQxbxBN2L
hxyv2cUfuXW/AeQbWw0tPlWin4/l4YzdTRK1jHufsF6L/HgPz1BY9hJNow9cjMBypKwrlfNmssG7
XLPYupYvSlgguVF0VdbnxWkk8Hnn5De2idRkFLo9HJYqaRDIZTbi5gtsmLbw8a4rQSQVlDt6jRbw
zl6Za/52JqWX3P239IWslIAAl6qS5OhfErBRLU41/fuAJHxixQ2XUknDnzCrNJkZVCWEDozshMZa
JG7UrDLQaKRflPRRy1giGzP89SpHkXkHDhfBwwISFNKUalDqKc7O4J2RdotkT57UHj2C9W+OYhjO
Fugx1/pX6pBGsVffbWRTDyQKmKUQ0aHq0N16/phMIkqrjdNinMYitahJMaiGGMVHp1aqDlGtOV5P
6WWJZ2cnFQoCmcRq6m/c7twept1qkaFRN/ZoxjQC04kvld96hTu3JInKkujwRL8A36NBTXL5ypWi
IP94P8goaW4rNI0llvvf7Kwfu/v4QrCym62A61VsgtqFksRR1d12MfyAl6kyPBv9uLd6mU4XUpE1
ISJw0o/bAEcQrHeeOUuEEIoVDlRtoqIxKliilDkNwhRejc+VcWqWLY+WC52v93iZf7iHyqkPLq7+
xBRL5HsZ6+N1BDDrTCICRWt0eTK9+xWEilAXkffZWg7kTaDD0oHEGRfeG8XgF1O3dt3bjwEzw91Q
ATmZBg5pcvhyYdm/SzyMpkxTiJOdPDxOHjADTXN3/Z49ku0GcLlq9faqd+hP6ujMuJvKLOj5D0ie
y0Ew05tBPJyFc3CpyCYN8WLVOk4pDv5EZXoRYHh07U1ytiZu7Oz7Ct/ywo5S/10TliTMLQ0zpQ0A
0/7V7HU0QNTHU+yGeoWXTyxZg19WQIM2x8lGnTF8kvX5Fz7ipL4e5kzbgV3hz1B+Pq+99vR+kq25
Rrh7i+OFXN3k9C3B1HFDvcnTnM4AQVD3XbJzOnnKDCdX8MDzsPCP8RezvUtquBZwgKUVTgYfh0Fj
k851Vds1tbhql29xj2sgE849ajTPgJdy5HYQd87HSLPZa9ELPXMUOaOy432/rDQCX0MCZMJuvo38
Ay8hqAj+1Axh6M5dV/uD9zZjZ9O3rsnvTp5PEAsBN3Vbhxy9spe7LHS65HL1zDCLkVIOpt2qDElu
ReLhg+oVtJYSuuQaPuJZk3VEHc9UmwCmdf64/KcmvARDoGoSoFv7+ZtD2011t8DnKugrghLEJGGe
Ip3b7gAlb75m4TiSJ6q8G1Rm2uRV/HrmXGRLH4j5UktUZlJIf3DqnZ4b3aphI5yYnluaHfBGLnEq
ekwm8ky6vuDB4KJG+BDJz+8aTMVJPBODYyXAijU5Ptw/C2dE05LWbNs/U3hIDjACb/OiAMdKaH6t
LK8NAX6Ob+lx2VMkqV0dl8FMMfcsMq8NOKDOZKEBiNL1ZbHfnYI4GPp3M5CyuRTXYTpzBwZ6a/Js
0Yn03dvd3ccJqcknndeYAUQ29A1LTFXgUqTmbVHaG6vD12Rcq6G7IP1owHKwPEdfIVPNXKObGEtf
1ZeYniLJo4CcZLV/lgF/PvWTZBGQLJ6VpV+XLKGnbyRRvXHzloH+5z3Ws0eB7g+eAXdf+T9ZLJMo
5NCD6QGept5OgmYBMelbjGf9wn/Z8HRVy9wuLncrxSVAX6j372S15Z07VXG/MB6FtEiTLiB7gCqR
TbLVJM561bEN7f66i3QXAR9J1GWBqbjVlHzWncEmtFINewkiSk44NnzvDLgHH0XnzYHrEq316Z2h
xEAYYLdpP2drNCk8/AL9Dt+JZcSTLHZCA3YEzniugqGO05RQSMa5rO/IecoyWs0T0WQ9F1clkIiN
L2fjTmKXBn2GmCvWWnmMdyVvxeleH/Z2oeqQKBWWUyzg7wEcaXvmNleB3esWa7sj6pUWOnkvxi/W
SmcF1Mv9x4TyE9KjU5tknopXnZYE1+BQk7/802HLv2fLKF662+gLMbqVmUldtAYRm7PtY4GfyuGK
vd/7Eppx8udvl1/1i9PuCQr2deTTRZ1i9P5vkjbILjGNUGQpfrpMpI5+BXvrgpGyByhWe491MQqs
wCqo0t2d9Hgueq8WCB7ch9s5I+aA0rCQLmuf2Frb1t4CSybiCJAhdOFhbJ/aFddJ95NDMXZeMtx1
F/LWchbSxlXDnryxb7+Puz0znM7rrF0s3UX9GnjbprYOsJdKeIolKtODVnsPC7fTGmB8ohaEzRP2
DnyUyTPBK3+cdUpakQ3VRcW+W+ZBBB236cXH68rYedMiJzQ8oOEsicP1zfqsIsL6aItRbhd3rN9J
CTmBGajyy5i4UKLMdhhaaMw1w3Fi4FQBNAaJ+J0gL0/Cl4GumBenLeOJnuGzjMmqwgz+QN2vCtyI
Ro/a3tMBleUEScHHYfDY0D5BzKVVlLHPmb8HUIbqYRHInV2+81tEYUZJB549erI1MFYfbikywPzI
23/BQq9rWdtM2kRxW1yuE7QGsXezUQIEUOvBnBhuIqdORrf/OJShwCYb2e4IaYDJhqYh1qzT6MrH
fnhBOZcsoVpYHEFry8qkZeTUY/sY9KyaZyYsrYxTog50YzZejOEEifENvYDiTyntfxvjK5QEie3f
KZYHjTzbF3wFvmL9JRx9g2RvLXkZKzJaWsgFsy/swNaJljhGPbnH1HNmVicTXzbPdtjSc/rhBEiQ
PV95evLn2P758xvxZZoAIUnl7v7t1zj2DXP2W9GQHzDIEbD11IOkcl/A6O++2Ny2jbmk4Eg+lPi1
0eqcIVE1SwNDWAwxkFkWakyvtmytIfcpKPEvWL3F4FUCxzndvTbLHYcOG/NssnUokAMyKDpVt063
Yy51tko/b/5G4pvb3bcQvdQhGXB68GcOBilulaXcwoBMA0XvZRxpMR6VWJT8rdMHpHo2EMfo09XJ
XYcJvqv6erY9FlnJN2SVhBG3YDPNPIUggX8C+QpnQG1V/fVbg7MI3SNv7ipT+UEDc9ja785C/k+T
luo7FZJxpQqAdo1H2NIUOj3pqxacPXkw7NM3V/jY7FRizn2+g2g/JanQymsxzFVinW6LnbK4hRpB
ty1y71QNRdHJXV3zFss6LCQl1g9DUVQgaYQ9utlrP0SDJGgunYxKoiKbktDGXijG0noPwRJl9z9Q
3HR/F81PyfQUqh+WvGBMYKqdRYd4ngveP3XZnjyr9/tGKYEZZJay/c8fnd1z14lRGnxVMzop3y89
vyCgshvLpGLIwRB7SENkCXwjZR6JwDGU8n1qVDVAFyXYXo3Zd024CVeay2omiK0ObPkT83EeErqn
JETAQYFHgFBL13oQEMEWbcV/b7Rjo/JsBjkN6Kbl9EWR3XJl3GKAcbbZUEJBUd7R2zEjelfMGK6D
Wv17IKEq9t3HkD+0nMjrev8J7tBhJyo59xzgNgMSH3XmLeBwJGuJZojbvTY83dcGDqh4v8oTUBFg
qIPPw3TAM0KD+gg4ybLROhLV/NtEhPUfVXVLaPlWc1eEFvviN9jTEP/UYnTC3WnNASDmnmY3+Mik
E9qj9UOMPCTifE4UJ17WiPcx/mahFR4V6pIUGVotsJAhnVH1knWNqBFrVSph7HmTp888dlCfplRZ
9yyCRqs6Izb5piCmQQ8ZSS38/F7I/mRb3ud4TK7uyt4ARlurRTKnYZiyDuQsgUNlshaCAvWDlMRy
BWBsqJdZLW3KZp58LPZdhVSuC+3vSMuHPE02tpDxQK5P8+XKIGp0ACGtZ0kD77T33c+lp9Rw6SBQ
Pr13hmf1WqnZGOnd7d3LalL5NgEJLEveCgMvMm+QGdOiSb0syCexdDKNlZeOXyDKoH39Eittp9Re
GZaGHKNLb5p3ZU6ksTosKooVkQuJmT0LiEVvrT569YwBpSv36fKauJ398n5YKrrlR9HS/aNW40s3
Ch58cRzjR+6pSP8m21c9fMSOy5AtP9PjapGhSiVyd5bic0OYXHR/woCeyKMtRBxqkBysA40tvnf3
izlKsSnm+YWNALAnViFXwm4PDR513dhr3Y9kb4KMsKDqcMm5yW5YMsOLgLgTYlenlBIhyVmwKXUw
zhRb2eZhHsyFqVcBfavYdjObO7w1BjEv8L/5xDXHCxxsO301FNNKohtsh/ySGOAa9U1jawkq5+ub
VipVlWmN2kbFXDIoL7j37hUT4tmHtDsF8fmSloOpg7NwcPRviHuOcwz8rlU0CFdkOfclev9HxwIt
mDH+xmg3wyCvuZNszWpKTpOGWTCY24JD7msQlfB0RHBexDrz58KF1RL4abdqIQ4x42mQM7eyf0CF
7NR5lZMif4TiyjQw+xFD0zmWv9OMYEsG6d3wC1IS7kK8/bhyYOHXIKwlXqEuZaB5G6umOBLlXhv1
Sq+I5N6/e1TR96SWOdFKIwJRLDY1zSHdbkL/p803+da/5nmDqjoCdehweZ0rrn/FgA1vOyWABKKA
Q/kvrg8cI5R2U8i+41kwcYdHX6RH+MuH5hKXvDWB9LydqbptHpJ7+oe4zI/PGFVXuVAbQdNY8HW9
yySxuiABqzld7svIz38poEyDvGphv41l640ljZVKGHEhke5LvPFBtTF8ddg9pFj0O66Y7IDoRr1x
fLd9tXaZoxDETiS2kzG4f+CXg3H5NFMzHzAHP2Z4SwmV6Tt3IHfL/3lIzfrOYVkd0EIb+ZVvA5p2
WL1iI3U3O2eNrna8rqNnLK9guuER30FHqDteGmtRiXChXQeMa2HULJmAuseMRSF94Wuq5buODUqO
7itTsLkQRpsNgKMA9TnWAyN7TUd3yOLtKdKQHFIPb4NS8T2ZXecqWY4e4zI2JFODwagPVAxx4W3m
ZUN3gqgqx8bbQo5A8gZoypw3G2ReFcIUBxZQEHEBM2gNJ2VZxMseyK5Sd8UWr7JLiBRJEP5gyC9E
B8/xT1qPjpGKVOzr5in/zoxmhiEV12M9yOOIm0ef9/zOkmX6vjNl1bfiMvn605gqG+8yUzahfd/S
OJbF8Nrso2wZwBfQL8RjNPX2NbSwF9RTDGQiVaCQg0b/3ZwmQMbZZb8O7pb3DYHr62nFYDWehjg8
FGBKyl9X1VeC5GmVpNZMmSUu84gON1EmT73Bthzf4CSnbJl48ulmiY8DjE7KPfAdOyeb2raaH3nt
0K2aTTxfFmfaf5DivtAuJEYTbhVVnEoJ6s/sn2QBKaXBpMHuoNPBwCC8oHYdf+c0p3opYhcfZ7DP
0aLo+xX50o7tqE7YyJWhm/AGBmmM8VwjrysUSRCWeKaeHkozpZkXDrDhPgykyGDR/3HoX5dVgcdX
ydXjopOF3kguBhaK4mrdsbWKw0mvxDgGMOaTU1wkBa6NL5olVVCR4bDnzq/K3Jy2FxFOomC7zmov
RK87PSQKLU+eEEPv5S4UyLFDxSw/5iOjXKUAGG6GXKQLnU9yDkcBTpWEzkGT3gstn4EJv58zpoVu
U9+DAUSSCaJo99elNsME8AwEWyU8PUt8Su2ehYitnQSmS45fnsQO2wNy0lzTP+s3vJqvrZVmgczN
yRA/2ATdwMGjOpnqN3AQjHaNgEurlPZjYbYJas9bq3M7f9HF/GmwSjOHZdrX50ZIZKezIAnQ08Sv
QHs0nmvzhJmRYGuMbrBTiT3wO28A3vMgBKUWPpU9Bf8W1wFzkAyM2Y3toW6bZCxEy3dJ6pG0SrQb
Z/nq1901+gYEKxaW5Rmi3JpUIXgApNgG14xcp/Z1JwaJtz1PdfVAU99plPK3Cr82YAzVzZS1lt0f
7p0AoA4qqdglaW5grMAG0pz7UuelYem+RUQLjsux6bkKx6llmDTT+LQOTkaXepk58uOq3/uvqWEo
aUu4OUHqWWwSj7AxJBeQObZ98twxHM5BuUdPj0j7uR23xq7y7KKp2EV1eI4rEmeZk7KdFQatO/eX
+2G8dkuVZwybCWZc+L6wT5nLN3MA2+oXlbVmI0MVPj103xaVElg5hmo3703k57cgcvTmXhogHHAC
6MDp++QzjRE/u+d7Tbvwj+qFIg1UIcSY23sJPOHlfdL1YOvCIp2wz+NLqpsd4+Fd5/AnRdYGH1nj
SB20VY4iql0Om+9K2tSikjUNhv6rF5km36IEOe11GPNCIqg4u63Blj6x7YcJxc8kL+mlO0x6vweX
gFYFELeDDs/mjdFMMrsjqm0Id8gOD8oLZfHzUyBhezyi2EvCL4MoyRefBZnKrmI7eVbtdV4hWVIx
+qFZ8TgOcsBLNHkmat8zek4tx4z5c8qtA/skH1FR8/FMellr61+xohkSiaD3/jtCI1IEHNzyMTG0
ljYqiLxo0dUvPMaQaexW2jsgz8Q1zcHiFM76AYnWPhYKosnYu9Kgh1rHJWBv/GtHQgbF9FJHvdcC
MZy0ufYDNMirqyc7C8dlrNA7At/3u7kerBtHVSBt2jFyAihSk/0NE75dxmbQ1pzlbkVv8AT3iYiP
gqrnkGv8rZps4hnLb5d0Ml5saPc1PSOQYN80TFoIY9HY9HSg4EgNnHI4i/Exzimf6/sSJSrgJ+If
OAfXTUwX8R7FuD/4Bvwsm0Ib/ZXzVq9IqxfGLpbW18pbbKKCAXHNHcQqPfz5wyK8YXDJ5EthsYBF
36sNX8y/YmAOrO4WNoWzRvcjoIk0WkbcYErZknLJMTWN7MBWc7Narqmw8JGm5vYZ1NIIRxBJdZt/
tr/IUmGokaNr9wJQOlKxp3AczS0vqc9m2GrOsmlBWS5TiWU7LbRni2zKET+knlTfLoU5rxtNkZZz
rsQCAn2/E1DtzLpI5WCyBjb6c5rDS+UGSJbdNz0VfDiw9/9FjxD3/UWwy3nZjslHtl3AuxWyg6/G
mKUluUgaav8IJryRE5Es27P3KpsAxcKg1fr/Eb34c2+lKGRzyRahGEoVbQs0sei5dbtFLyIq4JOd
4rlgr4E5G9fBXCn1f228kPm9dML2hs/nb3JBmT2A9j3rWGBtXUTGyOYM1tKw782isWMSl/W7KTto
M7BfOhZVWySsaK/jANtocmv275ngx9mDv43sWCZBPrzlEeg9Njojp6eHaMH1RtUCIlY3XoMgkTIJ
5G2HKLGv4+gv+Tb8YtIUV+0UMvHqP+FajBcIcLAGDUEY27OH6gDwjIaQp2ARGjVSCsekwryF2Ud9
oX4GOxDhSNUMd9C9cSy1K2fdpkH82OX6MJTOIuqmi8k90qX3F+j0vQ6sR03OMHIeEFfd3ZFrDx1L
nEd+g+Q0wkPoAxy8cIVeME8pTZqRQIYCyaJLzcPw3AbTObUjekSL4LN2E58NMmL2Hhzf5wQ1XMCc
b0pOjMCrqK4fjRE8xvE9pfnKqKPdwWsDj7Tp3pHEPJwOKD8ijg1CFSFDVu9vGFlFdFvYoXbtsQH5
+AljOiGFqvY/IJ5gKNr4tupMte/CQcXDrf7Uyzp2bch/9qw1OSI5Lh3L09dl+qLzpWFkxr4ICd7p
djkm3HEhZRd5EhwFkotJkdNyee9/XwhJjxaarzQASbW08SJXEHDgnJPinKCMsXabg+JBMBRATvcS
6CkQjxNnBZdD1dkQt7PfA/rnqsBSvQ2RsvBKrXjPFSB3jomssmsNb/pi3k3V+6LMG5klZk9M+DM6
k7lJNg+Ju6bMBh8HDy/AZ5iZXgIPzslofLyZ1V1VnCeIjh2bqVN7vEOS8Hh4P8n1eoIRuDzD9XeH
K/DQDDfXwEJAHCxQXBYYpPunLLHSMPskg3YK7FSp4AGA2u0naIPQjSb/p1fce0spHYgogO+xcRx/
SRR8doOEm3LCHUat6QlZtfC3XCJeBVuZgXKE/L2pHzocjOVJpcqyx/d+hDnyi4z+n1CZAR2Hdi8s
eujwSoLIAWO0gwGnha4BX6/UHu20m0Nbyv15qVtcYCj8d/whzrqM8oXS7sWLKWkBQ/FV5u17Qt+T
hShP3TLkzzmcSTV2xK61M1+K7QpTd+k+VuBR9Pa84Y5Hyu553XCnP3SE/u4Ul42GxDKkniIqFkfg
GHCmtrzffhsV0nl68S/eKuHISPDglJeh/TvL/fcTN+wuZ489brljSbpcqyV5MMnpQ+BiA8J9Waiy
SR2ea8JRDrbIVrdy8gr89xrlaBKbewHAc8ccd0fEyoOQqTZlFiGb2pgVZIi0FUlF1/eJo/Q3FK6N
4dowpV3ffcP+Gkknu4Srn0vfzuvVknWEVTPESXOxSPmuUeGiIcuT0kFTMi3fakOVccQlYEpTW/ax
idDJG+BFWr6xBl0MqVq4QSu07cSsBN3S0eBcfSnDTKLjpnrTQgzLEJvbIgzJtmeNdmJuAArv81HM
/cjLNmWT/Gb75FMJapFlX1WVRK46vA/+udK29HVhYXO4dojObV/RDurAZ2tBiEwDzy1AXEotF8wY
FGSWx0iOGe99TBztdEa8hIejcmgY0v8jBlfDEdUCiVoC+05777KqTjOa1rhozjb5SqMbyxsGWRls
5qpJAneTH1sdbwfI2qJWq5x1OBx5Ty7MDZpZwmHkcYZC5LPJVXXdeeA+jT5WQd9UfsF9O4DRN+wl
CR0+IuXlB475cGR76eUZ7nqsssXms9dHnhsmI472TL5MZMJwj9BH90HM7Qlmkx9a6c7OQVYQ0LSW
jIvuqHmt/itXXgVk6ZOPHbxnk1GmlG0oQDKTL7dwv8RpAjHVplIYPsL+oJTCTUPOsZq/u0tCk018
JQHwVyPTUueNleGO7FZNg6y0Jw1e877OsdK8OsdaqT27IvpMCyGZZPeuVZWVWiTgz4XMNUEQCc9l
MsujNXHBvBXCntOJ0jQEIHv6/4z524IaXjMn5c5r8q8ROjsJO8DWjFj9z4kp1qDf70WuZHI2GmCO
Eual5vevfTs6WXY81Z2MvOIq0Vb1yULRRaZBf/9ITmkCrjBxxhPB795NZtGbV9z1U6l03vZ3Ve6L
OdlXoEZyg313SO9VG6S99qmSNZFVJfAg/zRdaSxFJpPh2M7S4X49aLuxrxgOxopHtmQmjgs376+p
/zc+ZQtzqbRz1H+B7SVrd1DVYH8E3XAOM7KjEEAEHZLsxMa1RuDLdeNGu7+KeCzF7jUypUXj2yVq
lPcjrf0XsXAm+Y2/hemlQd52mQ0H+npyVEoQmdczDKGEOq2yXXYH6MgIXPttQ+qKj2Qb/jPtuKD8
YXcIruOMJ2hT3umFNdIPprVnpSevIzKwpNzmTykIkPXB7Y9lVsZxOmG3iaamwl6pR5FLrTD03bRv
od/mAPpCrDL19pHwSyCPFEtwizGmk07h9l0y3K6U0/56z0fKcFAd5Ei9avjFSaBy/WAr6BGWvkWw
ihzZew1X/9QpoV4Df5/1F0lAGh2ef9HNb5ryz6EjkoGyOtTKFZ+zWS2rd+kjR/2xbBEoDMUzFtOP
wc/1xU7T2bstaM+6z9v/Yh9o25gRX4/SQqkTfbfamR0udJF0JCMYaQzdAhf8sPdgonk/Xg07KSNG
f33yHmMKO9+kwJD3t9Esskn2KhitJKprd9KFS+vfyGNYY2pAjCwWzPrwbL5yNqWIH0M/kcGL8dPT
qpnIGKaVa7K+HsSkPdWjzr7Sqe2h1DbOukTCqylBYrEdNoTZuVQ18vP9rLQ8x1znzeCGORTy2RI1
oMxVBeWF44IAcyiMTgCjOQ/lVuXua7DQK6S5T2E6UnKlUcPZbAQUIEpgVEjiJ6IP4NAzwtl/AYho
K++y4Lsk/nAybvVTwuc4OLTBttdVOHrFm86rESpBCzRWH1wcSGEIaCNClOP5x9WnEUiYdEN8X+jn
t8XAW6/NJ4GAzcPkT7RTrVkksTyfNxVwX+Jogj9GUUo85VabDMQ/mZbyefvLzcFsZUa/QLTboZBj
uSHq7TY7/svnKVJtV/14LBFK7nhubmjAR84+A6idWNpTb59D6/oHVLHM2VvOXXVyRRKpRmalfw8a
YLAJVCK02XYMuekmKPEldUHgXFxbuJgjzh/RlDldiaeWA7TdoRm/snShqUUTAMfjxpr7BkMOmk80
ZsGV5J1x/ROIGBn7bW+Sdf3/yxPyPN0QyrL+cJMwOgUYRTWkUGvib04K5J0Tn4AA2n1ob0PSdtKQ
A7y1wm17p9xi/+XlGyUvgSyuV2iiiHKG/k6OTVvi9x+6bu+HY8/EEa1+0+AVwaqQM2PGl2Q1ND/u
emoIZvtlgPUF1S8x3P0PqCI1ipDxkWZ0xt+LiNk4YXaOr7oPHp56XymrOhRnQoQE10cdkQYdVBwi
4AUB0m+G5eT3c8hwIajFXAY6q4PrSdsH5Y5V9BTvUGYHJmu/uVArDvV/k6iD+bVmU/i9ESvMY/fY
q/2uEnI1zo53WxryWuz9Xh9LkDlnzKQu2Tdif4YGqMMNvDgm2eay9/8wNwDC6+8loZ1vyu6OYgs2
vbZw6Pm0OJfvR8Gn+wRkabNuGRpEyGy7peits4j48RpuZlARfW96+VzfCppwIinwCLNpA+citC8f
OoESyLw+VuIdewLpFcHa5sT3KZfb9aFsW6N7pVfue9TZlY3jhHc1dsyJjwjIVZJRU1PZsACHUdDc
x5UupGNmYUNY14bhBhJHa23VXtixb0W7o+e/go0B/qd5zKGmguScpihvSUfLwBs76vLx1LtItETD
SAobj168Lm4QjmbFIZZN3oEdienP15tMYjQHapX8GUJVyKO58LT+Xoe7UO2SZDmCQd6vG7Tv+w/y
e67ncrJYj5kdV+YH4WK8Zuk2ilHErk7/cWIx4xVo6UVMxALFILKQzuWUEZueGtXalnZtiqkE64Qs
34bkUdclWkFWm3r3LRHwHLR5MqU+qN4k2zvBF1ef18yTzNyEDGBFX6HA0BmjO3m3kT8BHEB+Yq1I
vdP6g+E9USyFv1Bs3dJMk1iJ6YGqFhWtC+xOhDnqmYtdNZDuBjF84+bqzuZS0Ssa63kVlIxM1PwE
WJJ5fmE5T7joHxygCn0sz1PSKHUazbjZT2hdFfUbuJKZGWoBDiFzHm0zLG3arNrwqFMo81hfRN8R
aDmZup3FRRwCxsdBVG7lATTE9vITLqgQbXcxXCEE4jdFl59Thdjm7vVpRyjd2fXzON2zY4tLE9BX
xpzT+UNDeLyp58zpXSV0KpQBDDJrvAvbfXYmAvxqZyw+JO1Q8mYFWiZ7BjXdf4wVd8RVHA8MCT5n
EIN/Fm4uzDaho6lsiww+fmXCAfZOhLjF3rw+Cie6o6s8MkiUfV0O8rd5vipBiXBdkbw5Zt2niqTW
kOQOHhk+K3ACsAOAa7N2f6sNhk+EKAOyPEfSj12lGWTqfCm16Bk+HaLaAv2kHDxiH+JIqzrm+twV
Sr0yho092jUdvrzqmbV5b0RgtOCLniaW8augvLLtA2N6H5hsW5LVAAxucqjn/AHdRZ4GMH/bl0CV
HKAZDqI0IIYR/4P77icCGAbXb030KAR9hLzxBgDGAOhBPljETkqMpSh+wc3DN36zw2m+T5KiGmSd
qvxAYD0W2k9EymptDr5xmSesZ3ojnR5FoIWEPilkaEWhTwi1nUYcaH/c9KPzrHH+auRcQ/hfpoAp
6PjL0+tyco4Td76MmyPqJjB31Cj2whZO9DwJqu7vzgNTZ16xqQtjf/2sPKroTAWtk4L7J9qtmjT3
Y+6502Yg4aGUxqms1uL+6I9+b80U0dLwxs8e1UyMAsctGXaHhFWnm/8osvOisLKc2uYiFF6FG0gw
AsVB/mpE4ZbHbjcqAhiHIOjqTpOtfTGgfNza+sy8vUH9WmZtB7L5T0WNS8XgpRcpvI0MsQyvLjRe
lkCSCpIe7m9RU4LsFuUOdExvPvApk1gPX/eqJt+6mUvUts2wOw/ekU9nowQQDzzMRHaCyDS/m/6F
bjXICFIyEkEnza5gpUyA2vwEnXNV9aN77UYwQ+QchuQWLpchNLlYCdle+arvqci8dwbs1aofAtW4
jAcEPpC2onuKeYYKYG9mRGMb6WYDQhNwCoY246tNjmq9zN9GRpQ9XLX5L2SsRvkia19azMIIkw7I
fp8cQjLZtgD3OtMPZtT3OdETXL69PvGmnnYIZwvaqlg+4pHu1yvNJ+H4ELIicNiajy4lHwSUd8UL
/hpcvUjU9ALta8bUdhOKhh/z/pEjuttOnKoErufZ/d8omaLJQC+mcqS3d6SKJwjkeDlGvepteroC
MCGec7uVx5jFavAqciso/1v/7/ALt/a7PqNXaGzkvNpITJIv3doeFam0omeigO08SFyv4gL9DPJH
vgDp61tHqNLZffHKrY7nA8LomgyHJCUAOy1VZkcr7rakBbf0nXz6V4uI9iI2/U2vMXnA3naah4ny
481bZDC3APY+TwxW+IiT6vlP9vavqkcoCvk0TLj8WjxeaUuflbyzaqIhl8OelVA+k9Aihe0QK0bt
60Syl9xtaxAoixZDLt2CtcBKFPchoSTqqSdIxQ25+z3d4sry+3BhR9XoZ3bQ/fa1sJ4yDtz5FQ/L
c6voR6UI/iaZkxsSmflA42ci5Oj2vS+NSuvCB4hCU85M6FBa9paeSTteBkn+f9x3LZUZ1PKoYTFo
IFakDf0UW3wX5dVYzUbpvVZwvuRBAv6aT7X8ZxcipaITHUP2YfdoS9vg7b15g/sC9L5xqJzrYOf5
/JHPcbGrFyVJjJHyFX4XPEJJF99jzQxsr5GWFjxoH8iQpBXmZSPrMFEXMXUWDvkxMjK6M/ugkw+k
eo/L3a4iI91hCFYPZ4nuZoYDKv6tU8U0JIUif1Fd9d3HOg6f8C6fq3GVbCnnEkWDjsxcw17xQG2+
hH3lATXN7PYvH1fZ7qcjhRsr5p1nzMizWX3zYVn+056uj6COFkpULkaAtPo9zOGO/hZNk5GLLqNn
xlNPV19Q/nnYN/FvEP6lCFRoLIXSzpPCSCQsl/yRvYtKiUKYVocayaDSvPlo+udURULGgt3j06VP
Z6JBEARafozM9NLf1GUsD+sOB9tzIsxaHF2LJwr21IJJGm0oo1HRtL6uqckWHRSDzxlHSZe9kEez
8YOjFkFyUbKxZJ31y0cRo+Rkzu5pfkEyF7oS+b7j/+Wb0rG8JUc0vLlyNmu9qQHRwIl512h5KCo7
SvJYmfYaotmLC4oVSkmfomN1hVvrLMsYYIhH9UzE2mS224gMoXNGV2g9YvBKQOX6nqe+dNFUGLOs
T62RbtAAfpXDIYsDk/774WoGCBNAFwjKQZuJ8rZ/Y6MH7FkL4h1y9/MW+sb38pUKo+QsBl5+SeoU
QoPDJdedJXQ3wI/HQk51f+0RiQm1MXBqL+ucDHa9sdAylc+sjDuOTfMECzrZ10q6w8Sad/vgeFs8
vQkzPXAaxbkfZJ15AcMNGpKHSy5qCeDLvZA450vzG4ixFjr8i2Tuon2r8CQ9V5pJ5yXpRGmxYVlo
LrfMk5Rqp1lRP4lk5YLmIhF0oNPzg9hqaIubCLGopecB2rJKiedqAKiW8GAnMB2bAbvs3NhV6nF6
wC5AurbV/1bOPjRD5DxaZhKtAzVaKpap4fYgQkSffOqo1hL85mOQJfKO5nYEx+Iz7GtoeyyRdsan
nHOhLgv82xZoAh+utgEDLnm3eF4M1OEptnX3wI+Qt2tkv5y5HPH1qFNk21b1xy2si3FVzj9NCwJR
dzCXd6w9gaD7X+oOexMC1sMUOaHsgjb/IYTupVKiAYh1ISOPD+vLc2oCAqbQqYBJY+tPesL2ir6X
zyYqKIQheVFIw6D/Fz/c82fVsaWEou+mzDheuDcMy2roSpvKzCaw95l3bZXzb09x+6rG5xs+Ap6r
QmuNUXC4FgbpMhEpdSZVAXLM6dZBLw+d4l+53/anGOiOZMIXQCfC49ezxNyCBWzB/mm08B1ty4J7
IurgmMBJmWOvCCX9nEg5iR3XnBX4+N2ha/W+p2hnDdTMhiNviDqNNgCqc4m0Q0fyGp8EjmGdueGT
q95ZExF+NbpJxgMRvyJCte14Gye7tJk9hcnb9N8HueqD/e2VPsykaIXXWXb9A0vPTEHmtc+du4Vn
OmAYjhgApmRqEcczGRzUkhgypsF0g7Ir0JPnJwo5PKBdc9LKF71HmXz7l92miU2BNAaCroG7wf+i
lQiOfg1ZAJEZ0xe1Jxjgi3T7vcUiW8yYueWs6XEEThXyyGTlTYUFdW0LjPI/an/6StNw5l/BreZG
CwwWpQfaRaFDjtjRpkMyHv8Jd32+ogEBVL6T615IkOr5qla/LuLiKR55EBa5QozyFP2MV4VVQK2l
3lWrTntsPpGOlJNASUsw18mMXhaLI5ezPXoVQ427OSGvKGjv+rRMtxVGl0orh+YfUm3uY2fsAhRb
xXKOczc//BcAccTE3kG5S279PblHTjMPM+U5Xx13h7AMvylaQWE8XBXO1mgGAyCQ+fGM16w00vhE
LwZ01YItcTPTRkTd8JpK9SRg3YW0OhXZ5WH41BcfKiCmawylDjd9q/oipCUvRS1kN3HCRd8JKm6E
xK5Zy5PCZIWFlaVwrPi+rMHaqL78Dj0plUxl2/pS6rpF9iQgOMkc2sf+7slQiKENtveSElANaM51
EmNRfRs0VaGRJZX8ebonq/T53EaLA2+rIpoVW5KeBUvqQqalz4NiqFdIeFyV8klm0+6kc311Ld6k
b8/wBaXvKoRl/iGp7mHdfhHeubZOethO0zFXN4/uxe8omC27KHLuZnujPID/QKSarpsa0YJUZ73q
pZj/wQ7Y9jewDOkZtZ7trmGDLiE8iukB6z7P4XX25GoUAVJ9jZEMkwqrg3IGvLF8McOq4spLdbgH
9FI2ftFT28JsNXHs5SAd09PGexD0/sKEBoGLwHhEfVCQMUoyat7r1X/kB9y+grJX18W+ANecWkgB
8F/gdwpa+hCemdMqe8YSjMRcZBREpymULqwmntsSOpgkt25T9NuSqL2lJavFs6xUY96BQx2KoiVL
1mZgKve3rqQKzronPghh/suJDxAFKyNLf4DQpDIvqv7paMxjGIvCjjMlg4tm5JHImmTFftOvlgCW
WLmpQ4UpomCLgddWkaK5cl4ReJUrzqxRHDVy2KjxtFmqR0FuRC2hnQmKrJJ3mxi1tWIk/pdErMlK
+etIfCn8tEJI6H9sBmyrOx+Rh/yl6o/GDaakNmZ3PXbThJCUkQgqELX8NLwKcWmVhPKIzJoDFTuB
nZDRYBzuPX1/vSvOukHP+/Y0AYMbTCPPEo5X12CdOtEAh9I1F7m5ePY3vXt+6iZrVXqb/ky36ep+
iXDud8ZJF9uSKS4nd7MsfqketH+bwb9qW/Uz8euz1Y11Flh6aHHvIc7HRVR1/VkS4uXGF0KYU+b1
Vm4ffwq/LFR3uTSK0GXoxjCh/O1e5aCZOOCiCriC0BAxg9NUiCUrHxx2YTFhAX28Y0TqoafDQmF1
qAXYuYlzDv2FRbxzdWdV6yaS82Fe3sDYkGPDbKCxzWx4ySj3ayhcN8nFpBrQ3VKqWa3OFrldz7k8
nCXGq4V+kP5gtztg/5Oi0LQAZ50Qi/OhIS7a27bAW3uFMyFXZQu/qMM9MONvOC2XOTKdi1jA5AZW
+3Vs0oJA7Al64A9izWGxbRUc+6vmnFTIJWoig5cR1Pjg5nhcras3OltmXnwGkS1CbafW0zsArdJ0
weXPMw0Si2QPs91AzqBRvB3lk5D++3f8nfabfVA2uujjckE89rRSRVr01SyO7svMXT9HUPLvBzLX
tFM96N4w58Nj4CgntWrQ/RtTupZjXtjZxJWykV1wbnyKYC42M8XrGtYHzne+QesBndDgNntq2hMB
PH7JjWVwQkL5tjsRtf7//qNe3X3DEhSND9DvcjiZm0SoD+rSMp2S55V+pvJiBV7YiBC2qEc7ERrx
q81cnSWY4QGBAOd2kKhXKAx0bm0Qv6uysZvZYvJCUji2WsjW/W7/UVaszDtMAuCpS6Q1ZbpM679q
WRTxR8hOKaBEOHgeshDDWKuZJ+PJL3s1Ydf5YYt7FDeLWho5DFLZLlOnHJbkJL9EMvTWQ3Hw/r+G
D7Gahbal/W953bJd7diOGQmSNcSnOAB2EJJuB9oxFdvb1XlKZjq3X9l9cspzyL4nrifhEIm0znJ2
MqouaB1b0bbHVP5rGYlNEjQUyG7o+U5EuL0h0ENROA3xf0xZ4BZZqpVSTFJjciGCaMmcY8eqNZ+L
SwNeIQbVj31MuSLTAf5qn8v5MRuXmoPKdgcBuBP4KaV2Co6UKiRikDNCI9dVyZ6KTP9tCf8mSdRq
+7Td/ICw9N3bpHsEM7wE30xXGrkcbcXl7BphRGQXfki4C75TkO4HartosQbBVibqg117mgjyuES9
FEXZMpiGaffEPUqhHJtizrkyjrLALf1a59raJ/xjXTAmATaznLLp/mpC1bg0qN745Zpvx2euaCKU
VLiCyi8owJKTGzQBdcGPoXpV6iopvZ5c/FDOmcU0tQNs3S0Uvb1WXYNhckK7OEwO52tcdHsDbara
ZZ/Nruef45/0uHX+m31OuQ50D89yO8WJDEFaeQcZCyYuHBgFGd+eP4NOsSSpWFrLccS5xvENgnvm
468oY0DeMfRR2UIzmVtrMtFU9pM6BbS9SxmP98l8x5wsoc20CYzPeXEnKSvqNPvzsukefJ36LVDx
xDE3CH3WXG8GcTbFd53MrSfzJmeMTRnPwtvucR8YQrRSJOh1YMSWFUHNyq0d+UM//zGqORWXeVPF
/4FqXxgG6/HrCoXulP+nLppiPCed3IdybgUHX6lgx0CWoJhVcUrDlaCX6aOeROAmlMFfyv7PVCTx
5Z/pnwVExEKfuV0vmNk7vvVWhv4vLlEgbBWcQAfj9qMkYCQm+zKwJ1LnJjj6o7FlHnaXgWge9k63
yakCFZM1bcL0GM8zw8Pcjp9B4bKTsQJW3mp+Tnz3Xjw/DTWeznJDG2smbDwzgT5V/AJdazDhLmys
XHhWudT65Ym3kCZk2bm74/VrKEfEAMco1d2WoE6rDVqM7XefVd+0NIRznLEBUyLEBqK0PyvLHeMS
kOwoc1Glcep0WCLJ+m4TARmJmlPIOgbKe1oZF26vbnnUmZNkVegcJHmiC/4Uq7lamIhKFVe5IpWr
O+QVoP4rlGm1UYg9U2XIm18nYnM2FtKbgccxiPrAy6MEFL62mP9JrTBmjXzvKTtByzlVKG+k1tD+
ldJ5tF3d3dq6fjjHGrCOmVcpgECom3TfdqadYNBmMALf5OG0qPXOyo2gh1w1mOHoXzjF5pLAEzsA
pLcX6g9d618cwgcTwfoHZQ3kUyuVvAilcWttvos06Fu79lz5P/RQ0l2SrC7VjpqZklAxj2FafSMp
OKzaQlswLphq8Lc6GQQYuLVYRCY8zxuCpuU2fMK5O78NZWdBbiI6x7RGYouVJ6YLqtxwbwLyNWhZ
itDr4mPyU4H8mnqfkVB7bFT9jkiwNP1RWPgOtBIDwnTe0mSAlrJ2HU0BQ3+gFloEJGcqpOQ0oh72
vE7h++rBp1a4kMCnXqCdNFz3y9wJDd7etfk7xCFwh7McT23x9sf8xh0maPt23adhQNTDX+Cdexny
DoNNRBos5ewQs5UdlwqXHfCkJ2EGB6KypHcthfmiqqtYyKHz4KJtfUnMK/AGDHZH8fW5t8NcXmFB
ojnNdfwHy493AJ3vjtJbMQ1US/KNEGBVmdqOozIEOIDW9x/jeWH3BZcb/ABIl8tGwOswr1RCDLj+
qQxAFApiGXJKBjB0ZDIc5vFLC0o3Py8+vDJAuA13YtuZeV4H9iKWCVfuavMQ9Cd2znGZK5Jnkjy6
STbvwH+EuAcLjlyhIdmQl3dfTblVu3d9ZxBXjPR+e8cQF+3SXB3cOu1hPAUEvrQ4CNePGNf/yTyn
bXUfXcEANkmUdhjJ3EcDDo74CQZtjpXb/iql74bqnHn/OYxo+7SFOBp+LlDhyD+NRhD1elEFXp/c
xyVZwvqHpKquQsG5nFuO6KjAqPD4HkwgnwuvmwO37Ujo/qSKo40eCYdvDS1BRY3cjALohd6EJYQ7
ICIYduT7NirhMZxUL++/8yBP2EmZW8nmvIHPVlvq/aFUs2vJk1eEKAS2CKHqj1tRsnbSKVdTU8De
AYLV71oZnA0Z8np6krN4XVGY1zVgUDzW72buuAubKbsprki/3BVE6IeX6TgUGgWSSiR21ZbUqa1b
rnLcXy38Xwq5vAvuSRWSfkC2M7W6uTNSJwL2KSiLwoYdZwJ1f4DoG05ddqUo2OPwoef9CFdtSqx4
N0ODYVD/6dP9OQmDpzBiwFZmZ+iIxpW3zR8XI/TVwkJG11vIix3qALWS/0gM3XMosttz8OG+xPIu
wwnuA2MvKMFM2rbsBABFAo3+EuE3AgaxWe5ALeS25Eh8ljeotoL4Hfq17ba10Hq0tZxnySW1RDkE
7QwlrtrT4ErJqWz7ieAojlmL8uyEBE7XXUG4kM3SIapsnCJtJ0w/MckDj9N5EBzkAyNG5aEmEXxV
9BYFPR6GBHlaJ1Hfaqo+ubYTnjIrB9D+IP0PYd4WUgMCOOfyAHc2s1WP2C+GIhi/lQE97ej19FEu
X3FDQYUtYJtVF67tmA5tUBK9h2oc4JvlOIALlQbz+p1Ww8jUrO7znPsAMYZRvQFsJ7F0d3ADSjdW
tvcGpBj8xXScWWKFILnZ+jjKhEFTerR+2v9gmgb3tvFd/3NbhHFwSAkwD/7TfdH/5r5LoIMK83mb
PnzGFHjauOVCZdJrUCvcA0Is145rJ/uH20sX8E9Rxnz3LgNlapqddtdzc+O5PDDkOAuV1OB/rbe7
ieWSDtC9AnZ9GCqUrU0JSQDPdGpbTEojBZwiYTk5lLhp0zTYiqtDXUwyBLUKdQUOhdzx7t7Zsevf
ngYlFcxlWXY//xgJ4+QF8PH1sNFvaJJAKc3lPq/rVjfQwYYluNAaqdnL6h2cEYYOEXtC9aKmZkR2
0h402yi/9kY+rcjT9O3BuJpx+mBTb8EhEByvF3N3Xu12z/F5xdKLmsa5n4yJWFiBYH41pFLX10UB
Is+qCzzCFb7BGo8jcwgQaEIsEtZFb32PWmh1xNLIEGn24bmCtgSEYTr42zEThVWPuqsT+ztRVDcZ
o36hcWr5pIMIU38Q/Xag+pB7pTuMsNKCjKf5LsocnBKL1etT+dS/WpFnJZJ+w7vOikK9wS/VnJnC
urtsnU90q9M4LInfP+Y4OUn0IMBmH0qUYyjwJKjazxkC92CMORBjDfy9tAi+X5zskhYxfCJOEWeU
Gk03eCO4LkfQRm8mP8WZPY1aMEtHNTpK+wByPD7BEFc1V6ZVmVlqR1v9Kf2BT5Nb3k183YRLEj4G
R+Gh1mfgi33FCLiENBwuMya5Tdks2YkXGAimcbV9xck3TKmz0dQQmyYkK8hhv+4Pf2nnHqOicCh0
3lT5r+oqLyZmyGxOANppbaYigqRRF01CgtjpzjS1J21BfyZ9kVLFRkszaYW5rEh0laK/0z3qPXMX
uIN/7Oh5rLpWnS3cY/Q2kFzCTka0lgvheWJ29xLj7roAv6ez1ppnbRLNt9BdXTxSCoDc+CYuIdEs
t4ZUVyCARU30xP6DtHint01lUR2OeFfPlQRuGgb0hxvNFoT48tXo1Ga2DDt9YwZ1tVbuLvRbTB0i
NSHR/i6dHyfJusgHPKF5ZZQ0PfZCBKOV+6fiaTDiBNNDB2DS0VBXvuifZ6ey22i3Q0bkc43vx0Ll
4KjEyk60Q9Wj1qxBMkKsfsbPS2fRuSOnf8XmSw65F409j65JOLDAHKcDEOQ8FflL6S+sd5UyoHCD
3bBkq8djE1vN2vM9Pa29E/8C26HPNsVT0hxwSmWlK+LXbwRa8tx69NMiQzt9OWtdV6gBYurJ8IqE
HN1hfU4WCQRTzEFtbu9cO8DNAR12gY3AAj8mqWKzNBmMA4ei09RK6Ql5Czs/+Hp2uALbKIdSEEpk
m7iISVLbVpRAuTC0rt3YdAnfahE2fWxS3uK2CUvjLLZi0rJWVQY0GLJt7joYfVctRChj7Y8jNbZ/
jAtlrB6K9WLEFbZt0zPtKcR5IV1fKTiOBe1Oj9CWvnBJL1ya32ERHL7344NvMhhhBT0jP3OTnbFp
S4Q1GWxRR6hxnQLUtWmWvpTs4/qP8JE3FkLtOign2FNpAFA7a6Dq1AqpdnsKwfflagtXEOWLyrzO
Cj6GIFSVNjRXo87I8yJk+l4v1OS0F3lGMcaIWAdc6sgUCArcdtb4socuiuyXHClICxjzLSXIcVsZ
4c1WwMlZDlEYbxxL797gsbT3TPvp+HZGWnf02X39vfbMev3oRo1bF7xT4DvT/eQuvXSPMr3kJtUN
rTAo8TF0zF4Zf1eEGMMx1hwGgcpHHWCZvGMLDVzgf/OE8ITLm99z4DEyPR/61FxJ0jKdzZBguGGL
TjCGzSBNOROtKUMfEP4urTsE8enIo+ESlQ8yrSnAoPoeGNwWnT8GSKpr6awI72aHAueQn352B77p
52EOJ0/eCZCP/3P3E7btE6gV5D831nYHgwIRrzgcYFnRf1H5c9j+STLvZ1tO6RNlmDG03+74ppi6
f/2a7TNyn2xH+Bpsv5HV8JAtmCXPClOxaPLpJrrzrt84cxHOUqL8231leuH++x7rPMYUp+Bxo6Hq
PZgbohXxcs6QMmnNWfhQ5joOpsjhPMBx67w0nthrN2I/KSZfLg9fci831caFuCa/jhRxK3y/QMQi
QUbxusxGpJiImezoVYIXqXvaVqWpyIHVdIOdlvuvWdWGtt7+Mr3+6hdEimS0vxyV7Sh2ltlX5bbE
kos4G0QqsNuMWfWPIRA5p/4Dv/nbLZyhw4wbBlHdn4t8B9MCh4c2iwCrz/ujK9kzNWl50sP+2Uvg
17WERM2it5ZQz//ElipnMEqSmZmo2egpsDQ/dInziX5mf2Y/aKZJgVM09XtxmB+fU+iL4MkCgBHt
Cwjxgp+lLZJZVUQxd9/najB6kEAR21VhT8td3cf8agCGJeq106wJQnVu7N6mg9CVx/hKzxqxYuww
SVYCsQr+CusUvyTB+Jsrv8+/gUWU2U6LLlZ/VD5JSgboXR/ERLhwF3bmfdCYiY2HUHJa/b6MAr4Z
kEo/OgcREYOKkYmINzyIVkBnGynNi7/8ua+jRM8FEeMOHMVz0uFjCjdQzNmr5Jamhi6YsMjeYSgh
kdP8DB0be2zFrck81js5CCbh5lPPaZx1H0HobPCSYkDR1bEZZKfqFHPZBG8WCdKiQ5Ox4RBwJ85a
CYwNpEjBBPraxBS7NWgC3bmRkrbeyURqllEXkqr+x6xJcka26MFL8487hBSDKKgPbzTx26tmEiA5
+RfkT2qjp0XbIDcJExnptUxu2+GxI1+3meTi27GiaM1vI+nd3LVlCv9ECe1kE/CDX7llM8kPM3Ge
UBoB/rzVgD25yTWpaDJL0+FaC27+RxY1EVfRkaMwZTS4pKSPTbdWn5DtUus9GlPWzcda0PBHN+Zi
TRT6fhldCyx0xLJ2TLE9fSfvkMHIioL2RHYTEhZDVNezbU8zqXuAYgI1zDyp4mkEhMTDc28spm28
8YnPuN2X4vis0hAze/BGbKDiqhXXzXVn8OE3Py2hb4VQVoaOdLD7vaKDkjY9oUFoeyXzfHl6Eo89
yFUhiwX8Ya57FcRxRJ1e2TFbIQouGbYWnlb4bnEOswHxUDlvp7TMYywTNAoBFQ9VvVBK6Emi/END
yHqqAi75VAq2y2TkiwS/2vO4vMxMkl6uukZLCdKuTwbJEm6owxFzfA18f1MEFqvf9Ss33HXDYSgD
z/UHFKjAc0buj34ymrWEYvgiKzPPeKv2MdLw7EM0oplwGGqwgqK3HHCDuMCN9e3kd4UZBVlgeHgU
PuHHGA2oQw3OpgR3Z94eoIXOYMzG2bKRNV9xVq+cNBOzMB5OgOoNVvAyVbQUDHThMt1vkXlaCP3Q
rC6/HaEcQUXnBND9cCU8YijLcDYq3+zh7cp8htIPTj+HiQnFD1zop3EdXY0k5hL05RR+cRskB4Hg
U0i9wOgvQA6ZHLqGI6uYLi4DxWTZootg/XUqBCK0xeiBAw3cKAiB0Msd8LdqFFwWxtsCI/pggRUI
hrXH4yyw1HpzJ2HO8LTv8FKTJZkJ2065v9J3cUhrJc5F1NGEEcz7acQiJWX1WT5dxbYOm0/S4faX
+MWkwjT58q858gGVu1WFxdw+DiTtTig5Qq5HJlfXbuqUDvjDrbP/uxpbHaRoK9vI/iCo9Rgs6m+I
9d54TL10uKh6PBaqUMo0ROo9/3zxFeqGtojQBVmnubJKGrNx7sUvOO8mtpmZikig2Wi9Z3z+bsSD
w44YL4XTYaJK1dfKB+uEB1MWwQD4B7uaORNFYBp05qyRsI5nH4ODN6LRCmvveoldD8XbRpg6kR5v
GEHzopKexu1x3B4RgOJWPYxA1A7NkzO/h3ZVspEr6WGFLKieQ3kLXbPv6N2V3VMl4p36pjiSpcM3
O1a7EugDgqwu+IaYhGtcki0VFe9f9HYvmcJsnziTrVGW95UiBo/mFYd0eKstM53fLqFfNbOXRFHk
1QI9gwenQzIeXz9oIJ0/JkoqneSdcUwXtBtpGK9zNspmCBp9bFQXnJU70oypRiwYOC+fG+pP4rh6
xQkRfMOsoNpYkyjekOGJgN/Ncqigxm7jhT/m+2gAsMH6jFi/CIrPidhpmzYOtQYDtRdjTq7lpBRx
M64c3FS+3WzO4MAxLiuh0jJEVuhq57RvtXrC6n08fCaGZo3nNYXBQQACo/+dXFudVdRCnATwymPq
jxwUVO4+NaACu9CkHumC51P8uXIpQoxhlkk72R2BjefIt+nJL0A6l2LDPC5m6/ADoEgr1H2qbLjL
2lcUT0zH+53pRU7qgt9YG3dLAUQiDPvAXc2VsJWaVF6pLFyNWRCy4xyEWLbbaFXyaP/T3AA0AeXW
5YroU/96Qfr5cMwFQ+aqNYCkJLEqhDfvMZxOaZ9Mw8e2/s4yRMFPbr/Zfd8vXX7BAeNsu9ebJHWM
zsUblOhj6TjrOhZ7rA98tLCSRh6zw2/9aUPOZBHNNKJwwer4UZ+1DI2wg8XGywVyJqZyTIgnt5MA
XJMLomWZOc9kP3h7GbrNi9qtoI5G0ivDbNUzhS1+He27m0uT2LiEzP4M5gRetAp2KfhvXHl8qwfu
p+uGgZ4o1R7zml0Cp2jKjtTOU5DSkNuTL4q0eLkT+i4W994/mqbjfNVVzvdRYdp8CULHBVsqdTs+
5dm4TFOeUrNfjfwYmjdh79fowgB+fqW+aUI0ibtOCDaWpg9lm0xUvmUGmCJFhqgKlN7mTe4eXPdy
H0jWVIktbDFlFqlkiK2KPkhkL8yWysnkOuVD+yBsC14h7sGAX4QNiVqHDkbUBuhw/Em89RBV7mVd
6X8hzFDitBFwfqiUnI/sXK1T02cDueOCtpmIMrem45senW+7QRoRXXQFM+VCluzzVEERHvKksXGe
dCqRcZh+Q8Y0R3th0cAv0VFF2ec3K8BJoo1eDz9I+MOghLioiRQdae/QcGJ7c89Oyx7kGw26wKwy
4gndRFTq09v9xohmM7EhRX0nM6qxPveR2jBm/QAy856gO+wslL8aYPCMnRz/P+vGD+qCSyTdkPN5
xPMt90Z3gUdq65jLYey/7k6w8wU7oQjP50KB0pjYrTibh6JqEwCYVpgITHFyy67vCTIEh4wDqoCW
bOMv9XzC1JobhxLuK1yyJU84FkI6YIQXlw0JAlvWyRZ1K7hschC0ihgokrr8HzVIXN4Ax5cKa+Pv
pBkHKCvuHjI6LfwbWaIB3eGhhKIwoUIXIN2AgXRCB2k5hwKgKvWccoZNgjkFG2gMf1n7+ENrbNyw
FxUdFezh1UiTuvKJcZkzXTSJEZaz6iKNbOmF6sN5II07jPV+rzowBA+B/1q+g2FwpYUa6utFjZHJ
ixFKupy/f4I/QgcVe9BWDceyrP+kKq1Ae79y7qG2LLh9yNAaM83CCdCfRDN+aifYfYH0MHsuaIPd
Cv14rv2XqXDsWguAbKh3KQXhg4N26i3p1BEKxDebJS97qzLrYnuS7TGcTbccvvhOwMFMR7YyGHQn
jNpkdyE6SCncfdcFNKII2M3B4iaJ9Z4Ohux/O+ngXW9cfe/0yW/CLRkZFdOD6oQoOKZvxtpRNvCk
ehQOWBVn6MuL4dEuBrn851ywayEydqn9bvWGT57+TepE5WS2o2CJKqkEYkGQaRjNKeU6vmV1rfYT
U6vbccR0WmlQCKmFqDEXR8t5cI7PczXJ2afUHqiaHZTXojBCx6Es+AgNtBdMwQBO95NZMpGPlRQ2
MsFIzCsTjP6aJTmnyRIHlgLxZPcu3wUNRlY4rcycLFYe4LW3jINDAh6uC0w1kP9FsQAt2WWM8HJv
KroeD8RSO0o0kelmnNG6r/31Ijtumx+od7uCbIPqdjaitgAsnYyOOhdIBRFMtcge/Xs5Ry7pALKr
DSQqpLdHKgW9D9b1dn66yjfk1CG42io0DI1hW3NWEe2/k+B69TfZR7Q4h4hcWAN8MrAluaikT966
ZdCUhE4eo2kTTV2usbYw+APsoCpG/UCg+FVKGCaXcLoef0oofTCwKKBlAZx9c02oWQIpUi7vQGUe
IHEqivgqLPiuqISNWmEe8e1Beg9He3gjk2WzciJFydEHNrHDytKl3Vw1whOFN9Ex+g3+IcxcWr8G
eXa0Ubpqxwzt8gTFsLrFwpyD1oX/OFOhscp0zRYJwtrpRXLj+lMD6IZwamZfJYush5837f5zQUwX
k5GXYQmxJpKZnDN4UOs4TlRydKeRlMvPxrdiOvNqdzHUSPm2rY5OXihm/o8StKwt37ufCW5s2pl+
sc0dr2hPiByD26R3JsXsocV8I59TEotU+UiJ59QklCLLQ3OkOe+RY5xvj0xicgqyXyVQDSs1RTfZ
Slz17ARJwlQQPviqWk6B1wB2z5sYTDplqRh0zd5JXcksNBqSjuVyUujj6300PGrVasLCKWO3x8t2
MZROxiy15b0vIuAncjkdEuZsGw76wQyOMysSGSAb5zprY05HilZABWIjVHfb5zPvaqlwBN0joiQE
0F6gm7TWSHonw45gnL27ZJwd3AmVFNPpiBErfC3ERQGFYgkCcv68slbmR71xE2w2pRtujL90SQPj
H9W9DrbTybEdiJ5/hspoV4y+9iii7elhBE7g6TEHstMmtQkqI/8yCvAnQtSFSzJVRV/LcA3KIjz4
DxD8kQSBHFGQnfk9b6O69ZcmgOkgNjV+Xg/47UCiM06rq5Ek5U3a500eh96IDvhGDPRBFFh9tJv6
+BnsRWv1x7XOPMQbNyMJwt1VzzTKpB2XmhrTlNkhfzsr2ODVNA3FB8JEmKkj9NbN+PLpRIWzxgtb
7N4VQ+r/r4oBuaxeDEXPh3jOAHiWjc8RWKkk//PG9fbH3702I0KGk0eyORUiLR0Dx1HveIIfIc4u
S55WwF+3x6nv1tSwZE354gltLhELAkQ8D1xJvNoyszCJ0UuwEVVseIM0r2g8a8HkE31avvrzmRSy
MIkwko64Ecj6Sqifk0pNayOPb5DYx6xgaws40rpePJW1vhAflWTFc0W8m2dpYSRcxgXALhNNRCWC
aLO3Wd157sIbaSTifbos3oBxHE1QIGlS8bXooUKFz1t3OAIi/8KQQ6gzOPh7xlpBC1/8N/4BaaAX
mJcm5KiDRbO4+ma3WU4pn/NDYtIOdTI8MCV9fRWKAbi4NqqFxoAFHMUKZGwM7lPRr6lRAX4FRvyx
UnrZQrIYHQffhPjDtfjqTOmn1jdMYEzBK+nmAfSlm/V3XkrvNvMKxLMbzcKpb2imAGBzPWxuAGVA
9+e1qH/2Ovn5coDbyDR+nBywwRUpzlrx4lpZ8CDXPUvm/U4BMlIGK0IhutGTzaS8OcRWs3zfP6bd
VrEsYN/+RsBRlKXf4pZ38aYxgbM671x1IBeCZZUxuYtLm6OL3/YOO3KBub5uSh90IWNd4mSSZ3Mu
qN2XxDhSdy2rBRXqYgZkB/+wwVRpzdfK5RxRaH4L+Mik3kyGNY8mO6zt/L2ZI1tM90+etLKl4K8V
BRwy3nos5vd4eMUXRmlXU7rn+HIhApSRDSPOLqRwqSY17zmx6FHnZZ6mmJUFU8NZhpJyoFO9Q1OT
z5VT+CfdOD+IvOMvFfWvNbVBpcacclea+qAYY9a5dC3BOCJS2sgooNEzI6mWijWbanaEuKO9NMp7
U0jiCNZ2Drp0J3+iTpeLrfxxL2yTbAWWJEw3SmJ3EWiJs9HGksHs4WWU76fbDTQgV3GuKVABaTy9
Y6AxHuYNH/XKSC4mEfo1ec1iIR/HdRkVUfCis1gXRzzwqWJO1vWMegDJbeI64nJNp1quq66MdJQy
jYAuF6EjvDvGfc3rEhZqAWrbwrcQt9OkBO6XfbaDxKoWv/FTBSz4rFvRHvNGrbuYQgfDOppsoWFC
bvwuzOSzL8kGfp1K9v5mkiR3n0SZmcbwsCvpEsw7p4J1saxtGJ0POE0o+9FmNr8doKQFaK9AHRvC
6PDzWNomK1XGvxOOe0xKEI5H7BgQQsAXIckXvfWeZi8nr/cW6BgKI1qT5Ik03tzANKgO6PvFYRdk
oqgmQ2hQHIZt61fahy0kif7wU9NGzQayNY+9+oWt+rsbdOl4a0YHU7Hh3lap/4rq89jY0JhEkw7I
z0V0sy5vzuS0OFl8/Dys41bRH65zA92G9Qxx3wmVWuZUBa4QeH1Qia/a+ba84Y3BwzVROJ5NG8Dm
Z26XGl+I4hbUp1AOxf851FCa0HegTTLp+TZuex9ys/qgMc4yvXAINJ93U+HR0UfB1i7mdM5AWtDd
AniDFb1T0JbIU7V4q9nSshfMD4nbA8472pHY19RmLxkWrUirFtSqOpMOBFdaYbo4yCQML10/N5GK
sZOfrIzbwJ2OazeUrIKBZOCdyqGgvLDtm/Viqznh6aHcv9gGfygg9f2+ahOr/vH9i6mzKpm8OMiw
e1cr9iMup9RNbA1jhmG6wOT2F1XCW2kQRogx6xSbpLporzuNiXDuGlDsB5t/u8P+kaNDZwMIojdv
mwp6pNZKKOCozspmNPD7Xxor1FmqYfPLOaJ12BnNAGTac4pj7pmiTbgf/e1Y08n56D2Qs3ZpyrKZ
km77cX7ZbcWDdTx5agc7pwUI+O5gTcvf9MCw/+SdwkN4aAA1kv6sWn9/9HhDjUHbobnMP4UlWxJL
hITVapmeYUFgjOsi9k+AwaI33pfjXzMBkOl4gb0YOVC38afnEZHCS8lXfYf8PosUcU5iFmBEQWZ6
XbuVAf+QsJvleTGfMNRoCEaDZswY3NblJ1fLFi6F9RXYQAcZ9FT+CsC9il1WRb8VlWAbYielh6UT
uuQ5ACPJzpJRBHCgg2C2MudbaSoTAtAxKq6U2j65I3qCcJiZ7OdYJvyDxCEvEEHJ3u9BIIA93QK6
9DKyNG7y9WsmDE3q16l7F22aoIvH8Z2/UAlWquVBmXE31E1ad64gXILXPW9jl9G30Jm6Nf+g/+tr
t5xQIjdIohOnW/CXfbgsejcXDCDj1XDVxBYGnvQYtE27noAEAaILU/hFkHa0DRRrkiqeRVRrwgZD
Dgxxx1OqUxul17+wFFlvYD8m94KqDaXRLrtYUXkfhawTmYcVdYVSCKaBoibrvUBKxilhq5+lvJzY
vgMjv5coVXJR6RjyvzHra1DRF4zBVTx3GhXhwbG/OaqD53oDWNmgUC+9RQ2+peF0/Uf3V/8IG373
pJNbAJCAotaKdXTPQ2ZKGMa3Nk7K68vQ4LWqsOp8Aovk0oQO8ia7GVPhbWL/lJWv4e9wx5bXXAtg
kJ7zcaXeF3UaGPL9Syc0HKjP2drUDza8NaJh/FhBL979Q3Mtsjco4JWf5pDw1/cu77OrNhllzDVD
3WrGB+SE1fSzISrSZiMLLQD/MCTH+saIQw0QVfEuuQT2OiPKnBKnWM/4KhBAeb4IgkFZRoHxIPMf
dktiZb0KmZkiyN0FMJaNauNGiHrLH8/Af5rK/px1dXsuS2mz3i7Yt0yEiA54+hPM4l2dDzrtQefr
GloCNZ/tX+97ynI8GwSI/0xLdnWY+U2kCGovlLg1kE3q4rxUGmvzNVE4oytILtDymrNT7LdB2zPn
UYFXRIwiTP4Fx6E6aZis6tr/Xy4ftajxMT1v+3GoRdAlNtjQTIaRq8hnyiIySTdPsGakeWtAu5R4
5J0DXjYUNFbv5n09t/8gBjhT7XjORt3O/Sr1jTg8VKmSZmlkp2pYVaLZiK6JYbrpsZ9REVLUy6C3
lbufLRpOEEstjnFu656htyTpiIWSfNnr5w0qrqwOfYb0cHvfTbx4CbpKdx5YIJpMrFFkB2ILJ7Pl
ZvA25vaCSHl9/fDWQUMiyyBxBhYYQu/Jvj/B5B9+Oi2Ihd5BQ7lonaZgE27LwRYmo29j7QJIVJSS
LCqdsnZ7AU1RJSpqeXJe54BFB7YIeCQrfDUDNXcPJsD/J2oFXl87Bmh2f2q5irUtqhDgicVdYy+r
Oh8WpCWhAr1lBDPIVBSUYh/YGUwHfJxFshmymp/H+lbwDVVKS5FEpEK47K1SZ1ITF0MH/yNhfvAZ
nJzUuaUh0CoEkm0PNr1h3YlVHepIXcl9HwfKhaP6aM32FxGMeI/SlMY7VtrvSN0U6daCX3bspiPY
3jOcmCkJ2jJr4xwy7QOprBllT4zr2dM+6r85teUvz31BjwEcXgFFTODw86yz9/SLg8xVTBlh6Qho
LjczEfyGRGenYlmhc+o42xh2CBYYceAEBDTVzSWEi8pVdMWWoeN5ileGPrfRv6z0S3ZUi/NpBmXS
Yv150iTXEAvXv4gn+pAi1Siy4o8hc2jChRmF7xUQyVmNQ6Sp0xY8XO97Xp9mm62DexoRDsw0v5MT
GX3jY3+MWZjGF3ycDjNL+e1JCK3jrRngiz+V/EPgxqxLLMoflsv7s27G3XYYlzTMxi9Q3+5pwJtw
uKeKbCsnAlPhq/bwaYzhZCOla3WHFdqGCUZe6MKKIGwQ6OlK6X0czbB0FFwaR2nb2YxNkTsjlRZO
QMq/FSFHdovfVWGGB/miSRk9rNB0jl/Ja467yrmePANsIEwOjanzc9UvwSzRGc+c2O5o2xBcN0tt
+LFjjHv9TtK7TR7L4gydzn4fb//SFr5LCuEGD8zzBWuatcR77vEN+7oWod10X6HiWbSDW5yrnNq2
/hKfUk2hwFAm/GpjFaQrbAOA0DTyB1/zRsmtg52NlM1qGDFtB3zHktEtUOlJROg/Y4T1a9LEzHOk
8rigD215uf4A2THnasHupH1rIiCLJiSxOUU2Ri3r9W8bPxPywXfPsC0CgD9owQfK51yp++dXUHli
fzxBdQLqGHickRgy3jKsmQlQjABlPvYWSLf+wLDK16OY9Hp6hepDUp+xzj5FEBumcXLztfy8FwAk
ss1qjDzvO29kS9IhiECj10f0reHqKAnq932zu345/TzukgVF4i+lVGKosIVwI339K68htcHJOZDH
dmisYVv0K+3agEHjBDdu+XXBqhVi5kRZMmCFyq/psz0MEl2RI6K82bPaaR+4ZjoFrQItpolmboLb
GtpU9Sg4MWKbRYvICovFlLPsXNDSZwn3AZumIEd47N6d5RtVAo1IPbkt0VoUnv9OQDQbgr+wypjL
mwutcuXrboOVs0x0/yk/orghIPtyiis/UkovWegAe2eQ56O1LiJR/nxUsC8EPJ9vvlqPcQkjn79A
Zd4NM5ohptoThJ9blb5zBuOCLxr4B749UxokZcNeJV5jSPkkaditgIvKrQg8TlVrPe2hoIcFw2g/
fR9SGvL3Yr5g6JBC53PANWczT9um4/a5LDuvPNCi7ow/xaAttUJIMm4AwZdRknR9saTRVbby+G4E
fvIT94T1LEVXN70L2bCKX30ieDbikqM+BaLU33pwxvnKhvehEPgrpxG9cbXM2diBZkL4A+j/Sxzh
U+JSp5pLUnwccyJJ7mRouqYSKH3QlIRdb34hXf4hO+qLUa9w2Dt91D/O0t1g2SHLL5fyL0HoqBNj
kUHvYQA+gYUYqaiV1eBKT1UK9l10VR3ab+HO+drnURRbUa2/Iz73qJFp0kT3GApJmGegsM8W/AuR
CsSTbajkFRWnCKTcYD7wOvqsZbsJvNWCwRMvCu374/JfQWqBgX4z0qon9JyDYt0Fb2dXM1PPa3e0
phFjbOZsUdGkTDypr+u/ZUwY6aEPYKbPiOlyp4HTZFfwb1BpJkbx1x5yspJJFZVlGm0Jd4lyboI7
DuD+tlCiRqCpRvnuNMLNPxvN5Gdj22lphr47xB7FbjRV94uQMcXHxAr2XziuXgYt7N1lsWsWzAeK
q+8k2Hr0ejfi/Vov3ITnS56poD2Hs7k+v7x+14SPUva9VzBhjxBxl3TjzczQv+qXyAv0dBO56Jkl
zSmaH7ou25NPCyrQpJvguBJH9jjlm7B1qXa77UdwkTIdvgqiWWxF7ehC6+8Xtf0/8xpwUi1K6MzC
7IRvNsyiepVpTdinUMY7uRWTCgdjZo58a4SEw4hSaY3McKgbII6AFBz/64Eh6pLnbXiqbqEVEvp9
dx7a9eIyzS3TGLFo++lv058Ee32iKizPEpbU+ruikGhvCI7l/vJ6XxjCL8LqvizVd6Nue1cK+V4x
suB4HmkEyekjSd5CYgd7WGcRxk3mboYAuvSImHzZ+vEO5sKMCdeg22TN9qih9iz3a1LQKpgNiGCp
AE/SmsW4og76RlrkV9uCgPrHYQQeWN/VXn8EyPkm5xH3aI+BiQ1N/SDqamif66bsgnnIyMnlh69x
5Ean4ziw81XXTKo+T2HR22PRWwQt0CBbK8ADdSZPLSct7Lz5WNQa5t0+3cbWNk5liqxxYKSsodb2
GrNyIOjWouoPJwdCqnI2D5yyJvXWW/FFsICI+YJvDkGtPmJii3tBDEiN+bKJTB9HoUk8JkMau8/p
P5MSIAWpROOgJU8hd9f+iZbWi7mkJ1bMUk6HlxxJFrfrHKj6s2vYqAzy/x9ApsGGpDQbngrgOZRL
qvkqbt1D5s1yF2H5s6LPo+CBo7ykdAEK0HJ9Srm5YNfuKCG7Lb2rpWq8WucurG6Ve6lGG5frnZTW
DMpq5z2oDJ7UeZugiHvQ+5FS7ollI9mLryuXwxj0FcxHR8lDKxUrbrAbk0EOh36d3dcvYFbSRRQD
FideQMDhziyG0PyYu0DWxTVOloBlKLh2MmpswkWfc9G2lMPxSzInmbg5LWuENTSsKAV3xk9kXnTC
R5MRc3yThh8RgLds+n3sSSCVNAyB68hBGXHaE5uU9t7gc0kyXKSFina8g5biIEROGVTqaObVomjE
oErmY9rn60ygYg5RifLxpoa5hzDDIHCAhTV/1sLvqpDQ6MDkfQbl+piKi1N5Jp6K7a+fPfOl7Tiz
m2g1s2NJmf+t/g333TePmx7L0zYEaRPyO0LTWQqY9alindOxBvUrfrGdtqTKwcFush6Y5saSDO/K
PQNE3OB9iALez0LkaaTbVt+y/CdDSYg/ybY1EDJqHMcybQ6L6ghKNm7jY9wbfprJXdIMgiLXAD5C
P7vpug0H9nQKQyHNL9CZ9bzUEH4JK0tuLoYikneXyWijcJYvkCgntxDq9PSYCaNE+guGDNJxLK+D
hlinHntUs+LLoGcHLHNl06QUkdBh1BheNIa9rYHQro6ptSgb8qykZYmRjXv38AF23pIyc4ghEb2S
Ptb+gzOY89zPBv+vnGAGwWPZTb8zjqDaEKyruHcsUKFwpvcJ0s4Kp+qvSN7G5O3HyRK6uCHYGjeM
eyZmgMM/fxvZUw0tK/W45R59AgN1v2HYgQq37hhHw+fRk9haeB93mxvGHHBSGsDyUbLYDYzQCwXx
zPQ8NrFgtcoeNjS6Ss7KIOkghaV3xuJnaY2FotL5cwUEESmgQOvoGqAmGEK3xtTCaigjlaldz2WI
oMdz4nU6rT391LbOgDxcjm9l6a+PSt3XpOjIZLVmbCQIh6Cl4way4j8/bk+BIoPUh8s4E4HlrI7n
FNII9FUfV2w2/NwuGo97ket+TyR1s8fUL3cmvhNPZJAbU+WxP+7fNiX1uAHZz0WSsrrujQXVRmHi
n60r2aQ7QK39V1P5naoo6Th03GLtQlLKUavr2SwkoIBavGlkwdJOOvMYVOlLwKMlFENxdVJaHmFb
HG65F7+Jl+FWxVNFpKbYXWaH6XMHasCORBlWbp2IDjCbL3ljQM9m3MZ4prsYVHmlmuPNd1XKUrFR
oBBZ6zJzUOnwBo9K6hUrE0hGy31OMmqMCjdc9rEO4c5EaekAHYUvpo98aVZ93z10IVSxjh6w3nBz
kxuokChH1TzNuVxLO4CtKVb+dJzVcrMnjzUIURxDDOyi0TWMYlLwjWVlzR2H+kFC7GzkmPhkByyN
1xvcod+50FTP6ONN0HNaqO1i1GagOx6Eurkv0zUQ3P+oXsBhAdR8w4w/6S2Pax5lMucWv59DiB9F
ueOsWCGYaDYjXGLeNEK0Rnx2FRbe3iERhGEa0Ta89KqxnPR7Bm7bmS7fJhHk87KiH0wsvsvKNZ18
BhoHiCMmnXjMNIIuJbGUGfsuKXAYB5cIHfGfLVRpp7SDx4A1cqRQLsY+1LrouzAisglGZfNRfZNs
RiyJRsjyfyG1/EiWdX9T7XNlUltlVEhgzFtygm06baP++sxRcFvw/YmYHDNWbIWOQZ6JBq4uJUr+
IZwCcMzN0XrHEPUXQEtQjQ+PRe0l2dyPkCpYh7fRRhajcA/3KkeeVBKRTjXaE7W/EKdlwPReR1ez
JAYWYHsvtFLpxPBNhBg1m4igI6N0D4Cvc88BHCjo61mTKFiyGPFASWqNQgY9PM1snZLwndTSJAfz
kWKeS+gnkA8Z/XtrEnxPvcIDZKjnWbVQ4WyMA7JDO9GfK8zCqX3iwUZsnjjy9zGlO5kHJThYnLDZ
7iK3g+0kRfhyXW6iZOICgrrA8nyRSvoUs6il8gFFXvMx/Udl0xYDRc8X0aToXNn764OXrIWuGTvx
m9R8LHj+6EVyWRNjI9b3HvZ6kp5AconG71ZaX4/kt+QxjBgOu/fy6CaEdNJOJ0LYv1VtR0fEFhcT
Zj5iAmJuQ1rJfdT1CQxGkfzFmvFql74dDlMxsHl08ATcG7CGRM8JOnAHpNMYwn19qQAFpIbMNZ4R
M5/8DtVi6RHjAKQ7VuykH/9ciCdx9FyUCa0BKFl0nRo+nKbpFr5jNRtEWlnLVZeIJJSpRq4Sn50Z
AibJN/PUIBEjlYAsDYjV5mxJM+3Q4P4RpRXPKXX2TcsnqtY2dJEpd9fGRi9RhVvHWs8UrtELxKA4
RblQyEvf7NYDfQv+s3UcoCvtuicuyx9h7upSrbE9lqOMk3WZlG/uC8FN8eI3NOnWgG2k4MCoYsov
lPoSb9YBLeLbpOGj8pelLIaiBcd7VMEQBw1fONe19ssNo4q4X2oL6NNj46WRObRuBlDivcqBRDUz
h8lYxc31QMzh8uyQOpU9s2LxHJlQFxpMLUkF+MEmnFXBHmm3TbGzzY8Dpm+igonrK3BeZpRKqtLP
vmHsxAx518WDl/cTswstBxtx93WGrPnxA+lkFGxBcAYPuJQM2hqfxPQJcpU/bv8Rmo5fFIIkb+nc
b70haJkDsVll5sIh6ik4iYPo35TQFaoiMSwdApOeJTKrXvEG8cR66scyT0kG8nl2hsTKgcBKboKO
46NL7NyKg8ZdQwkte4QXSVsyEPGSkLQIp5cnFOGRjYUiH72jWaeb3Xu0Eyv7EigYA0mh86IyRXv5
hXhAS2UCgUcDt92h5wpOiO0b8f3pfydfbV3sqrHZ0f2t3htT1UD3Un+gtuTafASOAdMvHpIsl+e8
ettV6nendbD8RDV1HJ6Y+HC1c5PfL4EZ/83WOZeKKcy0CtKMjAovOgKbo6iNwWFlTSfYo3JCHBKi
WeY+4Z3W7lGrEpLItEhv4YATmW/w0c0HG26rtbEFDorniie9HxJVodRgOujCmVNaC8+CB2CQkm1h
bPvSlhJgcyy2VcIo4Y7fEitovBz8Mum619rTkiKP0bwRUl6OOcUMimrm0ChNZG4KPjVBybMVmwnh
K87pdAKem/aZogebwBPFLwD7dPaYMCgLp2ZX09vly6i0EZGiFX6am3fEJbdcm6b6J6WPQq16HnbP
RQE5+KwmSRe/G2Iab6W7qrihTw8+XhtvQ5vWG3DL2U/aCniZ7I3itQ1jtuT2OLUxkZ7b7P1+c6L5
HTZTWQqrNF96sPSGpsFRT67I1zQCirZuuVWptr/oiM5yEpCHwFjgNAytlQVtBpklZFypge3m/Rjm
tZ+tHuJ+16FKvgCfyf7WDooYkE+7fBjyTJYEe9lRH1yZ6ulO+S9Zg9bRMROVojLdmPGGJ9zJa3zQ
aHH7uQtrHB27fQOaux2aMt/MWU9OROvnmeR63/UPT9vC4igVnqLW94UPbA0zQ5vHtWTOUeMdynIL
uoiwG4Y1b2GjhRQkMO+0xV3FNDa2QM+BrTJ7UJlEHSEBZLdtzzzEHGaHLAr+o3L9aS0Zy3UC8n52
+D0HyabG22tGVKF4rZhoWM8UNh+n2tQGPI5URg+KbNCzhcyjhNfc+hBLuYzkn46Wl1ILn8hQMjtU
fZFvCABQwIpx604iwBe7YS9+BhSCjwq5lWxSQjA4zsz0XbUCiUqeXYbZaVBMC6QDxkYyPkDihsqC
39NJpHVzl2eWlutt6xdf9mo0yQoSj7si7WD3AQlQx6a8CExbLjLJH0zEkfZnL/BNpllnJNzRE/ce
/qLHjoMmNwH2OahFKlsDSmEUiGhnUZb+H8GHt08RJiY+u/bwkB1N/Zb77XIe9TdyR518wFFcyjCA
y687D+gfhl1bGdDGCtFrxqeIkEADIrs29MLwJgXYQZQv4CeVIexbE7znpPasc700ugDjXzYYN3UL
w86xa5+TElUY2Qcgd1kmZwwRd7Zux5o4OAieVZh0BsRSCChSrnXOR7xDYJFGW5+TQxf2UidBwDIm
os2Y+jY6jL4BYet1q9N29fm5TVuEG1JmRBQjJTBcDEuEo//2VJBumu2Pe4sI1ipomlJka6+8lERd
csU+MMaByBad2t6E/Yq5klxdPhCFnm0BZh3yWvoDzmOSEps1JwxFYF7KZ1JssWjyAQ+4mlIoxVxb
Kc+rxW88jril4twLL7CN73tPU9IKY87lYhzrq4Rx8qDy8Op4pUM7zEQI5jEL8GvTXuTs8nlOR/a8
KmJ4aECho4mhXt5nBGy2T79ne4vm5mL/oRcZcXoWL1LJcghOmGB605qnElM+sX9SYtYvjcqtDnrz
f1aWyc5UMt6HXitxdHPnz4Bv9Vw2ukTfvR6CRpEZ/OqeVnSclS/fFdlTvvAzDxVUrWXvwa8ZoTxG
nbHlvkXmX0A4RXc8i2JEiNmkJUmFVuDsPuwZqHLE9lm4MbkV/rs5uhjOf9U0Sc/ajQNyQvZQeZOb
Ibn8KKMlHJWdiOaZNAuj7X8e+d8ZgOaZv8aGti/eR+vpUdPJaimjRYyXoX8iQGKxNCU3qn117UV+
eTvvL21j2jlvGSHKj6+naOs/JzvdpZBz9tfjutTtGZszUZjMX0bUcmA7ML5udOIqFZqy9He4Q+Pd
qu3/ZKWMjyUeqdlh9yy+JFnpwb8B5YZRtXiptba+q49HRIv5F+ST5G2uexev5lLHDqb5dRqcoCOk
CzdV/oQXIpzfZ33mJRNwJfArhLsk7l9FX1mnKHd+jGltTQnU2JebofGw9OXMVfuJjTgOpXhxSvU8
tm5VMFRlpn02GWb5Ap3JzmNo9N2MdoSH4kMNgbQsgpDargDGSGLCIiZENMT0KHO8FFRzP86AWVeT
AoXb5tk/nSIgSQI3MZLEzcGA4bgZl0cX5eX2Wa9A3nnS6QtLKA4q+qc+U+K8YEhp1UEZa6Qo2JBR
wUMN2Tr7RRuIJTeBlemWD+JGdPnFCCcoWYh58crnnXxNKztAySz8WrzFyslaRtCyGTAHxi3yv3A5
W7PE9mPpk32xrXekRaelI8y7DgEFYM1vM1Jt4sCrDxYFZEGUMRYhaCKwFrBPs5PfnVNPdwLB40j5
7HOdU4PibF2PkgMAyfP/lhgaVSv+wW1Y36rzdKu+G+dk/7EgAPzA59bSYTc/vtH3FSsWRpW3nGNv
Ks21Spr0/frGYxITGYSvz3HYPigtfAu8W6UHERaYqcB7qvXi5rDVQbaggLKMsenhSHHxVNUm++Cs
oDVa0sL922wBNv0rIptZgRGb6qnxWTg6RxMJ6GNl/iw7oJchfkmCjion2nQTIO+K+EfkmgwBDq9U
KaC+HcKlDE8z5ZaRwZ9bFJxDEEr5F6A/+OesKSNYfhFF3wAKFcHKtKeH5jmlNXk01L5lLJX0gE+g
ZB6w+8/vgJufF7wtj3db84XI+8gf/OqEoWS1mdF9/+mzalM2Q3NutMG+aUyoPqyl1K6q53DewVT+
auQxeJfOp+k9I/dtgak8ZpPG94pbPKj/93oj+1/FTHJKd289QECiEOJDJwiJeCM3MApphluSMAvJ
lU5zFcoDnO8FIeoUfQu4Ln0ObL0B7KkdLZ4rXgQhXnAPRga6V6pnKjC/rc4GWtppjAam/TtNPMYY
FbPeBjNQNJQw+tEhP1z8h5gTXLnNcJFTRUwtBUubxhqQz2v1Hj5Fy4e8q8SsXxgjUB+M/wsBbhYo
MZiy+qrY9CuysGBU+4CfwBHkHtcVhNWYL/skOjylsz9O4sSUKFKz9u4dJxEjzuFpaxa6UqYDrbxq
fENJtm21XcGdRTFGqLGj+7KNM9YpRXJXdEe2dF4yBhdIp6qnrPZKtGViHpMmhAUdlJmU1H5llue6
n70DsimqHClR9rHCOiufyDujPwMh5PC9p0GmEWQh4qyEAGA2a0qba/06KG9IcwInMdTGWITmlqQG
6/TBnETEZvdcJHKI71wIMVR2c5ZI6APALmqsmb4Y/qt8bTJEv1GFULj7ugsPchnbdM6ISWbsDS4I
OqIRkJhGZQMiJE3PgwubZTR3HdS2bYu7oHF4UoCtPuxNSO+oMCm7+3+zFLR70Ma6dRxguAZqBmnc
QaV2j0uuVkBvRq15sPR9kiWggbBAavox8KuKSH07sVWMF6zUqegI85plhFgZqjyO1hxtwJ5asOTF
3BOQ4/punPIoZeoVCSGCg//Hc7iLKJMSmzyXv1zFojYWlQ40w6FejjB92bl4K5JNWJ8pkc5EoJxy
w4R3QLCOHFwSVT3xV846v2Dt9vNo2SgdyEIOwO5V2p9qUjJdleFv0t6ZlEUs2gg7p2fZ1FqBOb1W
klRVQdK3nSfyMFNGFC0YJEExLXxf/QUok+Q+idYotshrJnF2egeFyoYWpXkxUMjo/mXcH2HXundN
o6JRbt8htINPJuOyXM8/eRJhzQfvqlVSELdJmCE5/zMYOo+PtgS+wBmfNXU3ChgNYJF3U+w5FeYp
3uVHtw77ZT+oTeX3rFsNWk5GBJd7f/EEih3FWnMQBMSWP4woDgxSlfSyOIE1HKMS8NtkiME5MeeJ
ET+HX0oJByS3ckCrd1c8/h1II3439aYdOJpMn5xpHsU9hInv0MGFCY+GWQOaxtyRJcB54sAhaCkR
O/v+vL5F0H4q21EzlaMWPBmk470NMRh9W1bRvdFOpoR8BDDCQX99a/9LA+vxM7qeQRl7pVZ+4bT0
Ach0UOL2mvqCR4PFvzMtD3UPfe7fbL6Em9Ywft23WMuKO8um2ABk3x7GXLtM4aq1O69JL74dj+/l
kX7TJNj6lV5/OofBGaeHbcSthMjNt73ux71GEp/guSen0rHHsPkaA9RT15yP5o4av0549cYxzwyh
noldXIcdwjmL1arEPW/PJpz2QFL2QUn3am4LC43ZS6U+NA+FCUQy0TMZRsGw9W+jnA0VxhvROvFe
ZiOL3BMlgf44dZkFxRrxJG9cD2VZDZrqDad/eGoOhGJBQ6WS7H7qhlvclDxXD1lG0xPhjilsr0Mn
ALpNnwRHemDelW6iyhBvGdMx72SBX4KhQC0MV3pwwxviqcX8SCHos6MJ+b9J7ZJMpKgAyL6is5cw
ipZU6EzRTST516iJGGd8lISWGK02mHswJSwWx/hJ5xVLhx/0C1hg36xFQodfsppyud02RWm9ETRs
d3avpW8uETMWw6rSqzC+M3dsJx1Bca4JIFfjZk4qo7zVBpYszjhf3BtsvZyVzjvyrJjirn0cD7ST
Hja90vAZpHlE6mixHdqYgFLnCRlYfTC5xWfkf5DsPAaX0kNVDQejsrd2YH3sdQZNq1YWNTZUsajm
q6uys4Lt/UMeiw8lZ7VpRTuVd7osC/hG2hcfqUIamQfpJ274FkI6fThledjx9MziMgKyuAjqhOam
RYcznAyxBJ4r5CIN5Hh32UvFIfGcVw1qipzz/VpWRKvNrgapxsEMmvbCmABGm2/Ln9VPnIGU9Qxy
iK4ipCcjgPR7Im1SJ5sE7WfQ50OCZ4aFXOjeQ+JKbNp3rPgda8YA5U3Ge27hXiWFuPdXIuca2kqq
TZwl4NkDpLowOXefQ59cp6P4qfypWEXH5R9HLYi4p9QlEWeMa6wo1PA2B0xV2pIA6bih5JRNQ/+l
fzF9Hije7qx6/9woA2/Vea2igXY9kv0g+znaL3FwkobeTn02TUaKi7B53j/NyqmZbazpKhb9/2f+
Sp2bg8epISNfDFahGOMuAi76tpExWO4SovEXZ3lKVXLu9n9PBSPF3A1zVUFMMPgN8JBt/STxYf/u
VnRsIGpf7wPG3uXhoeNwGvvLvgNLb90u3xfL6prfPe4dUu46n1yvI+NKN+guycVxIRGhE0tEvLTT
lMKJdhUlYsRJ4eAa/o28FXMfoRXmpMVeC+32Sp0qNHl3z+QSlrsi3E9oRZBfjJgKFn0bBXJ51q3v
/nj/J+f0t7xOx8pPPwVEL8XG/HHCs1apyYcrVXvG/LLWyC2TubuIFEwOU1TQEylcLvkoof9q46g2
eZuaYNcfds4a2Ui8sz49shVFvoiUvLZzrVQg2W4QAwiaKORr7AokaucdOxI/slp5hyDO6sqahqCK
PQQTW6XOU8upDsKuV5mBQ25gAd2EhQ5xJsgxOFb+o69qgfW7pc50GxBNRVei1e6tWPas84//z6bV
WEjac4EhuXRnYqXIStXZNcrxASbAAFGqMzxLDskWQ/LyAUdiLBpG1bNRj9EfnZW/drihZB7fs8od
exYqflzr41owpEOP8m02YNW9spkXdNadLrsU4sgf9SurU92k9ZXL7SkuHGeetYStJDOyNnFtMb3k
NH9aIeVEThtAbpRjVWHBh2pxDbm4QqHAZsObtcQdzpQzsF574PromM0OZ8NGgDQO9qQrEpeL7zN2
iDswgvLY+X+OC/pzJDfiJBcOxC8mWHmVHd4ird2/bB6Y5s9J/IyqkWQf+1rYxt6Qjw1xYMvloOZS
cjKuse/oya/cEAC9veUwZz1/aFDqONhUZBb2ZNabjKXOneiKrw/D8Yfz8fuk3cTZTwHkT8W3WQL9
/OYhUifBBDH3p5p7KNLp8At7uyNTOxVqgMeV02+PM7ZLymvD2Bj3XURYiVu69hv/rtnEc3csAhDK
EGwaeb7EHpCDQeUS1TMRU82QvwTyA6jpzKAHGjo/lfQqJoaV5dCC3YylicSOX96duLyktsKkjXvX
/2rcMsZJ/ci9Xb02gbTmfFQ979FKpVGrKdBAK6jFFDlpT0rRvsRZ5gqLt2fmtACURO3gqOxtpBd3
xLOzgF5ENMgzCP5d7yXGihe22fJGrXFVmEIbLiOQmh1VlclV6/p8JCCtpJ59eYzsQwivwrGSnBhJ
HkkEOhowL3ZDA77Z/VD25fpKgKivVR9mYu/LZ2qyXB4SEiaNtmLI9vFzIL5IDMuN/noiaaQ4nOtU
OcKINaQuzObBKJZl4/pVSAPYJ8XuPHybbd8KkfvLOJ+bMwYm5fZyCg3F8vuxyWn2pXYL+qljQDMc
Bg3xgiwYt7zmALwdk6Aar8SDzsdbUy1dOGYxLSG7aoohLxaYF79zozXDFrt2lvMa8tZd0OUXyqj8
EQ+5M3Zv9pGhBmnbJnxTGa0d6D1wIpwpwysiV1y9BoEu5BnF413bCLInJXPRhSqIaHIhuAV0rCMH
9dzwp0BrUl+mnCmIrjWYchNuilv320ygtRTlBCPFbLBh/Kj9AxxwuXkUYoa7iZciLsY/6PrOZl2H
iFX5W01aVtQ8zZYxXqfUIVOhdCcuoyZ+K3T3jleMYUbNvVG0alsabowuZyzbb8uqIRmVW41ESiw2
n9BC0Q+/Ocdg8jPxY2QugBfJ5wSo30KVwSz1GLSXUrQI3JKYL/DQVD+l8SOsF0iIXsW8QXGb9jLB
0XffE+ayMS3DkScoXkhFn6a4l8LtqHZ3E6Un+Jr5PLqeCj+Doq3CJm3iJUPTWvnmnMvaBOz+yUyC
5GOtpFrc0t+0tUI231bP8vdiLdZbPEMGP8azkn7BsFoyva13UW/yCnJXRHY9lDXV6VzTTFmasfRI
xxDALNvYulm8YaHpaG12SrElCBvQm+T23SZ3oQF8MFHZcD0UqPWT8f8AzmyLR9g8kQcWteizzb+U
zQUyh/pSH1q0xmhmUAwBq1GEC4/axhlmowLCjdSR6Z33Ica3hA5GLeKS9LZ2F20O54v4RySN7owf
onpwcX0k/UcwQ4fdt+/3oqq5FkGDMvcRWkiHPMhI2D0UD51d7qxUGm9M+Nd+jisKGHdTAahDLqdJ
syNgm25xshE2Rj3aun9cnmmJc2nRU7WbO5i9Jl5o1Sqi3sF4dmTI6GAbUD/UUCpMvP74CnE+j5vG
vMxBs5S9u7hg1VSv6e6dWHm8LhR7vHjVmcYxB6cbjn75/V5JA02arGmkcGP+Ty171gHKwR4nYK+m
n7yCAYcVTJQFH11X9zUCn3pkWmH1XJw1mYDMZYiLl335uwUI+GLiITnRc5lu5FD70HYvIF+kWYP/
LXxi9GQcACJta0GRidguRdJyTWIMz09YyaO565YumyjC9PVYT3le5u+dbU2ledNU8x9rAadcQYO/
y5U1cp8HBsOaXrcnTSuxeorOcSzTnycWxRWDRlpre3Ae8olxZ+b9KOU+gZWniGCGpfkaIrMb5nVL
Vv4AZHjA00ZY3I2+vxvARormHNvH6FlF+uagTbJ/GsFkECuysZ4RTQ4Dnd0HQkWHZKQcYfoqU+vl
e5UcNl7poU4IJrSWO5Qt0BN+tdND6afIqJjk1rQwqoZRmewyDZ4tuT8dx/9MQ4OJjNS12b72biVX
35ENx3/aLyqUe1fo1YGoWFI1U2OD1ZvygXrodnuzVXsZJG1VsF2G96wr20ub5U+Je4zhm8hIAxcH
sxQg3fR6eMuNWT7IkaYW5ttJsFDOuJ5U2drZ9RStTSnMuXIUfPEto75abuV0c6ZTYUqt1Vut/aQ1
6zhUMC9yXCrpFDwUFEVGFwRs00xfkrz9GVdmUPLeM1GHX/uYC/Jqv4iur7Ug6c0eohvUMcUcNoGc
puNyvQMqlQNBpL7A/8e1cNJfw2jf4i4JF7X46CvTOGe8FU8u6DBXGJuDq8GGZWsvL1DBPrfbkkoj
h2g5aDvKyseh9pH8qi+/kXz7hzHvsX5M5tPFpa+X5pccWxXl3l96ap1sDeqV15T2s+ifD+44yL7N
Vbrkv9Y1iunbhT6eZ4rk0RWE6OqkG9hG9KeUa1QpbwG+jkJ6fH7Uhbs2kA13THQlq5mjiufZA1n2
puQbup591BzteNNXNGmzjhQsOXtrREBlSp1HGiOvP3FMKdigKuTX+KAoBxS5wZHcJR20XrFzmp5P
RKBBI+LHWbRqdI49lFF+D6K6ZmsofmX5EBnwg5cPNXlL3uYVn9k/TtR88jt9di9g67Jnz73MPqsk
9B8MiUjaVYSmTQg1PwI5WusT9LEn9k1fWiEwLdvSDkRhd/1F5r4taJGYEdWSnC5VNSrGgM58K+oX
ti8y/L4lGRrJ+/esrm+/mHHPkwND+GkkrO1ZOnRa7AvPcp6Z/kFqkdaO8GWmh4qjiDEZ+eOgZoIy
qdtMWqCwlNn+EeJDIvs/ieFHkIGPUi9YNWXakKCrRJ7UDYfBKBzhRFy8YB/N1N5Oo6/yK9XkO2Vl
lupv99eql81ShtFnAXjBTjJVxGlSmRlAQw6v9L4WZeykqtQPNzhbIKwHhluDuuP5zMBk69l8Xvcs
OfbuAOqhbwbS8v2l8RMIQd5+oY5t+2Rt48ApQGf2CauoLh51nCVNylL4MFT9c1sT0UygzRABWpbe
whz05jWcqN4VfxF7EffwY9BNB3Ba4FzRKII/Q4W9uS6nmNzDnk+FDgTUyodYU4AX7OY3NhWmPNux
w596gSaWWvBDrd43eSCU2Fhh9cafyQirhFjVq9ce7yKDfzVWJ52Ls+iYGqSSe6tHfT9JbGKQj4fX
D/3BvtNWpP8Oh7E7OggNcsNWzVYUqg6k9vWy0UUCDZnJQPCX5x6jFdha3GiLxPq55C0c0Ilwk2DN
1dq7R/jWlK4/nNZ+uqYIvZWbKKEAWlqyP2oRLZMxf5mIX30xF26USct26tpi9J89ZgGRfF3Wbdo5
9t3ot6jcHpkH1hyz8FJWTFzR5BCeDUDwE+C4oVQ2ttBYQlstsxSz345fHu7cGZ1xtdrKasOnBDvu
+WVY3D6lgLiUQBS2en/fZ2JbtaiGJq0j1RAsXwojaAwpypMHf6drqo4Ry2G7hxcPNL42GyXJ1ZYc
sw9mBRRXLFnOAfBzyJA3iDwrWkpeh3biGW/PiqPmqzU2gp5ylEwokDiKgqEDGKsaEJxyR1P98DC3
EXmUgWyVOKzYva7WjigkmwCJt0V9budAgQ4TK/hNaudQWKRdl4oFqOrUfo4ZnuwS2Kz6g0o90Kvo
5l6YEBE4YcwhOydgB/ljkFKILjpoPZu/UlaE8bprl81NIIC9u93qc06+oh4TY3QHEKoKqwaDEtBM
Zem8OGw3ESXoi6CEZnxibDM+t0oOVyQwjLjxmk/zRpMWktgrZyWJ8ibP6BHzxeqXX+0MWTs1p9bm
1lq7ghGnBBwPne59T4crvA0AWwNVseuVcw3sNlwtQX1B73XQqvPlYhVW8pdG6DGznBeFHb0eHOKk
uWUUF0BfnlZRbFEC7nWs61i20vDmRQ/8aQQtVSkyQK/bT4TlfLtoQmEQBQltzuh+qD5eIiC1h0vu
37D+z2N65xfMY3AsFbEu1X80uDYIqj1hjTPqlWzJrGP8FgFL6K11TRZQlwy3nNbzdw2P5gBlrtn+
eKKNurljIFVO0XAmt50k0o0LraVi4MS3i5IVv3qXm6TKKKqNUgY5aiLEyvYUFlJxrQMOitwJVLwA
TQ4d/BlH6L0FsGWzxOoPzqsckofbkNkpBJFNYPh8E5TCBgYuEOZjG7fZ3b9/bZD7OMmMSAlrk2VG
NihmZVoPR1ZC9IWciOe/pszsFDIeWaq/Mr9N/oTgBDmByQSs5Rs0sjVOYrH2s7B2YTp3cUgXPIar
e3NNGuSHolM6eHfoINik0sPA0FJ6tDzg/oQqj8Nje7SUharxRyurqCdFGCiY4B+9OU1OJOuaF5DY
VJEyAXBF0+mzjFvtmBDEgU7pmmBbHbYxbk8JsOTnBQVrGb8ZHLrIOhLeYHIdHXTDB6Y4Y4eKBd13
iRMwQV4kAMzAQuemSaYP8a44uYzYD80ksKgAtCFmazwGUSqzgXlX/zrzwccvIbeFM66xoOOgjp7b
C4CeX3asibSbYB6RELFWFllpEf3q9ViDNjmp1ilAIq/dkwNB4t1twOUlQCyu2a/DzEOSsdSrU/jD
ITuPC2Juc86/n94kzJOk9BBvmArOnpJYxnHk/foHmC/TsEs0rvnuylL9HBlJYChJBEfQQU890ivg
xyH9lNx1/0nzULNfIm4mZsIZ5gOWiDsdZqrD0mHXIpYfPNWxrV+776IVEwscfj1CQyxgrh0krCO4
mkz8lAdfb3WiHFRYy8CsxyHQvzZdkj0+0SR07na0Oe2Iom0xLEIMyflzBsH5gGmN/y/GWMhL2DWT
F/u+dbmXNjbLyZFW/XhJLdZ78QS892OpefVqJczbgIcZvGsw2TgmECc2b2qPcVsd9rTc3iYS+d+q
Pv5dNCb6Tp6wcXrpkzvPlGBJ+rkzUwj5A/e8MDTQeOPxReOOkYHInAnLjUj9nXC213st26rRVRDP
8L7oYpV80ei4uUnTY2ZfpPHElNQ+GJdHwIP5zeegeBkQynwXvtiAQ+KK2s4jIAoDKrHDYgB+UhC+
ESzICG8QMHHs3OdZXKSq8xu0L9n2cD6dNReEiN5WPI9yGekzZo+B1tPwyUUzx66drYCdw6zxSwVy
1bygzxNbo/aUfF3qxk6hz/UAb3PvYjBSt1YrlQsrz4rPENdotXXhBV284K9MCNUXCwFOh8gV8dHE
RtyFSCxOoQl9tSblFJmtAvAVN/Poau4EMX+mlPQ21b3nxmcTXDURcG9S9pC/LrDvofnnw8n9IpyJ
fb9NcN8WFpK7LSoa2QKHoIrlX827po3lDZi3/5gYnEqT7bX1a/ep2utInBrP5ROFF+uzzkHg4sMn
P0im7vAgcsxlhRs0/LxAZgeAJKqY1m7OXoyOYteA5thawb7aEZ2MQ0lc3UFEgFVuCcXraUcRrweU
rGQSCbYT0jOiBMMYvQw1++iW8R6gBvLkT9iKxbRTsivk+UTFJdl8og+OzVgSjOXI21xAfDTpzNZ+
D01A8lhKxqmvFrdp/APB1PeovwXKUXBC0GReeG/UKt5MRsZQr2oCZ5S/kDPC7iC2nK6AUJAcbIYg
OO97/B8/imfQlzXx64fOHafov6HQ8wMESRG9S5MyAH4u5Rpx3xVtq3fPS/rZ6lyAJAujiTgv54tM
kskm/WSZb1DJVwYTTpRbLLrkLuANNecnZrZNAZEQXxtDhhskK1WT1DTWc6M9OKl0tekxMiq3Lb9f
1ZiS+fF7xPSTLFK+eCu5KGDxh7srh+4xzB+VaRq0U4MkLAV0Kt4s0B/YIaFpg4Bfe+EqY/CFmISS
JJkb0I7Z5vKKWQ43G76RxcPYT5Ba/NTxgdwKWa7TI3uowE6xphI008vYl0cNFwC3b/NSXT15Zc6K
JvDV9e+vCEz53lQgiTwaV831xV/a+QExXBGJMUkS/r/WuNsBnWPxDf7fsoqAMdDz02QmLjV1Ig2g
sY9CMRJqEKHfGseinT+A39OWwlMIM+k0CToA6Sb0BT2UQ4bcHBnuZ6lz5MZklMmi7TzrqDo7GNdz
QKKwQVvPiCJacsjxFe16Gecx1xKyIJOHEn2dKmxH4uq3BZECdhpjTaic5pVtrgUuGHIMuQz0AQpv
W4oqrJFv4BIdZXmI0Ayjngnt9ZDHhpk7TzrY2aP+zwkrrLkrDtkRSbYvIVoTlte6I7RFD6X6FPGb
xLawxi3KC+DREFskcqGu9tr+FwJSp4FUfnzzwTPHka2jSUWfH3yt7nVqja2/nSVl0ks4cbzpgr9k
nJYPBS4L39OftKYRgod9bWbn+8VEMFgMlKT7vKrVxca8BQyvDS5SRCL/H5YhX/E7DCPS2MbxAxRf
mIvmdXT5C7J0awPOwtwRxCRKyrtKpUxL+JTDml7kzqIVaYcgAW5LGOsh9AzVfZBPc1f6x9EeVAs1
3PULyoBkm+7WTLTaxRMIMLrGSZ1syEWE0MzZxMq7AfSClJrsHomy7nPXT2duJ2DDhkUMdPQbEzYX
C5XIC4dGmGTEFoXH0a7t9n4zBHt4uCsMzwtf2L9mDCxcDaqMEsUYLb6OOa3JJD11RjCnfcXFDTLA
kbH1X6qUgFYzk7GZgEv7iKFNWvDX48aR/3mTxoGWZYp5y9b/OJSeRa3RbjtQRYtXYrxkOrRia9HE
2IzA334z3i6D18APDPR22kHBk98nY5X6QiICzMqyPhl8mL7V/lqgn0eGVR+kliJj+vvn6SnJ9NYJ
Lv00xoQcLdhg2TthvOxAIIrXUZxvvGnxxAV18s6euyxnyzYXYke3aTI1xbuglhvGFYadsFROpeU1
2k2jwtmYohzuRWyTLsjVgDnqMHo3u/scTzI1Csd1/rHWmgIY3rAOs2eCIta7w1yjdotBsc5Q1csK
13P6ViX5KhRRsGsUVRGBWPEbtW4BfnZnGIIKwSSvJrpESVLsvpYJZbYfGw2tXlZvP+/Z4U3zKp2c
sn/+GZE6F40OvGXPHcBb9Y1h7bN8OW846TSDvGnB230OQ9GxzTExmep6uulwwk8amGQfUGfTbC2N
NE/x2alPvmvYVk7PQSsLI+CI+iYxRzjp72DsgAXOEjlTxeR6UxAciYSqha2C4s9Tn6CqgZ/nrW4s
zv1S+mh+cd6DkaC6IJ13TnxaJbTyVxJi364g2XJqIIzG3i94az5ZAIypJbVM4nadmjFBnM9ZE2NV
zpc3IEtfJyrOIqWplFi2PTDX6b/sbylSO2hvhI7MJoGgyJD6k8j8Fa/ohEwfo/WbKTc3YkN4G2G6
dWNATmB3px02qxoNa52Zf7ypQRd0Hf7fmCMTZrTcLQkmvzh73y8U93uI05/k93fr5XkBJZtHSCsv
22MAQc5fxttzTGWmf87poD2lZ2/Ad2JFB3zpcbn2Yd+mI5cw0L6Z7DGmKhjMxbGofmtPb1jc29XE
fAyxvGacv4moMqinjJ2SXKyUgtpLHf5l0ubuCL0kGnhCeczieMq+NwpWNA12iKPjKSFnR0d9pqWB
Mjs0MQnbCENW74peV+oQMtbeMbfsnpez2zTVwAeWMgcblPf4282V8R+2x55pq+qjHK2WLcSlR53u
leZ8Z/ZMn0DbXHVDxWW+aQberQzt+fsWVNXkFNziedA4X2rODA2aDFJ/7O9DFATEqPnJaJjBeKAO
1BPLs38ukEfT3dFw+a9tKrzHXW1UxGq5SskeB+vGzU5OXuH4lXA+xoGZXT8FI3S3ZPOvfBHbl+LC
MARD0Ek0ye4Rh7CeYBacJeQMnh+079idnwLzbFxermrtj6FRBIndR42ekGgmsL3XoLm9Nkpg7JNC
FovUiSexqwkclbdhhCvnjcJ8BcLNERwxD1gtrzyAh5+t76nsbU61iSuXIK55hWFCaXDq6kFLCIlZ
lclS3vL9DDB0rMyEHPs0D2gc0o/oCmUdRdLvqNVosZDZH1p2Y4CbuTpf8aUWTkwxvlOS5ypHvhzj
TEqHyNKO/v7LTNriRLQDByaQQIbu/ultsh7+URINQS24j9HnUUyq/ZY10HBP5AekaH1qKqAdplPt
JzXbc+IJBxegKa9dPa83OtplxoxnwH+AJALXU8WhzLvSlPMr/M0lVxApowJltsgw8aCzG2iZUHbP
pviirP2DDn3t43Jje48RY7OHMwOTGcSNfYcNGvCcMN52ImGVz97NrzFYdR6//sM4wNY/4B5iNgOg
eELUFQgUoYmLQn0Dq4/NWsHJDbw8ytlwO7r3HFqM8zTfTgG+bS4Wy5ZfgrfraNaSrd9tk2lzcK0L
goi3LxzcytMXU1iYf3TmDRuuQ/4KUSbySOVZ1OFwQikcSGybut3kBikLQ2Yy8tMUzgMH0ets/iQc
XW11wH2qzWiqmeymMiCJuaquR35Lt0TfyFP+T9Dto9fYatf2p4huWfB5KDb7xjmegcTl7O3OMOxt
aGuufujeXwZwLQl86myzkWSHuwVqSxVW/mTBiM28MdUhS0A4n5W0Hmc14LPCwhpT/IDNarhCcoUC
IjictSoj/c6k78vGQr12fl4Ed0UqmxA5rw9pvXOBYzbcowDXwi0GYB4s9nb2tiHy1u93YCPB4NKc
ysQCZfgKUBLw0ZBuGAfan+sZ7mB4dyzvOygkRnrNlvBPajSPKJFsh4g4ThbEjZbfx6WF2mUOb5IG
9rH9gEtMho039PbDXcxAZYI95r9YECZVf0Veg4OxCVwBvRYhR6x1vkRaIKr/ntTLHWeCfmrhri3h
HxIikxSCs+4bMnFOS8Z+30YWh6tWhdwaiSaKB41BSZrF9PRQ2teap1HIR0EAbfA9tTKyTl48+G/d
5JuvRckfOfI7uRH3HK63tTPONJNjv/MYWpAvnAjmTyuv4zLtNWMvdwP/F17EPh+oxU4vHYL/3Fd2
BPiD1kJqes0mHHDhCS7TQP8IvHroYM2euWQ58FjjDTg5sDZlgyGvjC84Rf18VjIye0ui28e3VDH1
f1VYDl6GPiFukSi34jQepES/UbMFpzD0hhFAed2pPAyzU2jsZs/H/W6sLk/gnWZCeItG6rjzEG+G
IE49D07W1eUzCWicgDw/GDx5FzbuE8lVBpOUBoh/AdIqfjd2efhXRJaC34FtrdigdWrSKAKlzYUl
ju43kU4758I5sZbc+MfRcrVpETg2729aiG6fTbCjYjLyuNNQEUgzUFoZVpNllgIyQyr2qZWwWRH6
YQwhxt91fybg14CY7zXGpy5WKYMwjL42GHFaSTF8CjROWSQruGsQSYwyNHJm37W/IyO+iIpcXEEz
09h+0JJElApZ5Y7oWiIkYMUH40S7rld0od9418V63gLvAqO/X1vQ+9QAd0ZzJGE9KYs3q7R1x+7O
Hd2fL3NfOLeP+VTqtawda7N02Nn4ACUts2ky/yEh1Pdy/xjjeZeyK+P+TBQjepQ3wxtVLCUu56Lz
l8rVR6WPgSOrryp/JR5vmaA0X4uy7ZOu4PugavYsbgQ1cgIu9u3GN5wuX3jgX+INUewRaCz0UJUs
MJo/P+MkRqUryDGiMtBLi4E8o4M72Jf5GKo2PzO4ytbVUE6Z7T37Xz8K5qWpUkUbY4jW0gfB4mkj
COH8jLwUugfQeiW44YKMXp5fHCsAUdTeXBTNDKqBkmb5S/ub0zvXZygLP+ufylWcskS4rVSYsDN2
+EhRdbiGjrn4cSGcjdGRZfMWwNeHwqVjKtgGJmA0fAnoKZ0Hp6fuuf0d44x62zXo+s+sqVBnW4K9
Qa5BcfDMxvWFEMTnDYmqAyKfiZlVxMyhQxsjWaift6h+mEBYHt3bgedoKrlYx90mJfsrO+6QgYYA
J5TSbv5PRUWY3tA3tacOcdcaP6/kWTA4QSVp8tjmgKSDot/UmqpmAT12uvhvmr3JLNPg/ftK/qyE
wBOQO8PL4zu+wvXFh5CAQBse4vL9oe/IbTmRNcBGgz4dxiBmQQHkKjrS+y/2Ayps38QzrsLQtUFu
YUzmZQ0t792Jr4iVrsRmFhzcpXEj4051O+7H40eBa0sk6qofO9qEfq8fZ1jVndo6Ag76WJ6i+4rb
QdxbIXRO3MJimz5jExp7I5gZIQck0KaswXR92lySKqw7MpuAtZwaGs44N1G0k4bSD8C+jzHJC+DE
eRPd7uA24qosGtjIBEeWIKmB9rH4KgucEBrg60NDPKlUhY9+4gdeZzFxCCwImqB6kDRLdgcx3yZu
wPENg0i5PjtSQsper+vOBuno0SvTzpg68pPdnMHcKOC3D4KMWZleSqGV3zfWgocY59z9PqqDZOFM
adaVBHF+lBjA6e8pGEq0cLq0H4DG9jj0B+x9wOr/3NmwIXEqm/YVZr7PAwD5cmSAYUyIMSzOmb0P
JeT4hYl49zaCp57EHgsCF2CYlgYOV6dG14M0gK3hb/wEDa973/6oStZvurFHCANOMa56zvUAny0y
GreVzsdegW/utADoB1f5nuS6ygh+xMEWsAQXhmNwo2nRo2AVbJAcrvCjZI77jC59Kp+ywXiYbdWc
MNBFZy8wx1bDaYKauAMow2A+oo6L1iCykzF+3+faJUkOhVNYndPMXbTH206kU42XbKI4qyLbYQ5r
3qbEJ/5rqLUo2oaCmpLM36ZCLsiL+7bORykvA8tyr4DV4xg0EEcGKhyOXm5IOokuiUApgb3asiaK
Ls2cyKOv/dH98l1fQ16dGZsEkNxLSCHs3W5xSe9wZ+Z7yFN5PCM7eTompQJUDBfHYEov6ARNEKG3
fgqc3t3trFKpRX25KiGUWYXAvpf5SiaXxM5je6TG3hcS9F10yhVsYKGG+LsAk1vzAaTc73KZo8WD
sOAeO34XulJBieSQNPIifF4zWc39O0onNwM/v/5AYP2VCqnVOETXRqtizjzeI8CEc4+0TEdTnl5b
WeTtLEdeukkresuCJvPKVEN9qxQ9cU7j/Z/T01tPg11NzfwRmYejNtZaUeb/W4le7Alb6ZDGk4Dc
MGa04h3t6ShRDPgSOJQtrO4jKw1nF+/WrMKSt30+7+9Eue5jpL/a+OmXxyNOEBmMl32DgH9kYmR2
1NgTwU16e9aQQDwkRjTT82g7lMQ/cryEG/0zfZSspZmgI/jpKjmITLJH+DdTPAiO+wdRg3wp/g+P
tcWThBO+FBNP10UYyPCRrbKD13dUwVsuxLb3rm6gNsM/eqKMS2IUXeeNaDpDEDX3zYd486duvdPZ
pFdX72dS0n1VzW/EuGw08jg2cj2xRzZPYBOlyHOTpZZKOQ09EYCZMhcC3I5J4K7uBUGzRQGMfrn2
C53mDMOgalIRVZocbtryiE6r05jwGIssN5re2T5RsIwDfzO6+MvBQqijpautMxgg8aQUZc3/eYiq
MuiMt98Gi9MoUKzl+tcWsALRvsUO8rRE3kNNQVzEcncmUpHR8Q7r9EV7UYDjhVuDNOkZwPdqCuV6
7w4+Y5tKRpQghVbf0gD9gH/+XcNHAyiBdN9VvOx/jH5fy1gYVCGhJ5MOZHuG51dDBkFO+x0gWq4T
bmh89h3d32WE27bRcake6Xad0Kch2NuPSxHEz02F6wuSkEiTUqFzlWhfkDlo+ZQokFB5EJbDCUfu
P9TWT2uMMHzDe8gLxOVJz/OUbln/VVSSQcbPR/n7WcZJuQ7lWlY8/GHmMrQhwcm7FJQZj8+G74Hn
lhc1IpXh/gigBP2D3Ks03OBVO83O2QJyVZUqwfxP9+AmqK7KWUpZCadT086hVwa2KfsAHSlEdb/P
Yy2yh/gLH7opA1yhJk51N2UasxYoxbo2TeCLIrSyqeXQ+PKD6FSJ//rGBBM3LjgQIkxx8Y6j1SAd
XBgVljs24vxeCyzteDomfBMwqwFMIzv8GmlEj+o8JKvKqcGX8+ucKRb+jzaeXwOH2GHkQccAkymN
poOPz+Xgj+1zyp9dkJ+g4Iyl73j4+NGtmH6wbOtWdv+Zf2/z11HwjxQWx6Rvj82F3vFLB29YO6Co
8jcOoFV1Fl2eAgJXtLfHrjZM6pYhUwIBU0X3QaZy6cJuzdD/Pj+Bi/qF/XBEMG+u0FtZolhmsCjr
YDwyqlNUV9CUT7F0cTxAkjIF7RSv00Xl/53pj7C1LVJHQ1iPDJ7X5XGWQfcTxL2LDirVd5zA8MpF
ds77hryNn4Qcp6MHk7e8xg9k6epwojAbbCFllR6YASIIXeAfiwtsW14JFcwVe2l2i9/OX4Ylb3z4
ut5Boh+t+L8NypZcEMmf+Sqq3Y7R0VyEiXXrIzAmDoHaUWFTFy1k42VG3UuF2lD4RDrkLOGcktr1
V5HtmkcxH+I78HvoB3RKNdHwp1NontweXpu8Vf5sXBuJAgZZBRqF0nUlWiR6ohfZcuC3mpoyhjCi
/BezF9GEWjWp5sNJR/U7GXq45BCUb6bUgGIDCxGEnMNMJJrvNerScrrSojylrKNFSUiueQDxXDhx
5O/Sk5pAo4uU+21xSLKsp4Yi+aK/oXgB4LE840Uz8L6Z/t1QCOSgtqftXNjbglCEL3uvDfxjJCDO
3j83jE9zZXeKmpYQ5hbezHF0Q70BzFRJ1L3xWTngX4PR4ouFwyPS52BStOJTWRbkdqVpS3MSCCZ+
5yv+74BDW6AoIcqIfBPAqkmx2vMJ2WZjbhL7ZLSkWzUl60+PVvt/UxibkKrfSF+93jlOegHahm1+
lPh8OcQUT8K+UGwYL62W2xNfA8a+EcRwYlfPgI0IloV4aoRAB6Q2wdctUPA0isdCcHYEu9bcp7Iu
oSngaZwc1SOvkofEHrSk1Vk8EaSrSCMtT7byjYMzxdtoZdWqfsN7qxZVvlh0/7DQTntpffXH6hMY
d5IGKEu3KYj+wWcvfE4VZ2JGku1jW9gtfPujGt0aScas3onDzZc/7xKV+nokggAsrc/0PRZEVvRt
elehLcOvW6Gqx8KVCR6ODXB2wUUMrFoFmmXj7MTPpfhl4qHyTP/AlX6B71WV0JuFWZ+iPZ3l2i9O
RC6AEqrdVtRr240V7Hv5o/poYl3xq8uobfMoTIeUOpMOVCVLufpKZPIBlmCbThBlYawW4EXjfLJi
XKmN5ucw33NuCuuPHZLuw47GJZSNFUeh4uMiHsqMTreTv1K1nv7D9x7TSVcKlitM85Sws9XzB72L
whz3hiKiWMQEN9jqpdnDY55QqNPK9tBuEFEAf1SP7u29JBov4hk47uz/lBmOom02fFPFQSTW6XBw
407OxUEMed5SJRElmnR0ho2xUyuPj+bS1cVQGfVrqLtCkHwu3aKQ4A5py5s3K22/7ZVpNYygJoeH
3UckIjiRjFRuan6PW1r9/vWERuRHWILFcLUEyr6Vle6bnJe9G5XFnMmHjLVNz7dCPisdZFquHJVA
NrzHMyvCxmSIXS3u1pzesjeHpAcz+Dj7Vji52e3oQHhY46/yez9goMTs8rvbt/hfp6r84wE1hQ3N
hfVj3S9wwNbveSvnR0IyHr8QTAI/g7GAus1zFiDb9mcX6+aCcoRhhKh5qQRjHdpZDPv0+hng37KV
dxsQyDQD91KxLuSJMTqfiVaQ2NUIunnZNjiqgyT0+Um2cohru/MvlF9wbGU1fQnxZ9favUZGtdGO
J7Uco5993qdCbN/8noOteOtKxOS1NK7LFt0EEJooP31Wum+7X7jcKGasDT/Qr5xlEkzZSqNytVCV
8UXp3pxvbokhurX4xXgAmiRRDPLY/Nk+/XyPOltbmi3ey9bt13IoWpGz+tsFPpqo5XR3RRnxdqn5
oGFoHVam3Un2DJHyNgGa7kWVf60np+8IKXX6Or8QxTaGQZf6tqkU2hOZDMv0T6N7lslPJxFDpyoq
nssf8gZb+TrU4Oq/hPQ8Ra9qd6urN062cQo/EpYL7/cNXAL8lHesAjrJwiDpSGJGBqwZYES6Soxe
glD7UImJn7sIKHcyPPpH2a09NWZj/kUcsjO9gxLzLxLIZ8AFTjEhADqFDrGOUY6/f9F0bMxxBCzg
eHYziwJmR3MOFzBmaPa8dURajU/od+ZFsOTrvjVOIKb43lvcQ+F7tsuUHPhhHWt/Cru1zwyM7pM0
coLMxmzZCkdwKPfk3rVBHxG9xkUImbHKwjatvv/WapK3KJFXHL98XKIhol9KjNDUzTc7JMyS3u/g
ZUvtJXG/H8/AhM2IT9CauFH5byXYNzHoaxPp4OZBND01uYHe+BGKmisyn/hA8TUbMe1Mp6Jb/Xy1
sI8ArGhB2Wf8iWxj+sUi59jw89CWw0ICCPcFbCtGfe0lkjqaOdXViXcfZTwBVk0zYfdLB5Pkb8SC
bdjKs+su3lb/AUO1YKC5AJUwU6zLXjG0nOLSTNJXDncVd+zYWVGrNm7oar9/Mr+EGIrviPCsWHV4
AjYTTnpior18UG8CdMNvXtxAKztvyCfSrWGFMJphV8XqcdeldP8r8pYf9KeJyP+bC00yDZXzh+VF
Q0rScs9WQYdI4BsToaznAxs+n/hoN1PHr6EQ9iDHA1VghTYFkVXL9PjMIduCX0CpAZrXSJYJkE8I
KhvoWidNbZQwdAT0Vw45WV2w/i0MdV/BqZCPaHHaxn8v3V5y+K+7cjEiX/kJLO+4t2Oihgf6+dph
wUGi0w121DA8VZuofD5XTMfe/FHsoiGbA8+hEwe5vFzmxTQp7OGEaSNCGpSFUNKKaubc3IfNZr61
c3+5LpWvMDaqDKXHVEWZj3UZj0/IlrTc27qN8DHbMrOo2q7524wbJtUYhhE1JB6Xi6M/g5tQvNob
InNPABwdbxPb1827mcrR9OA60zkAiwBqaFK4wHVi3PGQuyyd9AFtTM42WEbX7CmpT+ZH9ngs2Cip
gzxrv2xnxYjbnBqRs7qIi0mfeicaVUkn8i2VblUArXR7b8FjIbOg0FvdwuCWB87/X2vxzv8s7Wx4
aJ/3/fsuUc9g9VeSqMjPC0qe2B2h6uBWyGdA01Fi7S+b+h4iNdGV2gUgW4XmzFU6VeRKrjdCVqng
o8iwYBMoso/+WUM6v05TGfvxlq6oanLVmZCyvRsKpDogkm8dqvY20ujrWEwHue7z4fMU28waHBo4
mhLq35MXO/6G1TonZZ/tAha7lfzB4zCJs2Oe/iwTINZy24iG/F+M1hWVD3Gjto6h+tWLJIx2l6Jo
qI8N0VMTgHDh+4BChiZ897NyDuyDq9rQBsr845Cyswi6lmMadi7XAxJen42kLb+ZWDJAI9AZnPKE
3hpL0kwIE260CU4pnM+2KYTZpFamRivPCN+2sPMQVL9faz4w3h+ftcDhwsGXCD/TIf24pDGkrpFC
A8pwZxYIpVvET0xL6stX3zXSZqqzXtQ353efdhyNwxWZjTiN9OnCfEFdJ9rRCi2ai7lWO8EEfnaS
ixJB/fu1nwj+goFg2iYtrPlIQSFrV3Gua0znLIKW2c/ud2iCIjISgut83VwXexT+eBe4TEt/Ro64
RK5YsrBvZtX7Ijc3tHUTm4JKAV7CenphdpUJcNdz+Rb6Xz7gW4Q7VMxcy6fcPbJR8ZhliEYMiu+m
EuiaU5lNl7KLJBIUJe87/oDgDAVxUHNKxSVNZno+ZQdIdPX/QlATC0Y+W7b2NIr+SupvTnh25UTY
vZeJgj7MSDFMSH53k5/s1d3p2eF2vhAuL+wMR73KTuVvF4EMDgSsHJ0LzZDftpNauJBzk1NtZEaH
zbK85BjyfrCjLKj+rqwki/AAV9SZSSgd/YzPHvNwYhmnpuHCCZ3AZFX3vi+EtxJQ5OBHD8rDDsQF
jCvk36lCV+U955phqiH1NBJh+jL/VFayWYS0IZ0fKEY1P38UwpD6ijpMPig/5y2YM9TAljh4tbG6
Wz8f39bgBRlDa2KXv6xCac+xJ1rE7lKxON1zOja57l4Gvf6YmU58RSK6i/o0qEfCgF+XTlwKHUZQ
yxa4nUdJnSqgSd0MvMu8fn0yBbooMcjm8K+J+ZP/oKzcgd2j5cEWy6lzC/18JiLWYLwag8e5ezAF
j+KtpZtbFQJAz5Tsc8Y81Ef5Xqnw/LGyUw3HzIeN0+d2PmD/KIhBPTRGGjpgMnEVPEB8hdvid9Qb
/WtxN3ZCu9XAkqN5PK9bsnrpzvUedS+yBRySWaj5qMO4fCHfdp5/LntzFl3nyIONTgNVA9Bz1RCb
OJPn1S0F1UnN3fzofwVYwEBNaafpfUbaDyBqqx5z+/u/yzczcscm/jTg9MHBFgpyynldIyRQ8k89
zz4bOyhQEv2NgnoctPwdmUuyDroshTtkWVuKDN6t+A20tMUUPGXaiL0FsjSXA9uDTVnhliD6lPAE
pQlkvdaN40byIIIcWKTiIBXsIjlYvb2jRRwK2npiZp5zJyePQSlDv5ch7bTC35RI/aFzMj/vA87C
SKzMMqqLQ1K7mUHwZPD5OJI2SvaM31y+X4sitc8P07k15dr/xYDvqQonFAaTkfbOPNqpgqvx3A4Y
t+65NhD5ujTbiI/4O3TCZG0CiDroyVYFPdqrqFCzLJq6ikObdStdMj1w+nsmS3qXeZ4oIbQpzo+0
X5byiG+6HxqZKJeiz2jFebejjedVUBBc2JPTrCqGrzuAjudKmrwToKTdS1+1hoSqwaaPM9uFyovg
wOEGFXOuRZQotLsBy/dNJiKXWNNMyBXqpG0Gewx2Cf3DXKAiOB58wD0spVBi6wcgyhLrMtcnLHIS
eV+pH/gtqnyNbxbqG2P9fLHkh9hA9XDtGle/MFPulZ8QrPDwoRR2GOYLqp6agzi4Z3Gln6FuJVIz
a+fwLfUJyPZuk2ffPXtIBANWEEz5AbeiVIC1wI8D/TEQLiQZaHo0XYxksJ7N55jBPpTnDCSVSiNC
gFm43iW7tPpWVRxEGStUzuaiD7nJEY3GcCSsjThVvrBmTDq9EP5h17RWYtPLFz9tqaih2i1A1rOe
PqzBXNC7kDsd94ijilk7pksTmK5qj6hsqdX5l2TiyDAhIlSAjjcXiGVUnp6SqKaDQ8gj0ITWeYhE
0vfG7E0EgtxOxGkiVR2XnUkRg1nttOaoMfJp4bPpCrIGly472Bzl01H21WFGp6WgX1z3jt2Obu3i
gCWzi2CunrUxxl1apHtiyvakzFzL+eWcK37P55v8NRz+PvFrQQ6a1+vFXxyInO8YFyeQGRMb233A
ChM/SSR7dsQ3DeVpm0SnNXuGq631qvJRVpxoVCKuAKwA+yQxzrKVB0Dea9HPyJWI/kk4Bjtx0Lw2
vfSFBzRi6mCzicJ/lZDcPIDMswLJ1zwR+9Ju7slzA0x7T/b3zwQrsCtABwcnYfhzQtsLiuqGjEbB
lLtrNGWJxorS37y8rPYBClmGhFwSKVpcGVCXfLDAImzdzYn+nba6KGJXbmjQv8xyZ3Iqrh01tKzO
IsaGTt1I35OXAH+9QfT8u2NXMXXdHR2w4h3BDRyxfdPJUh9cUslGqk5Z5JgEu8P6Vs3yPxTCUae2
sugpZVTLBt43Jr4Aw7D44yLaQPjjynTwCdMsen76S0XqT5YM9L7haaEQrF+Eu8sS29AsMooiWArV
ZG75+KUGqFMezSgGowaguZ0qhF57Sok5LReSNJPJ2rdHZF6CTMmpLWsACfwh/JoZmJwDxFU/J7CW
PS1n85THf3N3hjHbV59sg7wrKVTVmEBkRRU8pa3S/Rxvfp64kDMq+tzc3dWx1WfBCg7I9afTly24
9cr1kTbCk/g2EhXUhh3duiGPAL414zKddgTMcOEkcz1KMk5b83lKbm1N//1zZ44js67VYT/s5KpW
qHuq55AeQxDflwjwtMTobgzh/2BUT93Z4SJ5OR59mAwEiGA5VN8T6HU+zvnJUEi0dhbj4Ta2+OsA
8m3u/Vv8MBxrZLKmLW6BHpT4HYcTH/T2D65EPMsu+6VRM2CNpXA91KLi9jBmwmOSrlu6JKnEqYIu
LgYr2efzQGyDJ+48rExdp94X58S4L/PIwq01p+Las+n8GtF83xblGH6wevfViTP8xeAkZIZys38W
zzbH52wYL3WyjQt6Ysg8bWd044njBD3IMbB5iNjkErGi2kKod29M5pqTZPbZV1la6+i+nFx4PbPw
QwGDMkmXQQFLCQum6DQhVj5ldWg8+++9zdN63CQXafejWFv2YEalppohj/5E/9+Cu4hdYTXWy0Z3
g5OOmBbUBHcnFzF63cKpm4fHn2bhvvcCDmo7WrEOo1EBEBtfjljR/bL05hdDmHk6/jCfQSTfFJzX
/a6SZf/oOnX34dWKyHO29DK8+JojGfSElqaf0DuyYQ/9ab/SYhWQJ6ZSWDF7lz0zw5E4/LTY1772
b4wLqpdRDY73yKqo75JCko1bEx8AfnDwYVI8qon7a6jZwTHhfqoppMimMN1+7oUGNtZJxKXvLFSn
aWI5rU2y7bQDjpr2qDHVzrOevBi9qZo5rMM5mD4vfiCGfC5o0gBqdDQquxb5QZ+wnz4mDGJR+nZH
F7CW6oixO8ck/KsM1FTyo6oEZ64tC/BNjoJT6adSbnuS6dVVSmHf/7i150MgDv0V3apcZu9px8iH
kObxpKamWQV9eCH9IOHujIljoXYVZO40I7fpJ3AEdYAhhT1wSZAEMRy0xXNbeJfptAzKnEyYfRRL
KmY4RlXzB0WBezJgDQX79HGhL2yg1IqIilw4ZRRN07s6rOPxSivTvouvxXphRz71yY/ttko6qGMd
XqwMraC62R3QRx31bV69kkKGSybviQRjaaomhwhC1C6+Tm4XZy5SNIns4wPNDR/7FKKFXemCzC1U
QZH88aeMIfWF2IuQiJchaS4jFW1ukATkJq8qDaGgn9iehwSnSZ3sRizdpL7t41VV4cEeplnqFVfh
wiBbX/bYQ6VC3jnooLIx2k5x6RsJP9I/RfJmQN+XknxNr89YNW5yAvIAk+3HySoMkL1Vm6CwG3a5
ppPsMn26nKp/wGwaayFC10sn188CZhXfXRkUWfMNvmyQ0xHhjgVzGhbe3l/u4a4BW+LF0CYAqfeD
59OyWo44bK58K3tyGSHLFsZtp4D9jAK9U4eb+lQ9rq2UtrC83ZUx4so4DhH7JkIOCEX2H0gqIJ4o
HFXyxi0wStPGuIjCzWJc9rqnJcY0adC1k0dnYsnp1yOe+V4Bkn+vF6WvHSa7NdQRd1Zx6oyoX/oq
hxSewzIsrgKV+0D/e02fjnT11zfak4FB7+7Qioh328r4wX8u7AcuC7ZjAodoqtwwK5wNPaQdQnQ4
81oqBX+CITMXQKnUmI770SfdMcINBeqU8w3AZJYcENeTGQVZVSmbaKrwFAYpunaQRMcDPCFe3qBp
pxPVMIQhRcx45v2uLL90da30b2hdGTTsQP+H/qMb3u+FCbPA/5CsfJdxINkCZa/jx13FTsCDKmjb
aN3DImLXE86aiajNzBTspOZ5ZPfDzpYwejDpzIF++iKjVXD9II6zB1cvbnbXuqBc2mV4eLJ2XUkD
qStS9JHPwmjOJG7RLbu0k8NRzjkDbCWFVKjyUtZFh99UEvdz+6K28Hpx9rMMFzuGgh/0LAmLoHrv
DL4eV102z7v9HcUpOA4y+jU6tgSHFhqP8FhoPH316mkT8xcw4QDdRzgY1TFRbt2XI4U0zaab58jU
kPD//+lT3qghyytbP7rearTU7M1p+qg8zE9FOeh/4aIuj95imAksW5S7VWRNRKWRQAMQK2dnACuH
TLELuSLAzsVqEtRFs8DxQvpUF9uoys5WXAeFNxmY2EZjLBZP9tyoRyydQ9mfdklam5kxgJJxg5g8
RI2atELXznpvw/OfnpWdi0l7a8a+RWj1c13EoQZ0Cmyo1Mi8ieLE0CZAgZBqjwl22lReAmZsdxTh
ogSu2cz7BZZtgYILtrIoJIIPAZm/JorZjgCUpOJ/9VNTQnGBVhZ/J+lp1iD/S7qOvBatxabBhFUY
5uGpmrmdGct2/3eQFdY/NXkL2uDKwcgzTw/+KoEeUtRF1B8HnU8JeHLR+SvkWjwHkcbgKbpVBaWn
HQWprG4xG0EkOujF/P69btN3U6wTwGgLbmKQIw7KvrB8CXDrTcqN0JwjSzdFIdFKUSefLEAG7yEI
yZuE4yPY1C+vRU8UI3qO9+RlrF6MldNj6706LvE8wildVJYHnbJ1qmRA3JBD2DXIteb4INr7JPwW
chSF0BbZvBOdmYG5LszC+njzP4enTfxWHhwSjK5kTvv+n+g5wJiUXVuZ6haL5V+aG0yiGbRyEeTT
FDuG0uTyn1k2JHr77yba7bdqfrq8nrh/usKmUFmromnuMdLxjmx5/bz0cUG7jt+ucFwqjK30e+AH
HPYbHLAL+TuXGkVg1zi+Owgdi18LZnerFEwbTg3qU8TzW3bci/+aQOmIN+mSknuvkunBejfpc4CV
HZnH1G1u46/WJJl4RkDYMDs2W22SolgPQnbecACtcKUEu2pEdHnQTA0hA1QSHrYpP7ZGGjcgpIku
F7am/YQpWfjCJM8XxEQ7lR1Pur9dGL/I0FZMMHE0Mqak/0qDjfJ76QCnprS27SoBRatFdpuT2noy
z6mT5KajVFJ4b84WH6vQP0rmfKhEvDWtQog1uBr0iOrZmWWKFYRGO8pvJOTJZz6OZdQlIq022grY
agTLT1UT0cWZzQ3MSvXc/wtW195rh8i1TS16BQQbqkETXrIW943C0YRe6vLmelru2kMTfvT5l7uq
izglG/wHrs50JRHowPMpQd44alS6Q/kJH4KL+RENT7fRadnzkAVs9tlgm0nfEw8oezpTdvV6wZXX
eVXkiiF4AyhJjNNI8e6HtHaWtTGjM4YdKtmpy9S8Qv/KrdThAv0ecYqp2uiaNo55wEj2i9butk/1
a1CtQS0a3Ugeb8CeM/Q04EFC33NO48jp3BW6zOJIMMcQIcbHZuMdNBbFpNKIKfoQaANrzbwnP78b
6bgEo+YeOj0NfDzcteKhGYS56R8kZIbSCCS9mQcExiKMRo9wh58zs2/XUonZKxaQ5oWZxd6aOsSF
zj36SQnAEdwmdtB7Jl1IbLzG3YAHwGJDfVUTGpLlZ67i+x/+A+7qIGBJMydE8OPW7dwaMEdLQfuH
tg2bPNjeHGT1QVWDXe6g+mB7mJv6ZUYoG1oILtN8cuq3VrCBMc5Xic58k0vLzgaMZ2WrBe49jq4Y
Tjh7CKofTthb76rt4rHLIMGAtUIKhHyvApWwEajxvNTP7dJO9/ebHOOmJxctZ2+i1NH3urb67z+H
64wO7oBrjtonCQuSgK9ZLMG8spzPGeL7Lyhu8CmCHsj0bxVNKPiaS4ifI3GCnjVeTgxHu4hceiR4
LHkha9T3sEHkux0YR4QK8xUhp48GFZA04JZLmcamwLlNqKKvL7UPtiz51nCvtGU46+O/CEb84azX
kgMxmYtM1L8sC/4Eu0nn2mk7plmBMzNmvV8cffODJ5vYaHiTbQC05YJVVrNg7d3nr56Fofatmq4r
6+JMQNpqNRJIOd7WcSNTFbkWZsT8uMAj/ylxppshmIBrdVahtwvuHw9tYywUZ0Stc9K6JaWCSNuG
+77qjlzJK09q0ANZ3rHPADnbSxoBsx1PhxMSKLuXJnoOqoSOQ/n5tQkEXGdah6TxZ8Be27Y5P5eD
8fE4hhUlOh8tAIxiK4yiP3cU5gbnz8ZMAFn07oJQqFzVE+ZFe+bwPXwvsDLfh+rFQsXeh9FNx952
WpN2W+UsWAihXv2iMXzd8Y/WpqCtolOXL2GgYgADslFxZjstpMiSiHf0uxb5TfOHggz1EOOCJEya
YYd90GMNg2ctXtDEHt29vTzyosrRLRb35V3trbRMIAjJxUDVeHIrQallztzM5nfjmSju5VPacBqD
xoF0p8yowJEo9RxWCmuQgX3nEikGuV755j1DbXdpV6Wk3BdU8TaehZv7evVqY13KLQghYhvGBgsa
5H7TijgzoaaUKQwJAGr6vdU509YAF45uYBfQNTyMhUEcYOaKyCufPkgJ3rMA4zZMryaN2nS/WIeV
I2OUHvaAsk8LAKFXPWAFLBU1xpKq+2uFzDPTtSTUov+H8Qu01yGJxjxXTVlTqxaD9QI0PpReAQcW
FiO+EVhi7DyDHsNOH6f7HbWww1r1SnwJpxWC/oS+T2YfBBjsV4UIw0DH1uUP17TPFV0z1UYKwJzF
+vdWVNVs9ArTkMnCHBs39kW6wfG7T3GufxZkLjj++hbhtDFkgyjgqOQ+l43HM5ftdU8Bupb6A6TY
m9XM7ahE9KA6edgQ8WmTK5JKPpxDe7h4NmdjIDxQ016Ok2MXzIdqovKhg3q0BLjq4rVV8mz7xxJa
bKXV/VsljyAGBAyLiudDF20M+bccjdYaANbPRVAT4Vze71MATXAMHhH2jGjrAQ498S2Akp2rJYer
lURgIk3DFT1gBAioio3g/zyFaXZp9SYM0K/egZ914u0aywxCyXlTcnrKCYAWzwJTYwwyDcvc+HhP
qBYExnFfVZ8aZld0yhsVgWdHWD4ORCy5l4icxnzaLjdWWRXpC94hpCmzKr9sytfbfcWpZfEb6DQZ
45L5XWN+6MNX5JcQdDR1x3HAeG80z84mOSQLHxsGpSrP2CGSfMzOQI047Xmu9g2T8e8s5X62MBBH
8V8hvTzONCP0r+ulcZ+39dJuOUqFiJ0/hQRT1R7pIkNRT3n+FwTWJoW/aUmNE/L2mI4YMeJUPb/x
2GRrYlx3gYsjzpkXVT21vGGcpKKfp88kbZJfgjM7V2AxQJe6Av+4jWXeCD1qTJtcHmu/SjP5UrV+
e4N22X2WQAs9ijB845CUNy0j+ppqcHpx4yh3PLL4iYoL4m+DkEIuGm0Coh9j0LkbSPY1DV2H5Kft
3RD4l107Rgn7wac7Sit6zu/uepGg3jyo/PYF8kfL1Z/y27TP7V3jnV0fjuGqtddJY2Cv3zTlhDjG
P5raKR1G29f70zFKG+8wrenWeIq7qMK1WEQn5hwG3W724gPZsC+bKAe2+cqDy45RIz5gdzvt/YCr
XAUjxxp5uYm5CJ1IYxm++rdACL/bcgZ8Yp1U/XuN3VCfhnVFVTKcz7yglOF7cdUKLL8e98jYTc2U
NeiOetIxtN+ujdeYUCXf8fwjU1Nfkl6g8lCntsvNWDrdd9w45DeoQ1b2GEzAgkmSpNwpuClNaxyC
ACblZIz/z0/UVsXbDXsd3o3uHmh28uzrdjOZmT/OECnELzUeWqikyoorkTjrBm2wWV4YXkSX8WLp
BduzKISpCs6CV21tKuaMRib6O0btKzSMUl7VL6KBObKptAFD9M8PVy8tAMrWp7d+4NCjGMycrHNE
sphw3iVoC0DzJDMH2qDRgBuEVXCJwUNhgn3lqixiWmuuWpUGW0ZoOkKP6Wts9kNhExqd22h1h4Td
qB7AGUQabTUmoGUAO3YH9d48eajqi9LgJcQ0QBtomTe8KPJO6L39vByLZ0goYH5apF/MTABJknQk
5IJdM3JmFbKHq5wX1RqUq1M19WXjx0pADmcQVoVLG4Zt++xxN0rt+9ysKM/uvEtzql3qkasuhZ2X
6pNdh+KD2TYve5ywFDgq1W8k9DoiXtlXUlHwXk2260ks4FUO3Ugme3+5HpF1XOxm6gWSZjE4Mpe5
JnIOndoYRRZ3n5j3Ljj/fk2Qv41CFb4NSIQCDJJ1YUD4e0AkiPY+tXh6Jn4X95npRMsonVv8tfSb
KrABv45eMVUgcb8JNkXLkyR+UMUeKwZ2rWNxJOmCdYkBFzFYK/YKsbl8UXDMamHvRylBTGrmu8vI
cqTRQeQ1RQZbQQ2Vh0Px2tJBrBkwioRufCa5ytdOa9Gs6kcAb6Pd5x2/70tft8GAWLSfcV9naQ0/
MHgVqnS5Nm3+ooKP/uzt3Jq5UqF2pc6OdV37CW0q9xXyBCPS5OokMAqscBBjgO75SwHDkmLFnAXd
c4euGZjdv25lNHLkmxEe/+xSBrMMR8pjuA3onCKXx8mY76vH7ZL0MLHcrvPsqZb91ahzub0TKOUm
M0lK1931AXsgQYD8ZHy/0J2t67Ti8hBy/B9fI5o4yF1Er8yoVdkdEVG+43rfb7JXjIBSCph4GmmH
LBdLSkMlv8ixw/NldJ/xiblrq8jBHNnALPTH4KHY4TVlh+sbBNUwzYfCkF3vZNbKj9wwqugkOwTr
eskD6O0Sg/3nYDtcmDtRsOxHGc6N+n4o4Opu1yF1nI9vF424jL/z8J83zHzhD6wJZS2wq2iYjAR5
/TSS3Ft0JeFVbzcPiaZw41ZCk6UaqcR7oO67P1+8cIpKvYQ2udt/dNkNEEaC/p2fBKv3H8vkWfte
R5zCYCWSXlzD39+w7HlxHe6/mvSxTqlT4PXrmBGGoEmxyA9+13p6R6U6t8WEK459yPOhFTbSy0TS
/VPzD2AKCoHj5/ojpx6g4K3xzjq3Xculc30ZTRA6UELVNGopaY2x9zMnBcYiCg0rLaHWhotG73CA
kLs0rU1Gu1lE2mBj86Z76YaHIXf3tLlx58uw/c0sQ1+wSkfGtzEW+DoYKlQfzkMugx63zhySu2JK
yVSMXpMIfoVLwx6ZiOshemDQkZ5pftMO3omtEBtrOzLOWJqnYGHX9cpm/JEvyEJl98wNKoEk6J4q
PbmNk2qBPULK+cQImiA4Msrlh46ki7XLINArbGSX9PgY7DO8/tLEKna1qvNIcAv2Oncw9qhq1nrp
JmeSUxbokXnWg+pvHCnKkveSFpvUEzkiKVKsqmYu+0ZFVNyu381yXmAyeXJcSkpAhcQx5S+phyI5
NnCKTnoJNplzaXitEXa5NlEiNGz08/iLORSYZBgxUH0EB1nWuAxfnMJnTNw4FHB9Q5OFO6ipzD1s
4E75lRP/t1FMbeCydFkLx7GvfwAhFzBwWohFeSEjbYb910gKXeH0GbMZOAMbb/uwqY5J2YQpFLL4
q9hjwvTHMTn58MUoe4WnDg/f+/znimrkXQOhl4y5SNNDfpdqgZu9pK07K3XQ0z7RKHs0keMrjdUF
6gZsKD0KdeZ3SQIZbwIfwtn3KvorRezgBZUOxRzaIZKptJnaTCDJhE1qJg+nzEDH4sTd1cPiTzUh
OVk/OjZXaios2t3A2voV+0Egyj0OZ1+5wickSD2fZrJsQBZBtNwe1uCY8mPr8e6Bh+1oB5CvGlWQ
dAyPA/q++Va8CZa+0zkN29xBV7H5ZNd705LJklsRJGLPBlk7eXJOGKWtp6KNaTLWqO+lIwMMvHYL
iTpY5nCFLD3zjdRC5lnkI/DmuPWSbO62raQD23v+NRxnzUQq4UBO94Qh7OnMG3Ki9+ckCvlOs6yX
cQ4Pt7wenA2i39oqQJiFA3fVotUY+JScAzb2Wiuy7WJeBO2M5Oa0bL6Nx26LwXMzVBmaJzrKZ2hl
Wx6+naWYJeuaSQ6XBTA3i7/eJ3BQ2IoVPbwrVrcz2S82abSgQX1pS+ynp53NRDii/QR25WPXAMYM
XTWDwIsYTrop4O4+QoR0nCjm718xNrMkC99v4tXB3VYdNkg4tXFcCFtZLdX4LQR6i4zBwdS2IQHA
0sf00+1GTBaGdUXWHGds6ePkxeVLOxA8L9Gdyr5XaabVAgW5Uwi7lfxl412+RmqU9t4yT4Zvl88T
4C3T4OI6m3wuq3MdtDuw9UxHqbfZZblHiDK1iCOKvuUy9y8Bhajzot8C1ZQRh1iz1mXMR6xcocaz
wE/sIbO76cVXO1NteQT8UPHDxoJDUDClnEwOuA8EoFKPfIHT1KuyisrhLp02Emj040w1Ba3hBCJI
gbdiW5Gyaz06q03eO+UYiHJHC/107ugckoEGtCyEjVYuSEWSO/7l1XGKB0TGCNZJXeVZVJPlkm2e
pCPUHuRKz0EnF+1TNTydqW8ubxVZKPSM3s7Wgf66DMbFtonfuCCGuSuw98+MoEfHtP6TMIe+JBjR
2PpjpedU1O3l3+joJyoTPrOzAbPlFRehWvC/9foryjQGKj/oB+KU/tWWljQ2BjWcSo97ffzx6iPr
Lsy6cBE+M5At9WdEy0Ejs4DMPMC5ToBWAxvRO3F+K3OoMGOkT+4Vl8zfJtzr1YuqQQ7aVaEXb2nl
M1wetmKvY74rm+EQEajlgjzIjdWjXwvhuKvhdfThxC7S+/pTLPNTNhF2vXt+O6+VqI0mAgaA8yKB
gEAS4zg9Ufe10N5quckcYe3vJS1KDoqU9D6tRQl/nU46STeWzu8pQ5ybaJHehga3lOphJWcLT4/j
xXzQBwo+0EtmnjfRzb+p/3oG8S378PuRl/hDe+OPx6BOT5VAxEsUA1KM3Ur4OJl+ZMKWhnKZ+ocO
6Y1DGQjeYTsm0104yJgKzl2eY1cWWfYOA6ZxXFEBbdV03G85YVNMzdwJwTwy9eJLJMIV/8TQtujD
X/hy4/OXYSqAauBKjMTH3eoH9urEkG1SQarDjcEGJvkGEJkziIQ2/BI7/6W4yP+kv5jvri1pnhhd
w7cnHDqf7wS0jtTBWD5XEfeIzypJU0fJAjElks7HabGgzXmqL6fUTjuulWeVSV5Xew7B3BNIAC+D
q/gqCMPg4cWpNR47O8PGLW4wzh+o54+3TqseYpjsefN+I2yaoIYMQhNdZMQcpiRGl+BxFVqAD+Fw
aj+dpbDziATGeUq+1fdwojVwjqTKWVzuK0uIeFLjiPUn5V3KZSbb8P5YHCeW/ZQNdWVI+JAcdTZz
VrMGit4pOjQnQbiOPT7LqIt+nj8fYCu8yu1snezHxsYOgO7wfgRqmBLAROo5mtF41NKt3wLoHoqQ
qCi0IcPMmCmf0bHihK46rbn43NZXGQPEAnzHFu3xVCKh09PX9I6PFbSGqara9kMzY94yV1pttMYd
izG9egVRYmaMR0li59w0+ifYH/FgLRmw/BNWXqDbmp+TLXF2SkH7glCkCgHA4lco6QaEy6gA/kA8
gNtg4VhOQlnqvPdAKs3tIX3DU9/o0PdIpAfTegtWj0aqKzyprrrvHvDIRwCyZkCIGeqjXsTCQyVv
yU93ESrAHa8s5ZDuAjqPSmabR9bdJOIH1ixFr8b7N7mftg2lWenq0eHN2HViyCjJHgG1YILzLBi8
7K+DAEDUwc4Yt9+GTgatWfQmp2S+338oVV1Nfe6UlRB8F26HdC2V59Sx81tlr+zkkWscpCea0s1b
lIpJNZBMKI1JI8WQKeFndMXnDAhgakwvf6mZFGjBsf90rObbs6rtKqdocc571sHv8HZUKJMPtc/v
TNKyP4YdQ+01iix+9UNYRIeJODTP9LnZHfgXGdqNrBIcByC4FwuHDunQXT8qInI1k+P50oP88Rr+
G1gS0gbIvrN5Z+FKFLnn3clh/hCVE2CFPjyPjIkLSrYDGELQn6+tzWoKJNQMmZiyUmjFNOFnK7oE
Dr2FCZSNaCAY3/Or1wZDEnXHkzqgK+lqtG1RpImoH+m85EyanetX6YTHNRT0yIdGxS7XjtzoG42k
VPhbQRF3aKkc+1axU7CZaEVsaDw9zQPec96YV9bdv18RF23ENLayykIHR0bEVl0skxlzsFmZvVDB
dKPB3XwB1eZfyE81HyvsuYIf0ndd+5b/6de77w18+0cruYGuQk5cy4SEy75ehOjLtb0b7sQSoZ3E
1BT8OboIEWJ44SppWJzAWf1bZKxBUstRdlvbDGxha3YuXwfCcwYmWS2PISDMq08saFar3YhIhI4v
RxMuDH5ap6OSBWIXmTRsMfXmqcxEELWWrLJPRtJneaaWPL5gyRNIuD+SDFuQbve/LJ1YXmSbMJ6F
RfHcmNxAfwi5mWtU280FGKIM8d3odGHXq54I1axTC4M/l7CMUFWltAeArpaQsQKk2jNhBJsUBGyY
/Ar47NSP8kEWvuoUhWFZ/HN5OP/RHmQe10np8UYYPraPhn96Xs68/CZvoYhtPoAw0L+IuH45SqlG
uOeI6hfwkpPCuGGCrzFA4JCtEX77KnEhkp6UalojiA97iuKjRcOrHoNGtgbFRfSarHTgBCqq49l2
aJAtNwj4PvXYgSXc3GruWuKRwyg2KAe/W346dxCsuNdaMs7DgWmP7vwCwYAJXZTn2IjYB3Y0uWmm
WKVvq2sXEO2xBF1Ox2erCc/vS8jkvBO6eNNsqLqMvStHOsuObt0bwFJqN0AIjQRnBECGVfmGSPmu
hOgIQbsXoA19HkopMYDCkdLEYgv4mvbw8AxJRxYinY0vLz8TDyyJ+Gw5TnI1UC0PasghVb30M6+G
0h+mcvZ/KLlJDSu6sUOuMGwdhpUBv6o+dSDvKpS3JTw2wrEBmJPFKeOGvUqcbv8T5vNA14s4HSRx
e8d2KFxUAWURHdSUcUA/fbMZq72okp1oWmp6Zvd8tDwimIOCs61RM2PjpgrQjpj7tDG/EaEveJFK
fa/2ziZ16zOK7t3sey9UR+aVoRXWAwXGTg3h0lhzlO0LnTfppN/UodYjCjPwA77RxLLRLTLIdfYr
FF0SI6RmcSAkTNK2JKaDAwwxjQzQmur7le4iecC3payppUVPDEOaxAa+c1BXxZFPxOvmQjytBDJt
IlLubcZdUJLadIbtQK0pwW+/lgoW2W6bhVO9OuIHiNz36o9GEHADe5w4F4G/L56QDLsfprtj6jb+
Bg0ZYLp556GEhFvL4yz8NXwQRTDBpVyAnXkKVHQ6aA5Vym5HT/qdjx4c5F/1057UZvZ1B/0GYxYd
qCzQq9bAndMxYrFVxftDjlH6iMBOteyTc/yUQmIi+/ybJ79XqwuySn59DTPlOMou7XjgQxjX/Zut
4gdgjbtDodjz6j/PPVln6YSn/1B5ueR2V6Yxj1uQ1KNZkBla9K/vfN/tOPGFXen84JCXd59edoco
8Mp0s3Xkchb/hBldZ05ZozYxKoqsWGpyrWEQfmh14rsJM3O10+IG4hA/nc3PYL8IPnOD8sC9NfTY
Hy/d08mkgaJseYMbFaynViYsmsfFNrkMC0n3/T6qqQY5TVCWn42M9JH5Asx43gory1A+/anRDxM4
XhySrIK4qKRtPgC3DMJd9TvCoxLaQMqTchXwB+e+Pss2MtZbbf/V0WnlyFTvzFzJi0H45t8pMpGu
8r7XkkSK9vn5Lw0rXDSgD9HCDm9TgnNZmF1yx5tPX6nUA186P6R2nXcOJDMyegiGhka7iHVGdNGG
6nWcuep17+isA/vYQvIEqRutXgc1NH6yOd/WuDb0CededobqG7Tt5/YlDnP+0dxdm2igBKTWk4yP
ptp/x7tngl0zrOCmVov51TBtBgmRV8DI9SdVVfoBrBZ9rhBkLyV6FDcCsaTbCtGCzuPVhTgPRIUl
IgLOQPJ6Iy3E00qSf4uiq5CGXDJAP9pAQGCBe4tts3lVuew6k0J1MLGXJIijw4XSM4sBoB1xDlPu
QH296vwvbG00AMpJDLbnD7aCPSzXperJ/AKJAOcXBcH2p/y9f8pBo2ArvHq92sw1LlYU8hp6CFce
/9zbvqYyKVuxbRJUWug5RnIzWY2nLyK6NkE8zsJ8EacLL1AEeqPipGNPAqC+L1yt1NVwmefIj1uI
vYKtI92ZYNqlIju8ebjmjcVm7//r9lqQJa1eXl4CVfLFJFLEtpgOf5+8xTJ+HbmbaS5lkMlGdH3/
QIs1dVTlyaf5BI+Owvqh9kL2H37uU1UjkHOfBZjGULdxHm5QsojSW7Dpe0qn7QhalE3xqSKS/xp2
DKZhqQF0bZ0l/AFH+TuVADDSgWC3ay5p+II93IjHT0/e7jFOCAp3edVyukhe4WqdZEprA2IyQTVU
SqnFdfFwu6hnY31nrSCW8kni1HgNvIIipSD0hVBNRDieEbin392tlhdcdbHHfH3oJb8d7AvpCYue
Z3OCKIYkqkDhX/7npfzFWt0xToZLOTnvx0WI6gVGSXyHNFL6OT/KnDtFFTWHkVIf7A70Ldft9T1H
S92Qw14HI7Xff12W3Jn+z5rcBvAUPCMZpbE58vOG2vo141+yBPf+/RlQSM7C61W9zR824/KjGTll
HhbZhjxw3h0m87ODr4dGZb8ty+yOUX+cJG+q6q1F1MGj/Z5HZ46ETZUaFHrJ4fzbpTe8VinLNyiL
GymFEjq+DjIO7iiIC3En4HADCewj/+L3KApsBUPyFKqRm/04iw4GCX3CEzFKrlQlhBILUNuW0jTZ
EzpMU2zJS1em1oiLlgcWSptD685VFtjGIFb/BHCO7xi3J4GblWniqlfYv7F10kQzfacfQm74QpMi
EHzFE6kU+GFuBu2YlAEP5a54aVRYdx8BWK2HLrtRaoQSeDtB8mFpE8jzCO73D9clyJhzKFwaZfQZ
6kAcnz1Y3Zdm7EokxfFnx4P0ObH3yZPVWOroTThhJ87GI2AsuuJPQDP1Rpy1VpIPxUczPZTw3Hew
otmuDbkiAzp5bKTi8XY3dKGmNHltjy8zpMFnA8AQpBryefGan83Bu1fExkcsxPTW/Veoj8INlLSf
dTvTX6jf79xrZbdI2K+R3m4DnO/HpWfSJGLRaJwGJAwqSaxxIM5ir/9zNS+ZZ4aIeyZi69Y7OySI
baTCovpE3nvDn+QZ2zyqL9EzKPlCzI8a76RpxHEaEG0sj6tAQI0W4CZJYSD16/7zDfdJECcMxA1T
sT4p68p4fkFv+gxLE9uI2iX3MnjTizaYk2z/LXiFzyKmO8+NFsahdcT212w5ohxKYG3zlEAos1Zz
o9mqzt04E5w4Vpdy5TVAxSv7acY3Ia3reCBzV0EF9T2SYJkCtkE9SUY9t0jewzJyRNjIRAufB3IZ
Uyw0XlcpsPY1ZxfCHs+UlZ1XjP+MhvQrJHBN6tlqZ5aZpu67FjeAx6TXLXAGj92D1iKNqCATt0xx
XDpKxfRXw5li3TsX1EVfFWQT/QA2lZkFsj5t93B78dQT/KzcboLPLAKOWHtCO1i+pYnNcuHRbZir
NbivvleijuacQR6/mczBqhhtd2aw4vAAUqrbfJGb1CU1ps87lZ/KIida889mmYkD7nwOyyeQmuac
bzn9q+PrP4vb+OZJhJgAp2VQ+SXkzfDdkOtYEcLY091PkbM8PHU7Vbc8yLFNVRNTf4oJO/E5QCKr
ay/e6nQ+qxbyOvKeqDr9/HxJr6COoSsGQn7qNXxRhUmMGjuY7l//k1TBChA9z6OXGGaIk/H1VbPS
Jlbmu/Lt20QRUFb9NnCjFpjWG3D1xN4MYWrad/AoANMztW5pLjWLiNLW7dIfx8synPwMqBSbSR1k
tnmPLVkQzH7IQtTlfW/N984+V+FEKcpehABe5SF3gJbrEM+lGIZGGe9x0DEqLupY252YOwXzmfO4
mKj8D7JfJZouiGfkNl3a8wlE0dArrKxpoENgTo9wDnFCNK0ybp9OVNLZl1qp6gXuQOMsJ6li6hN1
eDtPtXBEiBHPIV43T7qkJ4aw6XhgefhtA2SiZHQiyKjmdWmD221l1YWRe/WNjK6qOxW2LXcyLty2
5Y+s+ejVXVyk1qh09IXk1YCZIfjwiqplj0GxX/4MCJQJls+76ewlppo5V+P8EYVO2kevxoXp8lTz
tP5p7juI9DUPz3nVOG0RrXa0zog5oGgat6y3gafxJfCABCb3Bwsqq/ovOnYtRXyk3uPDnuZXChQD
J1Szen9YQA1QHZqh6j0xIj7JKmrn4CypkNYTQrkua8DiK8E2RlHb6fXzK/aDbemXhRgriTVu9F95
2aeIFBG0A11T9G81YO0FPCAykZJ321xb/mmkykQsECXEaWpxbwotPTqoRLe4vvNYRariLDw5MZPT
gmyS2Shc9R4aCVpDq6/8lUrPtmpYg4U2kGe6nsRv09zk62umcGM0i/n/bM71dC7BxE16cYJLVcN2
Ri4MMb3Wypt2tReQrZw70wzauq0fkxK9I8G3LJPqTBVKYBAVyvuTJ1QmX/cbZzr2z/dJXQG9Lf/d
52yd15yQIQUvAwezXurDxSYuglfmmv4YFzzq8+xfIqVwSzPEhkww2UNFlI/S1xOT2oO5amvJi0NL
S4NBejbtSV5j0Y8aZKq7x0XV3/dl8Frau5ed6DFa+2wfRiwi+0KOtyXC1I6S7stx/BUQT8ZLP9uK
GS325wRjXyphbMhk4YeLVY3zrYbi0kJhig0CPKvrCf37XUTJtMkX/mBmhSIm/oGMjQjDIa1heJtV
iRqct9uTAPlRmMTDEIsKI8gFflW8UnT/UT83CfukZGtA8phNGejqFgNpllKDKDzeWhZs2w73tWfJ
YaVDl4goWhg0BVf5dXWnnIW2is0p+Hg70p7ic0X/7Z6wTJKGIuaTrXOkmDuQSZoPASQj7jsvxGxF
9JeI82ZiDrMy/l93gjge3NtPFZLDGWliV5fHfqLka/lTbsUE/pVBcQuAwneF4vzLDA5URhahNqiU
d3k5FFU8FqdqqENOZiLiYpJIPatbHMx3vgFnVuyrWGLz27Ip2mD+JAuHI5Z9NzSx2MHKC8S50/Dn
+hkGvwv21sPjWDVWgtsWit8YJVmDAJN7J2NDhuYtIGQeFdslVgevjXGvzYcshagUrOwKECnL6UOJ
fHoLm8AonSJAKciH1cMPpXsfXgLTO2L5td6/Py3tP/a5HGgKjzBxft9UY/u4TUqzGwRSw/Y0Pfzh
7UQ3eSPq+VGCtHCD6Q+/102YQcu3gAs/bezBYD7BXxbtYFZb89WhgfsFCH7kawlyF51Zv9k0fDsh
/aaXYkmVCNm/Svad/cXFQ0HWMOvgSe8S5uMC4g1VFWWisek2uQyVLDnwxfHnNUif8lzRMD4PrYqH
OGAHD/rA4w+IxAqk7HNEcANbUy8W1D1KDNgPrsq4JTy8Kz1Xc6cRmXlHCGbZmnX/MS2TeiJHZbZ8
ncJ3L2Delml5UuKHaDJfTpyv1CBbYTyEb+4v9QRjVPLH5HSPLRzkr5MlJMauyNUdHvOusszrGjBT
9neoxZlUnbdlpPb3IGGLyNvfXfvL1Z+tAS1XcgW528Mrxh6zrNTyV1o5khkuZm/IDsYnyEq+1L/9
7Hh/4xyo3V5Md9sruCq0devZohicm/HacZ9Ur+QQ7zq9WzCYlfpNizl5H6zJt0sGPKxVVfwyoD+g
ncLAD/PhKBmnCu/94y/iZ/lPivvBQKgyDQ071QAwCjKc7U+sjie6B89Ol7Go2mH6Tz9cgR9EmS9U
0OzWn21fQqK+huzqIRPFdUTYuVvZrBNLV8WrguUlw0XY/yy3M+m1YzyXsiW+jn4Nkid457E9rMVS
141f78zvMnX+sAZXU603gyx5jf8wAsD4X7OjEHaPUkQXvtVwc92ExbH0RoCSywempFmnwEK2W2Zj
dX5whBVamFitA4spG1JorcMGewh2gmxylS5TshGOQhA/XOgBewXFwNugv0T191JmUDai8z2kmz8V
16hgbSpn2b9A5z7HD24PMbzX5xJk79Hiptt4fslvyIEy+QU71Wjn3L5o/h1l+uyGx4OCemO+hjKN
7FAEq/5/5Wybx9807SzOieKAQ4M26DuTesry5HzQa8MVsjX/+/bJp+ujK1XlVOXKYQnOYp4sVrxV
Sgv6FteTnpdYvtAnWa0TIGy8O0ziIjDBYLwxaWgjvi65Xv2fFcQRHzgTHUCmbWnSitZbfKosLgXb
lrACGY/YeWX8kd7UuMCFg2ntcVxB9KP9bw/snzIkl4q9fMt0C63fnl2HApB6Ff+rqkBW4saDcclL
4W0e6GRTCl5RzUSovFxElIg925YcnzMl4zS2FNLZ5aahBK4X6ogITaFZ02ySgu5Zwzj8RhEt7glP
5tgGqf3C0LwGyY4dImV+pZ9VZTcjZdhyvAmpYmdl8f+5yBfhgPFf3MDlPj/AglaPxQ9PIb/M+y37
LZ6jxNni0a30Rd1oMQbSFeKNXIkc5/AOR8LmaGskjnLSis+GyQB9DbK0Aa5vfD4Iadzp2Z77DsaW
1VqxDJ6WVOGmQUALiptuErPSy9nB/Dn5J8UWtegxjWaz5IucH9dvClvywTynpUVE3DyflO/xJA0E
GSNBHBgAfrT/9XE7jx69mBlveLQ5Ci0SVJ2NbDDqeTYmXV+JmXrMPPMKC+KwOR3DCvIt09VOja/s
45vSiWPfzAhauVc6C8WpRuGUrNeDlprj1EEavmVrEJXtLy19BnfiAJB4kjwPYYslEXEywkIJ5j30
zc5B/nYL03QOqVDb+euoQ5bGtVUdyk6OukRZJEjxsn43q/W/plk7GqfwWwQElfA77jI8lBJr1QtB
iv/ArMM72OpucBaQzHGzdeQ+XvMCL/WNeykClOTLXBucu1u+tIN57z1NW76JzU2dTUuo7SMd/YzF
WBYemsVOQdXFphImNlpxzFK+WeI9M8DDVP6Rctm03P9gwUtRIdkiduVFR7hghL9mQ4wUe27HxXgH
ry3ofzoDrUwXppBHRsKw4ahTll1Nz70R+9j9l2h2uMb2pGiqjdqKytECEi6v3vCeqeRaoO+3RaJR
Whl6kv3naOa0Nk0RdgSGzQ6QmBTT9pJS5dS+VaiAEV8TGNKdETx/0NZMbkyvqX/na9tdCrqP6Ia/
cJ4JMcf1gkBO2DyLmHG8/G/o9hiiy05/pjNehA0A/IPq6AisM3ZSipVFpJ8ZfP0DquNvROW0kDBi
SvKExLbvf3UBTmRVfYoahr4FXcwWtvLF6JpllGbbRynfaTIF1W2v2UH8yJxnLsJf0xh1pyeuRtJt
ssLQ2Eq+zxzWW+STpLqAHr/be9QEd+zPxzk3K+FnmWcDKvPDC43hE+1x9gRFlEBX3PjVR8AO4IWR
WrusI0NIW6N8CHcu4QdppOcJ8hsNThSYsnwyg8MpPiY0EdMoVPHq24Vp2GBKF+7mkY6sJdqB9SEv
OqVr04/eSoUTcqkIfTWDa4K3JUOSzBXWpPl7zR28q/5yLowUP2FnP5DTnalOhPiPClU8rma+jUhO
1Y9gd8XaL9EpUD1rYWWZfOYiHIOrpy9f9PRbWZg9bLRZ2XYqVGh9SJpSC+zZb1aON/iOcUKfB7hV
hyZvdkl3AhtzKud7aCq8ewzyIqfeMHUW9lE4wByBUcndQiKeA1Gwo7mE2m/7E6GRGgsdTuysRCs3
4YfLzhmKSh1r9aGmvqFiOmUPXwRwwShPzQnAwSLySh7CxbiY5XzKpu76CqxZyqvcvDUTVecJAcb4
4tg2O+zcyxsJWM6vKiGKDQRqzmnvzgjYu622kuO+EA6hsvSxpwqazSK942pXz9R2pcvY6q6r6SXo
9+WSt9hDxKbYVUTAlkyCssqArvB79lZYM1gqy87gEawFT3IGE3pAQcDS8XDDBQAm1OR5bkXBCYRF
j2MecpyCPix+X/Ay9a40CSqbfJEtZHDr0N9s7fQ/V/ebo0euvMb0p2pC1BevYohwBKwmtD/q+qM/
NF/xo3pwbp8pGDPg3r05qD147OFkL01akm2YM/9v6FuCh3sj/YxSYHwmngIsTzkCuDL0xl5RO8+n
oqHD1/Z1hGFFlPolZdGrusDNRIyEkrnznQvGZSA63f1O5aN8ndHITAVLxGNcNu5KgB8sgcJplc+F
M45APHtITyagBPOA/OeLxy8vjAbMPnuX8vP/W1sNAviqSGx/cwIBSPL0pWfCOQyXv2g7Tuh6/I3p
LOA3jLb6drawq72xKdKIvHja4wR8zQUNpY6nQlGEE7byY+azIhpovM86vV55FxaUy3rhyIIqeJJN
fOUKEZ0E5ucJ1OMDYtVqp+FoD70z2koPgNmqQ4wo7IKPyS4dVWNIK9Kf1kl8EoJ1jFjtkdkdEa7j
bFbKMqsaxNW8A4E/mvWhxS66uJzDoB9pp5qp21gLvyiDC2qy81qeENkQPPR5YFltz7AfxczxGLCO
nx+7ZfFm8ApFP0fHbQ3bWA+GsvUjPxKyIPwhK3foWElCKv6z+Mb+Wlmmbo6RDLWQIUNGd5EzxYX1
Y2dzCr8VnCdL5aOc0Iou+ZV8Su3iabVSirZ4/UJzILizsHOlU1CXbS4ZkB1uvVYgpCq6qxzX4DXD
Mt7fqt3E+VYk0dyxHR93B4I3yRLFCn+ryCoDT/ZvHg5NdQb71QF7rvUtrLlr6k481a+h+072KYFQ
wDUuQ3MLfF3gFLZLFyuRl6pqaHkWj6uOKLgsira5A4wANuGh5Hi1Rd3NszDdtQOniX6WP2Fs62WK
hMR7TJjOHhf1Q474LDajYzXGXtxwwMKjoY49CD4SRFdW6EuQYAZ4rRUH5nvc6LDYE46DHIvXBpFb
3zeGYdsMi/c5Opr01C2zrutWj0juNP7sDYoMEPPpg8xjpnaI9IGyLRBssQiuruRMwGd7CzO0btpz
jfif/ChJ/PNJT5NqTwjQh33lR7123y7W+W/qZ5MzwpZ838tzaxolWk8CiBCRxN6X1TSGFkORZlH0
rINVW6OTYpq7prc3/Q9LCsXC3Vom2W/6/g6+flZ7UZGp0hglQ0PEqvBeQAGd7ZKNVUln6hfgXjU6
V15irNz4ZUuLV3vkoTY35GYY7jpBxVkM2C8i4f9SdLGtCUpvJZSyjd0249IaQ/6335gg83ExiIg5
hQUTDiPPkVSGJOqNBbf9Q4ko/DpYsP2cQnD3a0aMaJ/l3Nu/RNPPw5t68F3Hodw1esbPAAvQHySV
4pALmqSJuAq+j16w0iwBk9nt5kTx6CQWxmRMVmdq44bjAybRp65KgudZJw2h2qU1js6KTSj4x+x+
NCqFDnAjKCzp0lsy0Z/2ujcw2AsHcosL3+XWqYT/iTD7oyv2SYL6UkQblMuiFjTSyhOOuHqSwRPX
00EqTWO/B2z7iRXGfE1d1HkqnqdVF4ndQNpzUmRkVfM7sb2Un+aiTa9bDflEHnMbLDdldVFNgR8S
10s/s+Mu7Lgb5D/dTwclC+a60AWhFpmCuxCIvpfkx80uYWfenjFv/dr7pQ2dwkvgS2a5lMaMNVbd
AZiNE1mT6zgc3t+MB+ZBtpUAh6DbPUrcZz0e9x3ZsWqJRI0n3w2YH3fZftuiT2774Gq8lrvDh0Qf
GeYVeLLqjcAL8jSlngq09raJSsqqffgoAIJE9k02QSeowiFJxHeQYvz34J/UgrUzlftaS4EUc67y
xkmMz/rTRLpvpviDdEDGBf9v9g8rtOmbRwluVovoeMGEGoe9ZfVWUW2n3srweXwtvaoE7FTep4nT
5iufqedpT148G8gX3yERzHCClNzGiBH48lLt7V5Sufm1XzTZ89Cl4n90hGJ4sStwzix4PH+xxGts
lI71L3IsXKXiud6GRzdXZ1nvspEQcEiCLxBOaEYiFe6PVoau/AUWbkgMcDzBwsmSZEq1/72/wzkT
vs5gniHRN+AEIWMykKZNqhVadEp4wEFPaJXXoszRiafnWWkqFsToN3DZxs52bjLLPVzubUCoDdcE
3YUMez8eO3Y9SFr98yhECS3nEBEI28NhWDytInNgg5StLey7KSPdwUcVHN2roccC2G0GSERrGZcS
ipYUK5y3fDGgY5eaa6+OFn56/rmBUG5KCeN4AJwz1Lz9nHiVYQ27a9/IYcNifBg5eHs5Hreot9HS
wHEodA4zOqhAImXg7ql+kzUmNeOFb788u5Sm68qog3ZLsRgOvSJiNkMVg47FbkKghLHEXfkL0F8o
Z9166IyIledHPMNibx5Fn5AtE4+3Vza8dSpwvYApfQfUtlrAqrvuvA9PCsFXf/FizEb0AixpLvL1
8chTNglX6H9uqx2/0pbtv3SEmByzjk8qe0N72+EqLKxNm22th3Gule6XqdjQy8Ohc5C57Z9ENgwl
24IeOoTWFnXY+GplKbBPlvfQ+FARGNiH/F70Ls9/eK3vpYwq3zv9Y022f2VNhZlZLQNO2a6zgdFS
dydF6AobAXrtH9Lmd3DlCrdkvgli5gvQh69IDgExW6QKzT8+ufTGFjU+dW9BSjwgJhbUHkYQ7Ymv
C9v241Ve3ypBSSJNLyDI4DB6DtV352/wTkhEY57Fq3KAAiB8DpKPhBq16SaBmTRzEDeU9ofRuQ8S
YIH0UUtME6ZwDBr51OviiH+NOHHps6n4GS1pk1eJq4ZKaZ5RGVniohn2BqHKcH8QU0sow/L1EjDD
IoHPL8GOqZYivUgVdtGEgHgf2Hne5LRbEHfeoaygbMV+acJKweCdnkl+EteK5vXtvsMziVOaJPKQ
XCDcjxUTJnNQtiBUaCsJo1xnNmB4JIsjNg6AfE/fTx1AB/pHZP3a0UHYVYUq/HNzcFFdAIooUSkJ
y2UELrHOj9SZTRTEL4kyEe48oDImepqJGxGrnYs6GqmHGh+5rSSH9pxadegt35dr/W5CPcIP+VWP
6EH9VOLvAJjZtO6OmqQqdfCYN07xkkKlVNNH7ey9umZVb/myZjXO3FF7lq3SwGWC1KcqA3blobxC
eZ13zmooBaYsNOkVqFEA29G8X3Yez+Ze5HYOTTckPQrhsW50UV8brnvbR8vlFD/Bj8+nKFpQ2Ctk
VhBmh7SVjdrxsCTOBxD+SJAeZCWEOvtv/rxkQMBhkY5v+1pMJPKk64LGNCIUxmKwBrW5HSYxH7bY
w9kSSuk6tggAHdiW57yqSPM47PoEiADdHTqiL/9R5bvn7VQ4SFAwFzxysRccgplVX8ASUoeAOjfF
tmIqX+8qA+NBKAilgV9XWnaa/eouKQ31cHRiyf1S2p+++rsPgI2c/n6XhAXg5IlPCtWvwqKu83aw
iRyoGXlVYjaiWoXuW3AwilOC+ILC0H1lxqxq3gslmnJ17zbwzTHF7k1LaDEhxnWmbRKA6sw4srrN
dXzOqRIdd4qmQvmBi6EX2+r2J2zy3aGo0Gk4SooSWXf2BL5dazfEjTiOwelD3pHLYoXN2xj20/O2
id9RH3TA/0ZH6CzVY6PYJACUPN2Iw6Gdqyt4/eJ40mJUsMgOmbCeGIHRJwaynvaEsvueIcG22j1g
KIUmIVGXpmP2mQgqNqIYqC/tSrgOlzU9HEhEVYjENPuM0QnI0dCEistt0INycnOUMNmsh5/0rcDR
E8mLPOY3zwsaeKxz0v0GF/9agkv+qLetB38jJR6I91cp18PHqoZMmmZOJh/qtiWzIoSl14ljOpBp
pXqaOeiqFDybaOiHNx/3ZmhQsm0tZhrYFkw/bxzz7DSjVOcGbW4VKMeZ7pXi2ClhtRilv4lqn4Ww
VfmjtLNwdv0Js5yQg6M47WNiCKvlrykdlwsiIQ3BN9PHwtHKCCNkV2pVdDGr5cw9yF2UceAvAidK
GC6ecQLE9yqEeBUldHdzuybwxsJ0CLE/GAw6xAip/nZJ2rd0i0T111IBu/MYW7VaLAztu1qfHRZi
DGG8t37JcgL3X1NZqQioRHFG9r+mBKlBfPq6eTJeXZSTOx72ynpqMcipc8+zsXt8WoGoy+c7GUwE
siEO/phShbzuCwP52mSQX0ZxllUuPnU7QtKVFR9yndSokIaj7kzZyCuAQy5nUfnjnIluiFNo9fDJ
8Mtv8Dvv2+dZzHA3VET3egU4w8uvDwhr+3x9R7zXz5IF3y+l3j5+Z1FjWTSlWOEr8iy/X53D5P5i
QDZax2dFa+cGDxqmWgJ6LuppoiK4Mpcj6oVVPgF6reufujcsqNwWVp0XEL7SRqHXiLbDGlRjwZdF
ZgzJCuedqSkjEltHIDOIdxadje9O16Cr4LfWEHWpRyHQBLvVbK8n7+zZO2F5w9OajNhYLNMItYjp
LfYvXo/HerciKCESNbIKMe3L86zZnWOXcYNc7oUQAqs6yPyFmpqEOqtohhzZrtA5ppCJ3PfDgPRi
VETqlXsrsylp7rNSpIBGMOonYsD2Sw008tER3afMXU1VVqcOT/a4wZ/8B4hZPqLK5gpawAEyfz/b
XmjvsHMBoMw/Oak4STOAZZ+IS+ZfK3NKCfTW8SO0N//wj7sTVztBeeBGtsQMld9OIJTjjK8eLfHm
yfm5xGPmREs82L+yBidz/pPnKXEJ8wZyQg47KTvFfMi1XdRVPZ54lMZEv6HusyBKKCzzEn/5DQla
i9uIM3tKmukNoABsP8LZtjvPfdqkgXWM1zvlWPrgb1YjgWzjTVwJqzvhAM4G604jB7hszNK00l+X
y686cnC+p6d09CnbUXM+DFOsW7evZJKmlE7kGKvUkR5Fc1VwAMa2vIDNqyxbZ6FG2MfqjA1HTayP
xop21vx72dgIWqkUnreWonsuKq4KXM2kSusWqpjFO56qlqh3vfDab85OxonaM0NI7WzReTMg6Ay4
/F0dfm0Kz8Wc2T0yckqK8yCTXRiZEH5mlgWKEzc0doWggM/bpZuz0qczNgCX1cB3YYMBYMGJQy1H
B3ieTMYC22gMQ1pkZH83qeoAHJSWGjHgaNlHPTK+NmQpYTT1FOsUYKUaTG7X7u37BGJ7pWdI7Kn2
4PVhf0qey5r5McDqJsdlHmn6kky1Bq44vXq4Gm3YiQ3/YhRMh6OBwJRnX76pr6XyrH3Rz8DkqsAQ
9/T0Jkos2qeH+rC9XymYbpevXO7Q8k8yQEZ4WvD2XlRepKppCEaAkKalRZ/Bw/dAtAFAh0OoMoTY
4BBJe3w8TgVujDE2xOpErz+KV7JcQCaa0kTboBalxU49z1fAoNAuadSHUk/LaVi98k1ORrMpGl4J
Lx79cksjloVm6ITPS3EuzNPgLBpIwcPCWKLzrSbP8fzVxq5FdpWNXSiUq7EJgbhpxi9JIvCBYbyZ
SEalcx9INfUDpxiqewmiS7fBcvXANpttVntQ4GRHiAjYHFFWbWYV5j3fo6CvQBr/UFiKHPq14rsi
OlNVdsSqANTxbZjunMbd6Yk3ORcbawDV0jghK++QqHgXH3L1GEFxnQ+11zNsjmtJW8v72+VD2uG6
k0l/Qy9Asof/mYaZMTiPam5rgoqGFGNiRhMhnrM7L7XSsMBQvO7Ml8ZS/gSeOYDl2YElQhlECni3
lldln3NDvVpHikhKOLi5B+CngoRbZokFGGfzw1vmiRyJpYk/N7+8jY/mcW1cgOxsWCmrUm+46xRE
UknKUWZrU3NYM+ZnrXfKJMp8Sie7remumIeL0LtdYBbSg/PLpR+dxEZSrH8G1+ycwts6k/kkAnGf
EjairBFekhehSZiWt22qYIzTHtvOf0IBgKbfs1BZxXatqX8pt/2GX0xeScNAli9KtEJlPAp33Raf
cguFQty5wqGzKraRwp8ZIvJ71/EZZkjolVQj0dVecqQleRBrkoFmYxtrzla1xj3OmGvFV0gYo6Rc
XwQQB0odQx9X6NhFFrvc/jlXUcNIvT3q99dCaSsWzEtVV9lJSz81Tp+2lxs3gqfdHql97ukLsvrw
Fhj8BjIRZZ2JuvSBWJ9BBX9qsbzGSN8TfNE78SNwn8+mESA/iEAzNSqQ97lAv8YX3iYXS8UxwnhU
SsWi1ZCndxW4yfEfgcS01BTFbw/reVcznL4GMt0rzCxp3P1yyqjp+Sj3ZgqarO8GGv42sY96e73E
2bKzL2O7OGk2TlpSWfamP57BcklnLwt2AVNNtUig/UjeIm4Ca/LmldWMxxDqCnfjlogZmY58sktv
m6AWaSWcDmROs4cF5jbaxIJR9c7l8xmU0zkCwVvdR7LXo+BfqukaGKd+Rj8TSP71hDmCsrZbjSN6
+LgyUQlcM+hmUkkohrgA41WPFe42810Y2tHXvZtzr7EVVRavzO0BYN5r/evpisKgmklL3KSnuDRj
LS/FkU37TH+tnAOamN+VEbAT/apwv5ZL7dC+AnfcZCLR30K2J9YfkkdPBXZlCAJ19oDD/8z7jivd
htPrRmQHplplNEarBcoyYlovoVrSq5lpwBf256x9BP1Yr5QlQqIDLImJV8b94XAUEGcQ04MTS2rC
srs8aH+5NgymLAvprxc++cXu2FEF5oyhLxvoZ2WkroORWoSYqLGtnnc8UkqHFO+YLqvd2DhXzZpA
RpsjkZcjk3O3aeHE2oPL3vLLP/ewIjUErfUT2JNT2cB+Es3rz6FjZnm3VslLqw8OYFhTNQNPEj+c
xJlG+mqAkTNAdnFaK182iHIQ9XjqzIhQufk8V4dt5JDfHqdxZt4QYKMKO1dOaWbYROLUqHYggn58
AoD7fepmvPWUvxr1XBaO9u072lM2Azus1csLb/rBWOq46jU2BkywevwRH8p2UEhhGwvUZwB6dZlS
SnLKQtalY4dIfJfoiV5UYKHMml/QFE2B0WYVFVCopLiyvhBzgAFiHomXzcCIKWcq9Vg0do8WV5xO
5STLVugYK++d/A3Yr5XhywUm8bbkWEMm+5lVBJBpoJW8naiT9vH6V1lXw3u1s3M73d6fIn+OU5Xl
23h1KlAR5KpP7J2rNChCMvtcDhrJfrqOz0nkChJfgiAWPneaJivhaXB39KdHEBPAHs++VNRNPKzL
qteb6BztetufZ0wlPjNi8N8VpmmiAV5OCn9wSARMzEeCgM0EKJ/0jmInYJAtlgS4doyqjA9bhc/N
dm4Q0/LBj7c7fn/Jj8w7J3evlUWGC7+ifl+DPxKvP0PZ+xa0JSrCfriLfWHRSp0prBi+Qr4SaoTT
Lbjo41uRdxhWMJPaCtEhI6j/icWPzjoJAJBcX2vK2g7YH4G7AJaKKtlUhvR/GXicNtd/LxyMU+hv
mclAHOsI6rxq8fppxXZkZtdvy5ygBBLGwqUOjo8ifhQ4qd2jy02sg14fNB8TxiSBLswxpfXK1IWy
kVbOiAbvDv2b6OdzXXZofJTbcSshDR3EMgexknHX+leODgMM1JYaagWsnWnVpSCt2RXL4V6/xshk
I/kUqowPjlBBdYUgcsF9ExsbVaENACiHSGD1pgx6t52RRImKcnW9654aH3m4UEErbRXvkQp6foXU
jYgQoGFRzake69jJ1jMmcMWv5DxLmnqT61MgZ5RNWgh0Vg2B2TGxPRFuWI4HhOEk7QnROmUlqSfB
VsSInZVOKSWEA/5HsrLlkU4YfO/sIpS0oOl2WEtfabfzNrTxFMNbJ5m7Hl/pXwlpipLvYUdSbGPO
wY4eNPFNdqDQ/wqH+GmQ3o4NNhKfvW1xBYxlj+S5f+gAHq23NPWOrPsWSpcMB6GRsh/mYnkiitUX
BGFX5lZfsjoQtx6pnbeHeGxCGguvbmY6P3KRegqK0tcE7bghpjd2ZaU2XvdUZoRchDP15s6sW7rd
8zi5hHND0X9bvQ0Pmmg1K+fCMUvTpsut3CHLtgAYYmV2Q3eVlzmx2v8VW22OgOK+pbw5mPrOMASv
0NWxfTO9wSBOuyYEKThpRYyBLca6xmaRlWuM3Drhui1S708dYzaf138hAo/1LVCrn0wyOx0/5zis
NUbS/n+RzoMPOYeZRk2jT8oS5Ls8BbEWB0bcxZ6/Q28NclNfRACOhoSwUijEQzzUrj7pV2CZM8/y
OuK05ISbI/abem7N2r6Y1aiR3lV4mZHQFRInde2Yc63N+tFSZc6gYCQHQWk/VoIT7z/3GF8ZHreA
e6BxiHJnOvYMzKMy2gFf416EmFzbiJ0W3+J8RZPYNVuNF1LjcwOZ42RJrnuxSQ18C9LaPozF4pmW
Pi/VfxzKTGI//2Y/o5GFhb7NMbKhTS5kez6C94fMeo9PnOXRdmxha1PzKo3sxWL23VLPIBuWXMYf
oC+/tdSaGGEBllFkEQ5JsXjfKz83zkghr5w44E1MdA5v/7zjNpt897Hg92G2OBiMVqi1sclS0Q3G
yN70+B2tPrBdymIMRH7OL1X8lV0Q/Y7kZyIFhDzAXVC/q2+uZYzC1Kv90C6X56xl2jHU0G+Co7yr
5EGHzg/QY34R0Sy5rroIzqEGkT9+mvqHlAVTgMN2I+xEE2Uap7WUcLIah5ERj0Atu5hcUT0RqJrP
PPmYMDmo2T5Pwfu+55GPzLT0TcwpxpyAJGWL1KcU0n5+/TE7K1nD1yOP406vWyAitAJBMDMgl7U5
04h2pEjwaIImAvbJqf4iyMs+AQHk6DSMMFo9BLL60blKklvlUBkXFEU3kehScgVHvzpoXaubDZfi
fyuPDhIGO0PE7BN3pp1rY+NMJfpgLZyM0EOivPoEn/L/YxoK9Z0XV0u5wV3NSRscTT34lfyjYSyr
xi4vj9gM2r3uLkn0RkahZISDJXFkWSuwOP7WN+tvm7jy2mJ8rcPgGnfs/Zyb4WVH722I4oP43t/D
8qllZbinlLE675fczQjwFJviG2fuKq2OUrR59sgXXBbKL7rfjsAVA9NwqjrRAfnQMIYyFCvUg1su
LEQ0s4z5UExNkpfovGlBEkR3YWREWSjQTr15MWCAvtwCmknD+BUFDM/mFLWaf6bBDeXUO1ymd7LY
5notipxgDw9qmAG4RKr/N8MfeucaPiP1a53q5zArJ60MxEhw/zxqcJnROHGdxmDNLZx1z7ZQQGyC
VemYE6j35JH0I355+zmypViPuYr7jvr+LOb3up9iuoFOJzhaxe5ofEGZBQzRxVs/vZ4rBVD8INWR
BMptsnyFmqHOS36bLnfjm9zXUUMoDhInuk6aXvKTjp4PkY9FS5/3QS+/nP3d0NHyzi97CvWtkPgc
fIz4bnbXL1RV7l4bF8y+1/sCJLexgcfk4Qbm5f6MUGA44jh/XNhJhxT/Hi2jZSKCSHsu3KrXMyrv
Fc1KYPqPNsrbSJsNNljJnCAWe4NgqxJjurN/DAEJ8VXT/tx25qXbECJUW8ByD9efZ3IPzFaKzyxq
YcsNc2S3sJ2hjQQfp/j0uDaOl4j3AIVm8FHHq9rrwS+fqJWag1+xaf2s9srTcpbnnikh8k65yxI+
qeI21srhOp2ATwE7XfkYrmom8PoJvEd99xre06kzistanLzF5TfrmiDbzVKa5/m4bXs86P5cJizu
Ka7m9AV8nQjbcTh2xZmCxCX13BelazZPL0liWNSYO/Sz/m7/Gj2etfvMe5qTYKTpm1M872HlC5kp
H4YpccGki9gK8s9kKPzDi/ZMSsJm89zvpW0lH+r9zSYYV1F6XA3jwhqFIw9X32wcMIzh0psZRhAw
Uw+cMrdKghRXazcsupmAvF7n3glRA5TQ27EgflFJHNalo/TPczTw5cir5XXzmE5hmM3DtHWWnfOg
kETJiRb9jlZr0dCHxQpRMI/YHB8BB3jjRC7696muvY4AC4I4AsJ8k5hKq51C/iWMOam2MJJjOx0N
EqBll0tAln7utnz1plaDd4h+rwx5QCXyqJ02WnKJ8VbFv93vf7ZdCLbQPjyHEkbiZSb1exM/AoXP
6vNwdwofNuUkuh8Bj0omLDLUCH/16eSIfRye90cqcyDAVOYU5P4M+sVKVUoiBpCjt0gEW2PHr7eM
Gwpvx3QL1A4ozx3ohaKnaaP4vuBiIsNVQuxE0wMpatnxUtpGIKJ1Bu1ha1p11OEx1LrxqaYLwBXv
k4j/InM0M4rpiuCfoDA8qBah7pBQhe2Cs1xlMQzUFaLO3/PZYHNDVTNNJz2omWKJVE2Avs75MuM+
KELAEZeme4dlNa1tjhSudmC31utgQINZdE7Wh+qXehXePUzy9L0eOdzsiVGcpejTVjFvcX+v5FuR
7Jl6bR6trWtRcW9cS16XYJt1RHlHyeGu+TzKVgihqApdhRJgkCQONVZEtURHnoccX7aeEVmnq0ai
THEVp6sRmueReBo5dVcENBoJtB04N7N0LnqonfxLK9M4hatQOWcqiMEyoAAr8x7YRQ5BpgTuqKNY
fz6+VVdJBIRDcTCRtHqPrsgpDsBplGuT7UoS36b6okMhUw6sZYKftxlIJtzsaRvjmyeKKr8SHZQY
xmeUvkK+18fM5LoVKSGmgnWmOWMa2XQEhrJ++QQUeK3VpdDCuXRcUt54qhzEopAwA60QBrY2iea8
7GjY1f8XcefO1+D+VtCXJistm2lSGrr7WxTHjaljOy4ncEkx/fgX2fOK5hFzZ+SA1oEB+bV64HtR
PyOWINrkcNNYk4ZSIXF1P8b1drreXpMMJsFdaHPq1XaT7P54dBCwR04J6kipb/ECNAXHFN+LLJjF
lvPvznCz4Mm10Ez3R5hG1RNDDrrNJrdLYqF3gfrMo86QyIH/ZVht8OgsEmVAwEOHiD73vBFQV0kS
U6FHI+NKHZ8r0m09ruJuTXosjWxq3P6r7VJMgkOfsJMOpo031eKwW1Sd3MmBX/bdblsN7JP8aphi
adqV45ru5nmdEf+Cb1i2fwEY0a5OSJLrOuB6qXnuDIGqPrupp8e1OVV/ayWDSl4hVYdk36ObC/la
pZVbHl7tR6F1Z3DpDvxpC68WNW8j2VhgNqY2dN3Bkyiu342Ze2LShqpnWGz+9MVp6HaEMvVjQj7O
0pk1WWcKzwbjh+FwTgDmuvbojKsBTxlsYxXb56qAwDwVleizHYxOAj7QUJbcZsmeur1TTzU0uU6h
zNOq+s68TgyX3N75dgCZUuQPIzVvtyXmWMBl8hIKF+RIWo2gqfb/BEebJXXbkk7CmgNCyQ1jbkJz
F8dTG7dWOwx5unClJyWzKODdBhgG4CO7cKbzz+yz5sQfp87Cu47CyMUxjOAsAQQ5BbObVFQliwvD
TJXQP1wjV9/tqq2Q60wnHoGbDO56RJwfz2IBbTAGrlD/DfZiMo4m3Nyu4l0EphkN6HekTMlsyBbY
qkC6XUyboU2I1RjHpc3Tn0nDFsVeItzh5ph8URdVSYZ5FvgJDhznfuVOPFYGp2hv8+qrarWnfr4l
bkc95GGsobvX/hwlZ/tkxSHTRvweOnib+fPC7n6z37pTNoZDySFtE+OMRtjZuD7gHf1PFYUbE0DS
R56Z5KTxCoLqMg4ACOgIxywnBjYWVy2TGPDs5ISQXqPSZhEIj2rzH8sIAUOjFYWM5F06dIUbBhJD
AyJok6q+fData5C/vbqAA3ymq65e/1Asvq2cLnVWyNTDRFSmepoNcPhhhnwlb422HCUQ/2pq+ou0
UGT544dstTE+1HHHnbfpy6ac3MtdxgBJeoLrSPKXbIATVc294bgA1qph0KHEqEuMX8P+fDSHZqMm
A7aLRvavZ4KqK8juJdUwZ7QE8y59Ejq+geJA71gxr0eSEwq9KhxNcDrUb7qGmxWCjTuXPz8Tf8kh
mcKvVJDCKEqou7RHPFswrokYjr/16BRrLIwHnDQos5hsPy9aRWGVPew9dYGGwyOQCMu/ln+Ixe+A
AV0Si4MH2GvoN7qLpfPBjfPNooYUoTgikujmZef2Uu/yCy00qp08PnvHn3IrSfJUs9MUhMGtn6Tj
7Ujiu+qBnhewi99zMBj805WAVSyRc8zp2cOu9ggW/TeZB22u2OQcMCJ2rb0KdVo5jSDKXsdt/fCW
0JAhknRNWd79xLcECxte/rFDbNeH+JlykRKRLQQgFeEWKQDlheB4Zqi2xX6YtMBWbuJ602puL6kD
8OPYtxI7QlvtYLJGMkkebKzNW9MBUD4fX8/gCXST1nLM/EczX914H4buAgrRRImPB3B9Nhq+Yb5z
rRi3ww7h7uLUOQE1oQMwKIT7bbc5dQueAfAfHAnPTzfYdHj5FgHFrSAhciaVIrGJkFv0rskrRXso
2Xm66Ytw6R4Oztn4JxZLUUeygcG8632hY1ez8guQtvCZWlx5M5HJDhn2yyHTLvVzNcaznYL5fZ96
0J6qioWiXEn0DCwuApU0lXSLneWnIEkGcNQNMSptiElYkkSMiZypM7KKiRCuA3+ehgw+Qy0d7ztj
EDIgSmMGl6tPpgVJs89MCGl6Fatd5/nEmTCeU6zpDWxQ56DUlIbD2NPiq+vShdgCWHLHJDaPZxvj
Fo22zlIoT9tvoQsRjfJ9XnFdhi4YTCIl9eZb4RhzzrZCgXIDFCJ8fIR94vGP+YPTtCM4cA3ycgeG
q4o6tnFiBmVZ+OumNuD7DAa6BvFbyEo65tXgaIb4/6KaxZPfrQjF5GJHMrxLQLAd1y9cboTsFvZK
3GDWaaV8PVhByfKfTVNVBMWvTaTVwDDLLN+kknZwsVV1zH43K4W5xwSowy1hr9mw5pPRskhWbMVk
qRsJotUrX4rny/KblNP/q9eTCcm20jbTPjSyxh660Z1RJQgjmnldcLSsYGUd7i/vfqLJcw9b8DLT
A8nBrQH5TM3YlqdmEVlzkrAdNcwYiLefV0c6rQmXCRFh7ZPX3O+qWfTqRWAcOwQnnRAGSid6kt92
uPnVhevh5QHbfQf+qfRz9/EfYAQK9kg3FSdG6+6rA8TarVnuXQPs55aviI3QH6BDEx0Q7U+NpdbS
4PilFaTb8zTnnAf1JW7ALuH2MxPr0jNpLN/QUJeCewfiXsDGuPNwvzsPjL9sPXFirrbyHfGuX1oM
zQl8TvSUZXQBShULjzouU0DddIU5kD4wq73mk+b7gDLuvYXBlSOG8ohzocjwOqnBU86PAHwknv64
Tev1VtxzRSVyQob1Dp5x+Y8qwObdh3RsblVuQmK20D3ajIaXX3F6/Ltx5xn0M77GVIR4ng8HC76I
l62keuE3rseze06KMaSu8GBH6AdjJ3jGcITAzxazO1K0nMOJR10rS+1cdayuU8+jPYhjo8Rr6IJV
DcBsec2cM6U9bN9HmRcKEI3/Uw2sekIdlxiN2aCOxlTlcfRRwmd0Bmxu0BbMLVSRQSQvoLkeOkYj
S+rGLWfDXdTVqv79pHdHQtrjpCiFeSw4it3pxpGjCtiT17tSN8Y5Mrsth50UZ4mBMHy6TDx3jkw/
OI+UruF60FBkZ2Zolo+d8SBgmgjUxg2UI63PlRiHwnNdtmGnqOTq8rawHeK432CbbiVN/oRfzzWs
l4u3fkLjQyqA6WtbRwswUZ+k/PvRjCCH+3awT6a5YHF0OcTL9cxrJEgYsFRj9MZnsufEstO2BwHF
ahU2EuTJimafCIYzqaW/rc2UOohepo+Dkdvni308CQqN+9jBPCtezg8OdraL+9dJNTzoQTm/UUzw
5tzhTWeYOWdGrW9Ca8KKuY1jbwwRJQTggnJLgquPlL1gWwgqy6uPjRQgswpUmhAiam0BTtMZ0Xsq
8Gnztpt4DIwr1gjs6qlhoz6XYDOOoQDsw9ph+39ryIctDIjVpzgVyzEMHMNrwQE0jk6B/T5pVoIo
HuRh6Lv5C2tbdm4fD4DzmEiqcdiycn3zLYL8bL7MRfsYURQoshXJKxSUzg2+kGGhdPhWKL0DCGGz
jxYDnIA07uj3ZuLcHWxkLcW2G2LFiro+kOqUYyYRoxHJxkR91RUfWBmRsgg5OTQILIu8PoKqtn8h
essiSbTI0Ab85MgETaoY2I5ENufu09moQK/+TjLMPmVOJMknIcLyFbBh2UCL0WuhzxZFxe+CDVUs
rIbYxLZvVAd57EfqONROGUhMJMV3DMBZMpZk90+7iZ+NGiz93Lml38USGrlKawiAUwzaduNp/6iW
n8sSh6IuHGDlhoZX5jLtQ4qENCX+1C+8X4ibfuTp5kcqM+ZdPLWPL9JkMHF6wxAidJahWVH1lMT/
1go030WhjmQ4YHf4cjIS2zJmvTr/eG3AqqiQ5LwSjrS9ZhG9lkMHVD8Ef86RzAMBxzEtkyUjc7jU
crCubRVLZEo6GQtJ6A2keYWaCgD/qK5IrnK1hnSVo1mtUU2JX7+ci8X/YngP3TBWZg2HhrvyI8fj
ACaJzYzmjrkvomDHLxouNt+hfm2EaLqksFD+Tgd2VUI+qiAY7o0hkB2BMH58e1cAg7iLazHb136D
q3kRIKKIInoYELOOjVYOiVpC/HMCEpl6mZedhZKB8XE8MwnOcK9jqcFMtr+aMLAEt+k+lmIaQUv1
0CZeMnF2U+2yAHnUftDBp+JIGDAGxFk5znqDmB65Q3vxniwb6FgCoi4+SYScwGAzbLVEyawgf5GS
RxcfH3uvlIJAp6bu6mZBJ+BgqWDlzxAumnHGx2YSwSBy866klCjpWSwcMlmJZS802i/4gp6OTapV
vBxrmLv5iBWvZIJahqfBxH4EASbfGvrYNO5VFpV6hpKgd0XDjqNbeLr1/aspZpH3ZeMQJJRN/Q7t
Wuy/Q+/x3Q0nPOruc2y6arGzRjgJrFec0Q57r0vP4qdnUVCuW+v7jsnQv6y88n6nDUnyDlmPB3dF
JzS6alrY8qF1qU3GN74BW0TlV9/dpJtWZCWnxS8kEDYmYzHRuolLKoKgPKYUMgl0SrDKnbw4pNxa
uhD3w51Ec64fAMBiFTX/Ezx0syIOown4faCDDep8F9jIPr8+XssxSZZVZSFUztYLKloGTzPHVSI7
0lRTf1v3dCBY3ebOwyk5/Hv167mEO6yS32bttvJ0gK+52A3wKtUZRcVCNBIHKuO1Jlm9Hu19YzZA
0kxw0ZC2N8SKyjS0I+brs8g//SFvb66vrnjgG3JAloLfHuX9D5aDq6X9ojWy/kRyP0jMW6f9PJFG
sLsTfp90h5QKRvce5mNo/Yum3tZpS9go2fkybB2xFms5At7Xfwwtc5ypBjcvbV+BEqKazbASM26N
wlbwaAC7K9hK/TtLqkcWGAVeAhei2VKqxXs4TdR7ZgQRSuLFixz+oPCxXHzatQz0T5f6A5749T8A
w86DokAR0YAbv1jmpsfV98JQcpCaWC+/KmHhiruFI6MPFrbXsiJSmj6N/6c5CDeNBgefIJwmLS7w
afTjptvnvML5QqnNGN8ovCEjnDcSHq8CpeA28K8GnIvQVyv1leDh60EWyvbBbTYGcjEyuWWH8MN1
utXD7LmGHPgASQ3Jqmm2LOLuRvgyKRPy8nl7bEulbis+W73MXiFCrzEAz71/MpmICA4/Cf7XJ/U+
Nh0/rXrA3mf8wyDUFKlzcfWvUX2dFrFONQ/p3xHOeNNiNdeMK+REHPSWQqmFUKMBlcLYRhmmZJcC
vq6sMG2iXnrcfg2/GCnum8pqZEjeKc+MevU4pIHpRAjPIQBLbGHcPou0opDHvWBCInwH8QKlhq7b
FlcJ0ivuq1QUrRlFEMC9BbosA9SEWwdsFXbW8TD3O+7HUUEEcP8ZwsxfUldY7aymXeJXyVRHT/Ft
WnCw6iYjAvWCznM7gAFruS7nXx45kTk5LFVJac/4l0thCSeGcSMSGWNR99eShY2d8tD2mDn5UGyG
XJxMM3+ehI34aN8ztcHcZjgqkFDOHcZK9T0AcMuiUP4pdhADsM++ui1AmK741LXfxBI9fbUci4d7
gdHcxKZOjrC3jt+XNIt94luLAp1E7OA0Nb4ak/b/q9piUJvaUqTp47bzinGMlTgXBgtjYjZ34Q8e
oG0L3R9o7JX7yyoGxMG4VoqU3l3k0iPGO2Au+XunoNScVxO60q95vaFUo1IyqDBAFQiXgzNhhApr
53Wm6DjR9pve6RVKZueDwGb2poUYDO/GrGoPsUG8hYFkzzrc6uoqmBswgDBqVMJZIC8HkyKFSOtg
an60oEp5qGi6nyZd2eazF8XuP4c4oW2uDm0G4D2LpQRA2PnimHziFYJKcVeeG+04bv4bd22dEYEp
tqcjZr+/BgxUJkmyOZ8k1YTtcrDgaqvf+dEFRd5pmtHTqfxKq8gvl/WWdytL+0vU6RYT3/dP1NTp
GS3zq7Tj1Yr0bMBRKhc4n5ISqJ72cTIJ/q4Yq13r4Ge3KvsPQI/FcFEbjH5csHerNijMUciuTeN/
WSvlB1viTJY/F4+jm+mC4cNF5iKiOE9nNchS+sWybHTW3GW9HTPpiSd0fAru2SWpAIr1xNchPY5E
ufGiGue36sSdsTmP3WP5NOOpvnFrE/Vg85y86OFprnwUtB7qDHuImFAeC+4p2vLM/RsC+9KMeb6B
u8ZHl2bsY3Vgr6dYZJwZJk8WJtFNAYroR9UUST+yT3bOgIqP7X4mMzUwczs67X++muQ3AgLvRwXI
cM6plYnfMH4iafqbHhBQBDN5wQV4BEULLDTS1ABv9W87RkAQO2Jg9BijMbAEjWPlgr7PvIaxfifK
jzFRnJfB7VkgQ4XDIceWgEkpt4erm3333bGjcQTI15rfa1Wu9QP/1eojvQCmfocotZOsPBeuRm9m
WspB1RE5cRr7DSmkK81r3MW5niI5s5O40ZGIUG4bfxy+oz5wyxNasXPVZQU1AhER1940CyjJnJKs
kRckUoUWX5DGmn7PuwWffnbJR53eghwJ1pRqIa2QMgjxyB6UbBQBoKhKW2p7viwe9H/6HMTirSgQ
ibgJO++S9ZLZmaSWWznp1BLWZ53pVFwk1YOx141zxpt2W/bI1O84IKsYA0+77e34nrUGA65oBOzA
+uzddcXNVOtoymqQ2nblb2HI6V6GaPyuFMdkbX1CFeNLfVDTxR2GmX9a2nzLttZJqhnWluQBBMot
QwV4ystxfhmoyM9HFgyGqLr5f5NzHgjIWxKJoilHLzJ5AB4bKKxHrGKcB1h4fxq1o4LlMseF11SA
H2RUZ87OSev6Di5jIwc1eDo18+rso8CJMCR6dNC/n3bDtqdp919NNQxIWSbDTWMOb3XD3TuzMfeb
PSB6tXDK+PjWRryAKRChk+92p9knAX4HIRrMsljXK4NJaSYlK0QWzu4DyY8NBYg/K4afReyUd4vX
kjEgMg8EWeaQGTUkrRDyGnSx9iOPFd0wMoE1acUE9haKrS+l+KBEHdEpOvdP62q1/iMgP2Z7IACy
4CbYlcqWm2Bz4WfmUZw5xQmb/DeOAJYlHil1izzmiUysIfJoaIGN5k7EamvOmsQwfuOM/pGuTEaS
rp19AQxCPQq6KjOQcorUbv2JTAnPEyJCguHtW3k3jUKBK/lVeYydJZs606nzcUPRN5nfW0V7Be/T
YuYedl3IfAY4iLM5HpLhWK2strb4IrXpXYLlxzcW5pYAmOsC4nEC6rH0WjYmIbmCLU6QvulhLCuM
nPpjtN/H8uKfX4dTuaTpbEcqKF6OTdaHcOEFNERHH6dLyJHH5gf92cqx6DXLsu0Ym6nNFeTTWqhp
dGh6CfXAWBLCC5YKNrMLHFl6tNuj9C69fAx/KrGdTkeWgbPkOxFIY7XGcHXcscJ1eKX5k942wKA2
SHk31WYrL6eACxwUeorKcX8GDbXW1NMKh/K5iLSAovkrCJKA1x6aPj6uJoRur5OvIEV0Pk0zdakc
O1NgQrW+3N6MlMroHK14SWZskX8XQY6cAR9lhWKRcosFTPLjyUjgxltZ5X2so9vqkwmo4Gob6AsW
fYpXcdxumycve6kDDmN03t/og0XZrIE4I6+gBskeZkYnrVbj4ShlubDPpg89JFmDJNXXPkbqZsnb
EBu7EYwV7VuD0eHj+aakYOSb7S+WW6uvevRqbO8hbgqVL6w6T+ydlnS32py/72oIqk6wIC9HPB4b
LhKcLAfa/KxMLHendrfYkeqOy9HS5vBmo6c/bs69lKmi1WJalik4OCYmPDm1puYpnXMe0fn3HkcO
KgATek4cLeveifFwnfdw1ZWE4w1PgE8HhfVRxUwjjt3TXIvJFUyGI2KB+DOadVzOhfcSJekJNgJa
a6xrXbs97/rRT2JOLF/DXkDbTCwBGon8U701cVQb0MGc9C/SK5roemL972M4xBm2gLxiTLx11BXD
ZKnlUVZGSXRnF0RBlRhN845rGUOUAGsZO+kWael27lsq4uTynb6lsiuZuxI+7EsYJINawn7MkxIl
DovHg63In7BdRGNVnQgPi/HelL0KnEVKe1Iu+aVwXUtNpvge3m22d/0oTbUNuOqFlxjIFLdqkYPY
NAzuY/z8rEAnyqhyuKiVo/GqqdEPUe87JTuKBeIqNw/etcNZvoXHDoDOewgcvKa4OvJCpG1B0mFl
A8AWbG7mIdIwjgPVocuHxjDP+DXZwIoZ8E7Gt3V4XQvfKk4OEYgHUEgHLrfbMR+wgeiHpvWLMTB8
C6CKC2ZTavELcaN5d/pLXmhuJ0D9pT4QO8D0IQitFCZeA+Y8vU7KbDdNSG7R6pj1YvAPzN0mFaRG
/1KN6wBwcz8SGr+OVBfvEyOnp3C5bUp8U36EFHa0OiyIwmUZqd5DAv8qbqZG47Atnil4L+jA9eqb
3MZd/XyciKZhShEi7iV/M95t2/1y7Ck1sxgDSzlq5jf0UEEWB2XTb8AsyujylMORTttLR5s9Bwmh
chx4iN1zY9fyGG74UPSQuRgsl8DWrwR6cMNLWJXQoWXyOqti1HNSNbJiMki75X4jIQ1ECz27FzA2
V/AyUHCoae/WPk1txy+N2pZViRlUrSelqauiGVTdLMgNYFOwCQLzW4sfZUU251Ud6NDvMmD5m3Tx
ZrQJE6VzQA2VEUOmMrCHbdbSpWuOrj5k1JPVUgwhRWbwYqRHWL85jABvqpyKatSsIWIOSDzjJuyB
s7yEhn8UuzVvfyY2+lCbOdLRUziQzNnybijTkgjzAljfvM3YbJsRHnzCC7nLBbKjT0s5nzXHZQxl
ZbNzQ2PpMgFo0uGBJEWSpwanR+Mg97IY7tegU0nOgMdkvRYnOP1e9WhvWs0Dhw7zquKX79C9pTYI
msZTMVsFG8ESjp0bf7nGsZ8L/I2eUVNv6sEcxJui4/FqaHM8BIMyHNUrTUN+YK5zdlV4wyrJaJCd
2/XP256XyZeXxgOAU0CkiySWU2QcQfFgdzqAwLnFLNT3rQWoF9lNyukp+i5fqx38ztWiA2LnAGg1
vhcmY6HaGv0xxa1gfsW/w+UWxrcjOjap3ko8oRBf0D37f+FwXDfpVFtpydGXrkITJRoZi//XEOEX
3lYMyiRVm/Wep51ifeRsORgZTtxWPeLErn29PAwPLjmTuJG7YkN8SfaNDGaNZbg6a5XIQclWWrvU
VJ5qAZK5R8OJqHTGcSIEigiWjyacUxf8xN2gteicmUFl22+Sja2NmSfpVS1ZDpEtUneEExXp3MQ0
N96nA9o58HsBNzi4k7oRSmLguUyUyFTtjT5CM2mSp9wgXqe+lP6tuNa1s6IVc3ZsKpccOF6zNkWC
lc5TlHzThY/sg8BCPmyiAL9bJYazbPMaqSYQTy8mcSAKoVOIq/GQUerJNlgMwpjvS9bhMz6e06ZN
zvkHGLYAzQ96iwwtgNxaBWwnsxw5sSsYvz27n0vgz7rDmKHKZnvbx2iRnNZVPIQ5uawQP6YWiK1I
gbzXM1H3ecbLaP8OLLvWliWev6K6D6UM9DDGad+5C9gbrNQruWld7vxAv8SFfmobiQr7rue1EpgC
zYwYpJqS9qTIdrLCGd7+ABlZUlmz/lsgot2BuPaqQE2S7WXiWOqosbM+zHYCJW1ALAgkfmZcIogZ
aotiwxkiAu8+H6uYad06BRgtp1pgxTBmMDZN+2fW/U2NhC8XWz1bjsnh9PKwEk9Z1Tt3oMgVbheP
ApCe6JJGlGLK5uBuNf2AJQy7jBYyE2fwoP8Hyd2HShJbeZJRN5PMpOzhm5swt3JDyef4tfPmHdGp
3SKoi5i0lMRWikefo/zeFFLxk6Gq2SQwiuDFDRygbwteORTVFjW3VtRz+KQ5BmVmJUeCo1L1QsHh
3922gn3N1fXMCRMmVpf7XJJu16isJRXjD8NyM/q3V/H8j+gt8HSGNXbR5YRrhLjw9BLJGLwTMAj0
KxXdSN1R9CSuNq1fE9Y7jM/M00iA2CWmVhlhMyfw/Rj+Hhd4nAjK0tS0NH7wRCFn43yGcFdgcPrH
MVcoh1C4siCsxbwqnYfocjTTkep0OY+eWMUyNp5v8LJLAMpoaSL7SISAENU1ikzDoCcOzDQYnwXq
eN4IF87FhKoi+2Hcgmg4WI5lJmYqcIZ0RjCBxjfIBLdL/aFPL7EHZI6QdUZUSjsCcjREclbWtUz3
zzuHCreeT0wil6HnslOWLr9rvlUwKp3KlG3PT+Lpc00nuW37bE+zMcYaQ5idUGGgNJ2rzpOCTzid
LjeX2ckjqej6nczdzCdx3G6+pbq6Y/0CZoywBYEMN+bq1dyc+WI+wRuu7mCLmptKBg8A7cUN7fCJ
PIWjIHNFyn2veSIkdr3qSDbEuGCdmiaWSo4gH6d/zX1X1UVg3yhhytkWybz5o89GCilxI2tONaYO
3DMwd/QcUwBPJH5Ipn1qXvVR4Ce0SMBZjdWLYYyrNp7tu9hJVv+JAP5LkmBHNFTM73jazFUtn/h8
nOkt2lsFVW0iDQYyA9wkiaRNpLGy6WxsbbNQJscewtSBAvnxWZ4ms+c+OABarCZYN6U8kXyE4XAs
haNGY7VA6h36QNEOnhxjNNQvvj0fmDUNnNdzm3UjxyWmwgSNLqPrNzW0PwQORjekEpnQcIhcSBRN
IoI1r/aptyzvLXyMcKto/IX+orHVbYqqHdDTK2iRYgKgYmhN/IMKOQdoqkPa5lewdXyC0ofyQugB
iQQkqdXq8Ud2j3Ooca3xQGpJhiTLDhpbw1H3xQF+7KONJuue6CwCmRvoQABDcV00JOPsTpY9RKYY
MV5Y5wp1qHxWR7rVBIT4Quja1ryr+eCet124AG5G0C0Qu+A+EFfOL2eDaV6GEALHy18aMIe9DnBk
mfICIe/Qlo+F3RuOePWLYWjZ5TD+L8x93YDsvt4uPOWeIR/zSTeTswSfO7CIZMWd1HpFpgnXuL6A
5KnslSWjq1FuPp4Qt/OuG1wc2T/2dN11+1wO9v0+Ey7uK5jWVN/+rZLvoFnvfCHhKZ4p052W31xg
Fg/SK85g54ehvgqe79VYw2stkizRBEQC8mvTCdepmJ2BcNzAT+nbGdS2T3wQz1R7gre+jiFOHLbM
2EgQS9aZGxrcUO+D+f00vVJ3Oz+7lZxYVa2HihA7cG93RwFZ8YJ5NwfZFTkKQYRT8gxLbaSbY01L
1O+EdYqJj2EUuitCNoEv9dyo5Ue6X69+9L7bBzSThJPTuyuB9aDuHIJ5CF4NeDcuhA2kmXlDh8o/
2z/b9Hlg2A3ZDYtLSo8YYvvhJj9TjU/W9zvtkNz9MADQph5UxwBMSQs+1YhAt1tj4/zS6mevNdDV
FizInIc+O13bLDwyduhJZam5v13RMNFIzj/ZUyxOx+KsvPLY2qJZ4zu/P4mN7m6paxhMiS94+vOR
EO/wvg7Psqy2M/vNjlty3poFyUoeTP0iPiLeEYdgaN7mh61MAgvxUqops4FqtyBdKg6d4Sh36B0o
N0wOGJCYlh5EPzjgsxOi/e6lUR8xt0eBX5lhHV9DqFjbHHZ1f4VqEuFWtfwSBT73t8i5f/eF+JUD
B5Za2CMmk88rv/g643mZLBZZr/Zx4Z7ECCH7Zp+H3sxhlbCCYpvVXrRJr+iYy/kahVxx3mzQHV4X
TWrJW99X5ZRyqDGRPN3POIKWWt8MTcmaFsujUhCLe4cns6AwStWWcu7aH/DOfAdElDcYD6i0UAhc
IIrSXsPweFNieUdq/KgmlLDrmMSLe5YE4UhiN2EtD1N5fR+Hn8uyBzTCoYIB2DcfmDoONcq4+PA4
5d4paXvUtJ/ugucm2zAD/XvdfqTYbeolswbxeEJocIRcja0qqzHngENenKjutc2b1q9/KzhYrsdU
EToNfj6XcIxnORffZ+DNk5oHttzuKxCEFpsTgHIEnYSzJ9UNPM7sRdw+4X2eIP7LsAwVpQd7cDk1
NA1j3lgNvDhrs5b1lTq6zUshTfFnPcVI3WuWP2MJM8oeJfv5ZamPzr3nQ2XKO8KJ1WYZD0aTW2YD
sQx8E3kEIRlM2KjVsIUdxQYI93u8zcq8pI5xnb+YVyVCg6Ff9e3ED9l6hG+bfnQvcrGdo0OBnO43
5/YER8EYPhid6/o5wkNQEnKyMcaSKRbOsKZoLL0v5/EvGYP3UFb52zUpzVOFH/uAHZJCO0WPD6gm
A639LCAZv80b/II6aabUKX06qfoei29X2/eqKNRDt1AXDMKo6yZ9Acu3yu6wq8s72xNV0qIOAw5z
7gN6N/Lcv9qca2WnT8Qk6dLa9YhR2HYqZ6gMgJur9GeGCp8akFYg+nBwHnGQOAvMiPdq3Pzk9j/E
hIx55b2TO+52mYAOCms0y2ckxlLNf7Bvn8VEmI3aDlPQB5+8eC0kyVjqUSsEDkYadpBV0wnofjyM
bmIFs78JaRS4l6knjuAhmFG0H2NCxdn3x7nWIvE0eVGIVEh5ozKmqDdU7+etjadVCDGrt/E2eZJb
UwUZ4asoh8WlYRIM0KPC9o59FLMBhxpVb3awNxekFH9KFEzTYqD69Aedc5kDachIMU2lrOd8BoOu
k0etyg9RkFfMndGdVsaGHYeEB7ThZbi2kzY8aUtlmkqkwn0yFL+exfhHVt35IPtu+g7uLCQeUIPt
xkzpsR9ezg7PmWLdQtP4EwsONBfbjMGyQQfqFh5KSZE/dpWg5nXdVN3YVb+R4QszxVDUyJ9AOF29
yHuKxrje2CScN8SBi8s69NMEvdC2U3mG63lLsyX0w31rCWdAOQJ26IaW6DsyR1NdJywNzHh14fqh
cjaPmrUldOzvCTQ5cXmOd6b4yxqS3WsK2qhNcX3TVL6Wjw+I+eRlsA0xvhfj3pAWwnbVAbcPmc4m
EVoNS+m9Y+dc/jgaygSjXNwyBh6odtwGIzuQDAHqzQL50PNel2aGkrMdkDrfe004t9VIJuN9PZIb
HFuuZv7xUmf48JX/MduJfuML4aLACSkkPZAi3eslEIyfT1Unepz4Qpo/IKCshM7vrIBir16IWgSH
khOLKZumteoj6NJDmeZ/fQtArG+ACT93RuX8Mh93s7syqkAakhF5uwyGZI+SujrZRX8W7DFj99SE
yp6IdzkJ/MZFT2Q+pKZI3Ag64koQtSo+dijh7LnfRDa9wDYGmLfnpCwwYaucuwP56dVgpaW1dVLj
bunngSS9vdzSn/EPijL9K4N5ZNmK1i7vflXc/b84aWqbYOYi/P7MD5KR/zPE+Ra88SzXVCyMB/XX
SqrITIyMy2/Yvir2Q01MaEEMvvYHIcYw4Hwdo2B5weO8wsJNgF0ofQgXnAe74Yi4y9aRCMA88kRg
VuwLsaIT52HvdsUetwvXMsZ96LAg40dXbjPNDYkBWXTQ5aQJArMXrxtdW6gkj8p8w4NE2gc11Fnx
WKtva4NAYleCb9OjneVfuo5ZkCMoJCNGxq/FcN9lHh0mywCPneBqal3rBR0ZoYa0f0cGnXiYa0E1
n0DI4LfI/n2ZAs6SlFjktwbeXJ61PGcH9OyjMgXnDlP9pUuWTCmIx086/VPfZS5lKBQ46S+ReMZ8
t6mZL2LkRd9vSPlUtkVEXeL2RKuM6r4zlSxJXWngfUEB+msh48yiOuCTv2Mqvn4xZPaE5D0M5JaZ
RXvoOjT6ebqrkpz+WNVp+qKzoBVid+zStjueIXBLi9/CIgO1del5iJYMf/VuJOQB+RwP1uCdK5px
2p0N1IkYspS7Zs0IVqp5bsuxb0HOQORgpxLxoe1m5eSu7hc8Qoocoj251rRYXxhMv3dlxWzG37eo
hOkAbBPjBeib551mjAylhC/dyFgSksCm5YlZQp12++Oi2pbJSVumQFRzeIkoKhqF9rixXaTXlxDv
Z7/hh/UDsMyDhTG8PMnuRFg78f9JiB2KxWe9BqHqh9b8vuQk58RlFoc2hT2MaolunKoOWafDBT4F
9rt0O2iZeJNfSDLJt8tw8og92yvNDtXpZhgcwTn2yPit2cs2SP4XWN7gYtKcOsVHske3hac4N/tV
1dkgrb1H4IfV0KLErHqvJKA1AYhF3MBw01wC6cgIr/3pEC7E2F2y6d4CxSIJdIxGWls+AZfDTKq5
u3RvCfOAA6uWcQmFb3nnYGn378W5JgqcNMSJxJfl/blCYHNz3m9sCkkPMHjfz1U+YQf30XIOrKvC
rvc0ZP7C+6Xwe9ET5+EYc5XHwsGhPFMXIycFrIGEUZ/iTVxTDlNGCNNLEkD3iw53qxUNVmAeaNBs
OF4bEEIGlrcROgUvrwG48E1T0PnA8VcvflATB+O5hfQzc+EuzuONoRZy+dXqcp96ldPaP5kCNPWJ
a162JFK0+4yPTysi//SubZ5bZheg78kBIDd31v0PQWj+jmzColepoM/kNCwVeH6SKPPCfqTaW2zz
65nu461LqDXL/kEG8Vd6A2pCWOkwAVpXjoosuWppatsCdS/lYFcwjtGLoOoRfX6QQ7UiB1LGhHTd
aztIKjYPSAJoEskWUnFrZBFKyV9zeNRyjkbLAkHXsHLZheznOp31IbuFPaTJRyViUejZOevsAlu0
ZIXqO9WLlZKP6n9CMEjS8ertZ3l9qJHJNFiW8RmeL+h3ZNjX20ViZcmXpdb8cnp8DTKwQOFf5+VK
5An8OCW26nB3qmRHWTJmeCj351uCwVkjmQxZs1Agu2kBds4b1hQ/jylNxVM4PdF/6BakcN5xi0pG
rk6+2wiVYzj8IjqcbnIxY/9BAfJ/LJpC7y3J5skavUYXisHFQIwLfIikH67fkItYigmJwIp460/Y
bLfKikQmtyMkSXHbbQAGLSnBooOoNJB/faY4g+Od3aug/5RxhOyf/U9oe7dsmEqTB1SXXLS1b1Co
POk0CmCxlJZQdEmOMu8f2dJcvJl36eEEcSTpVFKcQE6nBfJunyzUQ3VMVNdHIYxvJ4HS7IvHuSQG
LYX2mJVLcO1RYEOtuEUhA9NXZ4t48rZD36e6AQYDB90CXwqXRN5SPdKhtZzVey5glyIDLQrjfo2k
W7sbKTYYXLRTQiC7+2o+j2A4PTERl7Pf0hKZ+cheWu2QWP5aNCShbrgRxcpPB/Ky1oKxwrS+0+3s
q6uXRF+O1sbLCfDTE87ETzGWfoyeJd8inqfIYbxOns9OlZ4qdIfEQiT/1XzAbkncaBhsSW5yxwQu
kS4zBmbWGO5hk8yXa9EnGtCvQWdQJwOXwCGNDjiFd8h8btMBCoo0N2Zw1oa36guEDFP1/p09VBqX
IELnOgii5r2PmCbfmpGeaYpfgpAOftL/J98BeCSzDNNrPAMsbwf1l0QlIawh/p9oDSa9eqoH1ROK
2Bvdza2Vlv4ffnSnr21HRukWNikKYXzJu+61B+967FkC25b03qi/fwE1BaP6ypM29cAMf4kr1CVi
n1Dtyz8nRfE6AuWdvlh4fhTabdfnf17Iy4QJ5uGTKDU/0Aof0WPFh1GufwG8AQrv4bAtvUXrY4PQ
QzfNxXyT5xAaxNwMPnOv7dcE4TZ0UWuCEgSv3dcBR5jlwcd1vSU133H7BcC0D4q+V5rkq9g+Go+6
cTXeFLIle4Q8hfBzfQy01j2VSEB9afOXUV10D6WyUM6fhRfDOTqj6eNxPVpQWpdwNFrLg/EXpcsQ
W6uKDxJMAQEZXPtfhV5SS9q7VxzSRuVQ1D6lXzjQBvPmMJRC4Ailz4pgC9CxsWe2Hvs729kSy3ev
eyDxJlrfklB78J57FL5ZXq493sHnxu9LOde4ys3l9p6U8P8PzHVPIncmHNw/DyICi1FlBRMTr2lw
w6yW7d6dGr/oyK+1zNeiLwumBecRDwiPxsBZ9yYdPOszfsvpuIiuZQCx1fPEu9atLxgdUhctIdxK
CpJInyvpQqiLUmsas6qZmtxb6xHvCl8yZRdwMpMbQE/cyUAc6tDkLcf8MEUF/WqbJyEo1A3/9/tu
SATKrSzikva+DMbjBabvAbV/KXYrv9Ol3lWALjjf1mgSq+naaoo6a23ixk9nXg3MxvBMIq0nxX5w
/ZKkj9ZSkRVydZCka2WTUWC18uKDaZbROTK2UJMJ7/8A3I1UR/ZdHER0z1iTDawHjwgEiyhZYGjM
+dCnJSqZS0yA8uZjkhxItYNGHkyNXwRgaPgJeQz/N7hZVehbNGq4nQuV4+o5v/q0c8r69K6IXqWP
k6jb4mIkBw6qrUF5r/Ngj6WhGNcddKv4+mHTsUaPeb4oaIUha6fjZstMVDoBti0n+502OEPMLqSP
LUfJHK0Fi1CeEzznglMaJGvMsxYhVbdeS69v/qhy3kQ45V6202EEDuA2jhyXfg0vuZvxVKNH9vYV
AH18dko1arBTPeeKJj4uwnwV0lW57TwajGypXfHRlw01BMCz3wwWLCT4V4TBTIioyfuUagaz1+la
A3rkKV1bJbCIy0Y0azs5fK4k0qyBlOZ9TGgikl4PbxNvEeEloJJnWvWxLIS9gyWb8Nh8ken9aNIs
HU1ECPi2PhwPyBCRz1syGOtNNsk5H7TGPzK5xpn5ucKHi/55TF7N3c+4iJGe8D+vUn7jRheaRJDH
LShr5UcXnPo407tsJv8LH5Rxz0b1U3bwzb8RBvXR9LnIQZmAMEqaFN0F3dO1lsJSbuigQPLUTL53
sOYeCUbkoCXwXtkj3dXjfsydmhAkDZl2m/CuaF28Lpry2+LizqhcmYobEZg18khpNDDbQkIDaDW7
GyLonAAYNWGgfbErkswlLns4IFaIF0LZWexMWgKw1u9lMIJ8MavaNC1R7PCVWByjMCwWibeALNDL
o4KTdPMbFFY6WkpgKLB3ZYheik6P75jr2OQGZJxAY5Pw+X0dB6QOuNpDCx5jGny1K+QJxMGonOjq
fNDD3jrV7NC7L4G+Lmtuic3L9P1kzCjHA7g9G5y3bGO0gDlsdqVNbA5MoyzAD5vZNYP3KlgDsGf7
1msS9WwqvGSnqoJpgXUHMLowIgO2AGQxhK+E/pR1ipafjgB/G0Afwns012tYlkYvPOJy22jOgSu8
nLeVAdfJlgxlAcFoBQ3ZdtVwtV5HODglWQ2UAanLvSVKhhflwTmOR+lfN6QnkDHs62RX6dMax7Zy
3ouE8bMvTej3OCUbmQcpO9RGeiUov3roLF4ZRNzUHdu+lRYSzgCoob98OFnBPgLaZDKG/FqxMJu+
rx7Zx8v++y4s9slfCAlYKq8LnyVJbvOBucl3znW0lWU7cywaAMeLax0hGM0TW5Nwfvtk2eVDEiEl
hO7XyVEK+dB8r8VWaR+AfjqNpcMYWzRRcc8o2AXRgmRR11D0MZ2Wa5QIkSFpSPZzU0B8QfK2uLNU
QzFl2Piz3ajt5ciZKizMrhcOObXt3AUbENutLOQgRxdx9COaaPOww/kqKe283Smq8j/hFmo/oSCA
IEQm1jMaV7BAKm5CD5l0P3rHx5sFbLp3/jB21ldPXbHYjinUspAFL962ff3cTYk2/71REtL/QDvN
LTagW7G41HZ2xmROTZa1ardBYQ/7R+PyyEwrUUzg/AKSbjEXv9tnc5QHKqvuHmjxMan0q5+pTjlP
aK+6WKUQQ+gn7zbsOIIJN+eP/ag/SVZ0p5qtCJishLp9wrDu71ByAa8xlkdGwJje9PdlgLlbRn3e
pKZtQetLA/+eHfPZllfWGVGP34+rGYYt3HriZnW15Lp8xi/rKgPLXwglbNg6FITEpFaJaOOi7GBN
lhmLhICp7nrySdk3BJ2pcQyv2aXWYGBtbzUmK+usoT+UmUoqPGsG7II3F56/EMk+CbOQVA4hnZcX
CmnRuoRQdsy9MT4cTV3f6DAjTntAvwwEkDeA5YVrzfgH8uGuxUGm0IO5zPUY0c4h8ShlYa25qiAr
YWcX7lCGe3ooZ6udo335ncChZLk/OjpBncji8DNAiMKkocIU1BWN6+Z4fWJodQazg11+opPoFEUs
OEUh0Dcmd4zSCBINlSFLOmE3JrQC7H6JFvsP5vyaXcwcvppayACvYw6SG3qsZhIe/cBTCywlXwfb
aAsTxEs29aNfTDoQJlwHqX+x6dHZ5i5ysBBsYczCdkFNU0A6zoI63/+Ty8z8lba8CNXPHATW+hL+
AOkzk29gCm6p2InQOQB0p/Vlse4Z88b0w6PUM4JzMKPgXEY8hdGb6sGp21R6gmtaHvsawdNX+Iv7
t4k7mf9RKUqSrQQuP+t+D0qoWU7KJX31nXUxsmMhvcMWQ5PkEyFu3HjngzunfRQK/R768Jq7nkAK
Wc9912Yu1BGtl87h2yVGw8OWpk3B/WsqInHXC10UOgfk51WuyKXmnyi7idpXwCngGwFWHxrow9Hu
2Tvpj5Qj7fLHseDl9qkUYz4OzFKtQ+P5C9GnraorshVAyv9tdSAJP1v8uLcvGCLod45leqkQFcW1
eBjdKqW2I4zkWumZ3xG+W2n+lHJK03rR5YiE+xNn2sYKgBp5zyBpPxBOvAW5mwz+qeP0dOevB0Zl
HuCruCq0Nmu6bOn5n9IIz4WOFJIKz8g+ALSOxJjOCgB4ef9tD0wwRVtxn5uolifzA1f6zehnyvV1
M4QuHJJV5wbF3+S6Cr9+nWtpM9xxyTO9C4/jbTgGJZRX87QtCE+ZP2XG4pSmN7I62+jYAZGpZwg7
L6bt8iytPIoQHY5q/2yRl0iXOMaO6wrW9bHwQERttlMvKN8NiCC1QXURpCKYqZf4Xmg8FmRHw4Wq
OZw/hJ8whUMkn7bTrRl54bUj98L4KX67fMcLfHOHIPBucGU5fqgzntIrDSw5jLOkVdoRRfNLpt4p
BXn9AqDtdMCOOVhpJIRMgfF+yIOKpEnKezuy33Qk8EXNshto2clPagt+ZCsB72k+IzPaiI029PXT
a0u7rBFA8jycHyj2pxdtyHSVkvcWfzwT0SvA+9F3b22goaRFGf2xVHZMaMHfIa+lDL6ls0DB59M2
rvTovVLHvZaioUtzGiRQuMlUUq2D8h4AMSu5Qvr54fdz03g1uXI9GmvaGmpYhYsaopOD8C/A3hs+
ITLiUqba2sAdMZ4Hq90Ju1ip9QIWiuNziRCaUyPQzOcTdBXFmV6xfmAN6GO+GM6pSTy97ch4EMDS
rXwalyNDLAtFf4ilk30qeTdy/fLf+1LZTJeYHVdJaDDWGvpIpI26TT1WTUuEx4UpeAqLd7Q4X2mB
gQEFGePcLV2mF3K1IBPZm826tJCjVwDp7W1wOpg+9yJycKNS6c82ER3u28+3K9R1TKGHqNDqZKcF
JXGFUihfjAjGu/BmLie/3DDxF5qzLeRx/3p8B+CBxXO2eaGF6YjrflQRW9XxRKyDL0cGrvLN+fz2
NPqL0XMWmxYSyJSb3yWddSdOqgvkhgnVIgj+OaR/tj7m9B5drD2L4HMb0ZdF7d+rVX9cIvYB2Pgq
K5nJYsxaaRc7rZoNlgSTdTA++cn44P7l3Lj+fMQlHHU9AN3MH2olcX8VDJSYYNJnzMmSlL/ktDWi
Pa4nk3RLrwwXacJPsmQPTKxyUGkcmNM5fYyEjMen9DjOdgiin3JxNJLb54FUP8v/yjiSdwWxUqsV
SwSTmGn96aR1249zVF6i33tdDquXWM1zdi34EDqbEYxmPj4gnL8eVaT7EBjnq/27Q3rmjqKBeh+v
BQvtx+D2nHySzAh2txZMPuLaBhYBYgMlS/yZ7IvCo+tnCUrS9zze4+0flAXPg2wQH5M/6u3ixqwJ
SnO78XLH+OzY2nccLUvz2TyjoHicu7bQIZ56h3GusbjQPubYrQ6wNys4uLGAW6SP7Le3BPsPhwyK
CmFwcSY6S/KfaYMcZlbNOdIauKQQte9ZLSAiHCnfc2Opf48Xs+W/Vz2/ynyNqMJdjWSBXNGCsVSo
RMv7vmhHaxyVy4i7AhyFB3gXGVd5Aj91FkH+ZBXRu4DOP4eaNOxreJaB9QgQee92PuqTMaxu5BQv
q3oInT8wjRo9K7rQ0N0pfzfhr0caVb3/1+PVaWVsbeFRwQgat6vKujAhiMw1gPxlnzxQurBxwJRX
i4bwuVnr1aqBkNsAJohdyqc53y81o1R+94NiAbuJyf2sRraOhhCQE0cWPxPWpW054rDQN+pKoWiF
SmDJvP87Q03wZyUbS4dERfPIbWJPCB82Tstzv+txmUHH0koKT0L9BGZD5aL704d7TRnPeuujNLGD
LeeF83RzIdwZ4X6X2/rN4zufjxByJYcZsELMA/sBd8HsmlGe3BNxR5K0JUrTTwKSZkqMAO0B+Akj
k0EHRL/kKBFq3ECKL/usv1WI29krmWI6MFeRpjztDyiTgEGVg5SGxgIskAyCtrzEurM+6Md1xs6R
eE2fWLzd3i7cOj2R8cICkVGH/rvejKQ+acp8eqRY+rZZ6q728jkivyerbLQPnuD5FXWHumdzpl8D
3bPfMObQpk8yOuqWk+JoY+rAM3VIYcwItJnuMe6e+3/mSnE7gKIkVIUNYIUfhMk3GqRC3ZjiZgHN
GvGP1aJJnm9m9jPNTkXcr55M75F1jQkWod2kuDEWYm6A87v8HWhkYfaaJmdUrSm8eD5w6pUrKp1W
AifPzw3qeKsHsyYWtjjlDVws7kXal6XDULyWmqvUkyTrVqCkBzWS7iuBOzUXt1Fhxm4Rfd8eOI0p
tYbYN8GitZOYNDj03wggbc7RytaKNxwqtwaL7P21Ib3rPp3zEqcR6R8t7iZQTC7VNb93hyM8Jrfu
XPFxvAkfgcfbWcq36RoqBRp21jLpmbW0o41xzVk42fPsN0LeoWDwEuNiusZ7fvIpHZnOQG1Yd7Ho
D6jtvO9VAn6AqsWRrVP2pzpsO9mo+lvpYvYiU1i+42UUaLl7zE95ZRUsdwKLuXw47aEyr4mTUGs9
qwCd7nb8yfP3/iCBbBZEIpvJbvTm7PkA9/z/s0DA/OU4pOIpVCYTPeWUnBFChh0B2fO34zJvBkjy
J5l8XSjI4IdAEhSYFg/Zv0B2oBYV+O3NzrS7XsqI6GAP7Q0+3jl0gVKQF/vm9Bpilq6+ldziex6i
8Ns5EGHbwWFtToG5Y2ynW4jnQkXpcCz4SA0cO4QdWJ+kg3T5CpTAGpb1WCLsaitXwLi29FXV3JEx
3eBYR/BxZWnyc6kPt7jPYxi1D8DHjaX/0WDqFIlIDItX4NxUH04nEEbX4ZmWKQUGDzeaGS2d4NTU
S3us7u7QNwYmmqJnha4fqdmnanBqGOB21Wq6xvs5OCsctPtlJPlI9/x+7ig5UWQAbzNGdDqenCAK
Y1uycAHLbV/TET9NQNe0g0SWbre45C+zsQ7V/A5nuMPPb9xY8fm2NWqylGeJWuzocSy+qQY1uIsw
XTecq4cgnswT7SiuYM8VCmYrRrCkw++YbiSq3B7XfdSPHaq4Ms8MeERs6Az0+GggHosSTUr+bD0L
vntKUhgVAqqpwHEzwpESdlg66K1fXy3JbDRGYH8eYJr9PlRXao3DM8hZHfyEpDKf0cbicO024xv6
iJx+4RTkLnZQNrpWEC2aAxRR2YPwBl5WyCsAt2dvyCIZMdkskXZbmaQuyPGCFLWCpOwdSx0dy+uC
6q+aT1EZ1NDswbNxtIBlSz9RNUd7BR2n4QI0kfiXoH1E36oKaWha3HD2jFsaC2DtqloUb9P7HHrU
9DzetOU6Ol3VDkaAtzroKnR3nwAlvBNKVLtTbWd7rDJpImLkMo3ssWRvOT3ag1yUuCcA7lwx+3ap
44vGHB8zVD4c1USRUHJyX1vjL/UVI3yGLy7FT6P3mZeYCeciIdAMiPkG3AF8WyMiIqa+ObNkc4XA
WJsncmcQzyrvPPgEQM46DMS+fq/q/bEXhecDjtf7POA/cR3FStw9Xd5ybcoEKPzKRy2pH40IuHMa
lEBLvL7lJC20/LSEHghelxtBGlI3F1YNlEMG3MWJHkGrkHCcMZHgosNmvy06h+G+YvRoS/Cnjatp
woSq1ee+UJ1Lh+t79NSjJP6WJMyMT6mMFWzymoig6Gd0uOCTQuEdZYK4mlfE4U0466gI71epeipp
dRb+cXt8sYmJjZR0W6WR6wMXz1itccaAmSYVJFwCyX5OBo1po18IXrSynQZMfUqXD0svOq+yRfdK
RtFE/4atBvGV1AtajxowKj5fKbIz3Nh9PBkjw6MZkV1pvJ+sYjoTTSagC5HcP0FUSiNUZyEIgeQi
17xJB1TW18c5pJF1764d7ZPFRo205c6Kn//f7d9FlGkOJnwqC6ktS/b2hg6hv37JHh1k8Jw8/pPi
KqTyLf/stfwQW1ySERKdjw+zNUJRDHQlN6Oynb28EzNIsXCQRBzG2zMoFlQ6MxNayYUY7ll7rf7A
3r0p8Ni8TLg0k6nEu6O7VVH6pwe8RSdI7IDLgErKgEYK38K72v/v/IwkrfnVJgsMaAX5y2iWF98L
Oj0h1cy5xa1jy/pNtLNMGjkrnLIEQAn489zQlfOYxlo3tg8ZXh/uxlOMmxScftWJsLpAXHYz1FE/
mgccv0EYglC8alT5SIIcM3j7xy150V9orG7hH/EJ4v8kYn3xJBxjVgd273KJnJaV7qIDUcGEvOrf
cykkG0Kti/mtTvFPy/Dpwl+kAtqpQwxTVo5sYL3EKWyJF3/fTYnHuDdjHRS838D9Bk9FQG/bnXrn
JE75V9W1CRTK7sRFaYcQHoqVxmmaW0LAavtXXjREIr8c1u44tVXrQ/03Al8UHVoHTgkmbODcJUHg
M/8U3wv3XxzJEznbYjMLsdqq4+eBGElx5M/QS4IL/xRTnq0SyY57lIvvGkxz++a+SM0b/MdrIvgR
iMIxpZVsskLLGi/05HxpK3e3xRYxjW/m/G8WTZ8pKsgeQ3IIU/04UC6CLWfMaN3oFghsWN3ATI1q
wxfco+MIImbXGuxDHGPJMhHDZUspciBwvUd0kP+6uulPom05MIOQV+I4Cne8PwwrYvkq6YiG9Mdc
SAL8M55D7s6fgFEkbMpghmxbTPWii3sDqnVUQiuMyKzleyHCHNqrtbFsTtTAwPrlDrxHkhFLXfbe
10AhVXRoVe0lW6eaCFof/jAdBP+bXas4eUm6zYkPfbU03tgVNsfV4uPgUWl4LjAyE6qlUMI+tBHQ
oxXXtb6L+nvJVg3s5mi1uhdgX6pQ62tkcTgCV4PCtZ7Z+EYJGuBaN/lm5y3xXi8h+WOb3WD1tL4h
ffxu+sWpR37TSEBRixpeYBZMN68ygYOQbqNyOplzbPmsLzfpwsNbMLzAHyQMW4SD7nWzRigUEJY0
YVkllvTQsSdDXkvRXDq9VUcDSt8iJ3KQBrgS4/ytUs43VoX2LQr2VdVGgjXFBT9Tq9xAXWcLOfM4
H2HkW5YnKlzFMKW0O0YARjrk7ROVgUy7QUH2atvwMnN/f7Rpf/gjP6A3ZoeVF9t6FrDZ2XwQNWIH
Alb+uVf1xXMOnEqkCwcp3sWWie3aPWMfA76cDiJksEl0+BuhcQ0NTV5+UpH4giK/MUmEuMqxGHxL
HBmNn/DQixTb3rI130cNX7525yMWyYWLJqaw6XFiEdwdkD97Qt9Lu9weG5eOUDtKlln9oRuL21v3
YSyqDDgPK0163RfLt07XNIuhmCuRZe8rewM1/RjPM/hZ1hLqwje27crwwPuiLXNlDkkMywkOVgup
9rubingQSvR1wns7I5BvGGGV5TGW29umZKQE4TDt9EqBj+hrsfAS79cFNEnfxwsvlxnuvB+Wwgz4
mBpStr/oIiNCzk91oeebL6zpG8zd43r0enFwMFrKcvslvP37o9gFt6j/3xy1Y8aPmsVFvYg1NDzr
6+ZykdhncMTwjaJ8mywc4yQrHdV4T+skmmyT7jS6Js5zOE89aFj+M4lFMmZbOQ8iu99TzDP+y4PJ
ZHx3885Meskmvu05jwBILcvQ4PkpH6KVdjrDCml1PBA8IFppArG7JLqg6DcA+VxYJ0CvxVb5uS82
mKXeH4sqmAFDJ/pVPT9niv2MgEr2es2oPvfagnqnTcXpASKZlgLCGoyrZxI6aTktPaowTE5xbb37
d4Vp31Z29AnrHTOetyWoxLAu+riuyqd+9I1yMSpWUI5r66UU6Y6jj4F12Uk00O90bqOli0yzw3rJ
xRF1lCMsukJdD6XCyYtQ3YMVsiZzBu6Fb4N8q+uBe3Ja9+7cnf0cwHydXdhA8IMrHbLjI7755kgS
iFhpwygxVkJ6n6WyHS707HjFcsE/B3+34ky5uYO9X4DrHW3RKJcvNnytvHkphvTXRV5KjgBleOkZ
23CJ0bNhobwuFyWfElZvEzEgDYtlYO1YP52ll1o3KKnnN7JzYCk6TGb4/XV10Yo31pe8Qi8KG7qK
VbKzaCoBZbR/LWGIPPV5WKoYntYnsXiG0kPUGoXhHjeRupx4k01NztP6hQfyzU+hGDyqqcMqwnRU
1i5zaIZcAqfQlopfw+JvBv5/HMMkO7fpuhLTtPjNulcLnOqWhaYu6tsB74b3oJsffiAEOKIGLiZZ
b9QT+WuBnwyp4D0cG+fBu6SVcoJ2bZXxlCCMjih0S/wssAvQITYDkFBhqPuuGkgyiHdfax1VlsN9
6BAzYloUMwt5nhCFVxXy2qtH9ELxTnDe9ltV/5RJ825hWaHUAm2cN+6hnJ+0TD4PBn6kpPV+bSK9
iCipHNLjLF1EAruD9/uUvpxGPYMPea54BmCfDQYn3pGiqKCb890b/wBbv2CBMFrfiv240YFm3RrN
TDkMMkf3M78xWFGs/1onkPedxdNrWIWqFoQj2ci1Jwi11cGQbdo66JvnREOGsmkR/54aXqmTZB0R
ImFhKAq7hqd84y1mO9VzmriJ4cz1ueoDKTwS7KKudPJIU6xKtn7GWV6uBRGo3Q37ZWwcu5fdktgN
LpQI77av+YUlPK5dT6Oredj8fKWSK/p/+K32lWJSHuEB3GwpJidoxUR1Ks2yBjWJOOwTu/HNT68C
OdgeKNSgwbNbWYUvOXTHLwc5cGtETcb3uVQkL34zGKHVc3in1JuMCFouVTo/QB7UKa4Kwbm7O/wH
eE8N9bs3XFC3lvRePjKpnWgQpGJnBWjsbMGoexpSyDk9B/Fc+KDxZmfHikeSGJOxyX2/apVa1MwX
0HaaMAmYAAhxG1erD+8JiIeerhN1jUjyWCrZv23Yt/P8NByiG/E/q1R9+f2bNg7FpezFtdJejw/G
8VAauN7mhez37GVO03KZSsYoLX/bS902g9aiLY2DqZLrGBsT8gxEK41+wa7xwCimjeeUA6239/s/
6h3ncECrKW6vLZ6fpBMD7FFRrbqyFWMvvFhR0YSG+5st2ZhfqGkR6c88M+ChLpuc5VnrewzTAFsk
MxB9ffjtndrIIlfPrXsA9ofkzkxTpenxvwfK04HdXwFoax5Eq6CyIuFmd3uy05LHi9/Me13PFCT1
qSK5UB8wxd8DF2DumU1Cdqv0vXy3khabDCasiXKpgg5BZs1EIj8mFfbwzETw8LxVbOV7Qj/BUI2I
YR/0eDebCjCzqynHJ7viHVZfyNKyc5Kd+Bl68mqMhQrRWNpnZYDlWAyZM61KcwD3J/1jMmRtLcCY
H+DkZNQUuHFMInJ1bVZhBR9zYB3wldkSV0t1KhXMahVk4HmDdiLQaQgLKR2cBVZVqu40ujmgjtjG
+QS0dAFIvDnvSmao3WRNxGnLZCleuHuCxO+C+nWEnkSi6FXyL5rVjDymX5KjPRtZUzyP8aFvUDQ1
5mgaTEbXtO+Xdj4Zy2uB6ir4PVs4USinELPLADHQDvcw+NsDJuQ03cWA4KWwKHgZN4Mb5Fxa7wM3
2dR+ezhAkEZran0E7DCRBJP4lZVAdiXS6QHdLq0JUcjHSBw5CNbKfsN5UjUjSRfyHSsUZzV1tXqP
efncFNE2bbDtI30doxDFCkW17w0Y+sHvnhkusEVmhC4X+GyjKe6lF0bLRnIrs3MAjXuvWXq0YWjR
cmJBffXLT+TOesGsYIqYF7Q3+1Z9KM/NBpuWc/myxhBhwVS+REy0d+QBPJ8+5TJD+ob27PEtM2hh
VUvGAecb9ml7QO2RzeEc6TSlgZe656d0BEoPoQoIYKa05T1pPZVeQHOt0/QTG7YdXr/3AQKRDWBv
Dk9cLtF8MN2+EeMI2uQLj8G6gHrcRlaRPDQX6yExX+7Khd1WNqHt5OGBK3mKJcRiz+6iwRFFNiEv
TKJPuV8UvzhS4Ymo14B+pnvqatdBy6wQis6ow5SLZoYRAaE+nultID7uL3GrMGUyFEh938ggD7hn
0ifHzWcwxlI8mQ3wzylzMnbmTqmSqyUiwKIh4uxDrmbl8q5k5Wrycd5YDxIcqHjkXyt6KgJnwrTx
06LpHpw0Tng50UtjHMbpxL9ueBjDPFZDS7gyrZTo1Bd5JSKkXEAaUA+eYRP0Bm6oOo5bC+iiJC/q
ii6suKUAyEAG2XSHQhVi5pvEpXQMfEPoCh9KdavvXUy6/PKYEAIS9GBAligNqWHNXeMHCL8HPftR
4QMc18vYUCXJv12bPRf2McNgehBS/I8/QJaPBTa7NYWhoWnTMdOTTauoXFu3XRfkWvaBShMjwt27
aUSbxr6k8LCylEA0DBxbNJS4/jZtQcC7SUfSWlwaRJZdJe7Wc7ignVbf5cXsgED/9F1lzHW5tEEq
VIkb8hocv/XGbtHGepnBz2+pQhxvWztkejeZhwpG92Mt83JWW+roxhUAnCRQn2+33A4DWWvgSfCp
DENThr8fkmI/GEwUOEs7tY0QJ/mrESKNKbtxjDeqZA3hb+zUGMbfp9wwmmH2Q+syHaULXhIuJyJe
f0ZQxOeFXFnnwXaMtyfHCyhSyHa5VG5bX6O/szz50pkimTuibCCUMA4qb29HyR9OQ8ddXvxoqQCj
GP4qOgfGPQfdyhgJSbVae9x+4l4IJjWeWkPS+U3RXUJCY46SLwuV91UbD/Vk/CxbADkvNNtaglaZ
Xv+ZypQHV43vMEgGOhDMdv+Q7iWvVvnspi838e8+V58p5VBpBfNVye0uIHqhuIBqHcy+BUse3nDg
kLUjmd4l32ZV9uv2grX02Re/lzzDwEPgavB3NUOqtFXTiv07vpdOfzbQ6ZSqyfvOkupqVgUA0JCf
0ochAAWnRTX0DL68lov5YS41SMRDK8J9Rzf0VoweTioWLchyTLUR2L96krzlXkjySFylYg5ptA0i
j26ZmjUx2qMgRGvhEQgDXilUj2uRc9xddzFKGLlw+3TZS2x0LmZpSug5EcTOejI8Vad4jWmcStjA
9HKBVTKx5Uvk6qotExGNcfcVYf5QM0URE3NRVmc2md6JXKL0GiGns8CIncTISg5KC1+pfTo95AQ6
r9YUW7NOQWj5wl5DtiL8wnLR5PnGU2XLNtI6u+ibOI3izGKse1XMFMzjzaI29FzlSjy/TKtDz4EU
TJAa8K9+J1W4p3Zh7DksgMBUvCLsZWGcTQJXrDLpjIG4sED/0XL60LLHsqHkQXUKHjposuwGEi9V
p1i7C0A//NRVZJoNGsGcXh9tO77ZbibNldZgB58k56bg+h05ZGRm/9P2wul5xinXtKu80ElCc8sy
QuTxwc94vMi32zFY9I0CuOeZvAAKMBIizknNt8u6e+LCSEp4uqijxNGOtlGq7dT82PaJSD8/mVIJ
grkKqtyFVHnllx7KPGQ2axX2vRaOUgaeUkXZjup0lU0+AChVGgJ199076l2v7Bk8aonCcYWBqzlu
KTJENymKQuB8mQQ/Le5tXBt/MzSncIrz0AzLpOMY1+jukT1xpaHMdrOlKjDJU0+JSE8s+AhHkFx3
zgHd5LTjg+zc2KqeOuVLIDm2RGwcjNQFDDWjPF7XBsk+769HfjcjhKiw4acOPy2KZrJeBIfGTj9e
vfV8wfi08+vUSWMNBev13CGmfAzV2FQ53q0QD07VLB9taPMD8w7lAXQ7KikU8g3IqvBFk2Jk0vQr
QmB3t/bg8+zQZOZ6+4Vuck135UdRoZB3WvHLfGUzF/ffAMgG+VW60knBpNvyuF/vxxDmB1JQWjRl
i3ZMce5MoqQTXnuESrl76ccWggGhNM6w5SQsSLWgocr8P1Sq97XgXuPrpqO7JzqXSxBhuc6bx4T+
6LkTgTOW24zFisMmF43QG1oaZSOEbExw177k/UeLzcNkEzMc7mLmAhKRQ1YhupeWFsDCKnRStcT6
VStvA+RmJFe9CGicPi0ZaWQPVFXKc+F/zFT9wPdnRmN7LNwWJoCLg2q6JiqCuKHCA3uwgWv8pc0m
bp4XLe6IVU+/2zKq6BDk84lVQYlrvRfSCKzti2LiGPDqXPk/qO090MfCcYPdYzfjKWBKLGjfM/QU
wqGQSacyp+8sDEaRtaJiAWqh2PF3ahnS4G1j0nsrjEmcToqoG1lWEN41Rot25ngRU2I1/u5rbcYU
JfG+ztH+FfqGa72y/quLK1USOdLEX78syunSFW0qjfNQpd/UDyX2vczopzgJv12i9BNmRGuNrR63
RGJSwovsPNgh8Ve36eQKMjrSl+pJU0kOQsHZRZfYepwdONPvegb4+cfqj1rS4ubIttzzvZoviQki
KPZMHwRGaYnvr6AhdNUkZoGnkX3dJ1NmWuL7d1IQgTBdwJJ0mVocxjiiwrga5LLNBstZSd6vHMP8
poQYnOFLG9lUw++NF/xBUTAsTVXjN/0obTlxCb668q+f4Ma4ypgsUZ6cog1JpC/gvj/N+eQwng7S
+xeHTTbopxDYMWZjJWqouYjI56yloArbkEYYMDEt0PRR7ZpoRvkBIXVc4/hScKWMMT/4UnM0ZR6n
0sMIbmWGBsWwWHyDyPZIpKp3p9Y0O/6ogKXa2aRQrVlcSP4WxmuFnpTtPnA/h6Tv0oUpK5Qn2Wn1
XYXDQrwb5fc1j0+b+22dbCU3bi7XKvZ+kjR0dMKqSNRvw/Fr+Nmpl+nWPgDwiKw3ksENL8ovcT8m
IndU3inelDeksWQSPAEZjvAs2BYr63NhA+JNHE98p7quLaJueDUe94N6c9QKaBSAZf2o10qTYIwz
Ty1fB40CYIewDeuiXU6uP9Fski8vJ5kc/HpckSHI6uknInRl3ksWDzeMQjtpCDmnJOONLLNvXKk2
2csEZdM9Y+y6nhzre/CWv89eIqm6GYDosyhVl64sNwCHmeUJ8mUc2VRBQ9WJa3+6ooRrf0bdX7Dk
Yo/UyLRXFuFv4oaDA3eH7dWKPgJ7NCBLQDv8zUCdCbcisM/wXijGqhkVRshOkM9EBMAnWu+3GTSI
VUywSALf6nHUghMdlwZVLEEYprFC3g1E5grUQvvezkm68BS4D52n5d7IIFk3eGB0XXfiElIHXrae
uI+ROW6TjjPI41JEbt//6Lrne/fjSTczf/L/Fhn+Y7Zp4PxQKUFqkHsd4VCO8uukVvv+RKTx3Y3E
GG+lifXnl8b9hRa/kaSISZTEup8f3X6r3d8MX7W+kKJfmZrE2V5Vb3b+FKm74US8TISPiABCFa3C
5GXWRm2dW9oagZb6QEMF2Ru5UyPBDTMCOYikrqhYzvVNYRCR0W905T2bADqTVSvu8LT4xCX0zxGW
1lG6sdqXKD37QOrYoW/zcaVPdS5Kuw+TjEuLwvnba9qAzhfZ29ga9NqOvUg+5T9MBTGtgEi0MI08
6t9kk9ttKGIEtPebtN5hDMLokDyppHH+bsN8joX6AqfEUpGBjcsGMS4oI7s2Y0jtlqTP6Ao5fJP2
SZKOqmYL8LdGyk5B2idJAJaPcOGSYhgq7luJm0cp80VzSaCbbDUUA7pPUZGxa/ocgSweSqrYG8mL
ks52VPt0XZNwUsIDXCtOMKynJ0tHA+EmlXr9H/m7N8uGQCmTuPzZV4HkdQYdCPiNKqCOChJK0G3Z
0I6s1j/5uCVjI7ve0YGdJrpH1KJr4+S9iTwUvBk8XNQmbR8rqqRM6rGdwpdzqSWlQdvVf71QZuxi
VmeLwj4tM/l0DwDN/+A0k5JovNYAeYdEEyf0BruCROU5u01RXZ6TaMN9S7IBdRqFwaiHBs86WLXL
WSed9L2vtPz9pmMgWKej+1s64nXmoqqlozugmhukPtX20e//ZLEubPzSccn1yV6ePN8kbg5wETCZ
SNZARgFazT/Fo/MhKzY6vT/EeGXuYGuvdF5rDGPneNA2dypQSU5k7/EbqQZuJmVVq+rWZqfeiKaH
TZeWRYi+SBAlefIiZgaoUQsYeS7gBBsbH5N9vVggUkoTiGW7KTqLxIi3wlnxl9ndInTCs5BdPvD9
oPUCNuwChSwJHSH0xLh2oFj5uEO1piwy/xaQwq7QeSuIHmH/PJu8XguL7JhiV0QbG0m7ZjcF9TQI
DW+b5RxVxE2AymRYaMrVh7XzIuDShVp3HByLXPMOANdXGfbNW/iR2Z7uGEk8MgMbglCPtuxk9AOd
NOmRrjr1sWRo/zPYT3HdHsvj69Gir7Y5WkIYv5dDl7WzomEyzEAikSLJe+XuGoVsftFbVZgiC9vB
a8PZsUbtxoRFINJeUnpwBJdUYWWtdt37s829VujdYvg5oU3QOST+ulcpwIxMgsKZwOJWZt1iXl2H
cxHm82ADDTnpBfwRRlzykHeOrDyCHDLfz4sTtFA72iE260+QnwseCJuaiaPl2z1YDRmsqSd8cCEL
EeXKa6TiTiaTh6wgVyDCz1SMgxkaikwmznPdiuWwxza98o/CkXzNNyUzxWzxAXNFOb6dYF7e3amY
NK12y2OrVwJ4NpDipqhfgU1FAzGMlVvn40ZjqoWyMRyzcTGVGFtoSqhzISGxzD/qlMwvIFo7SM44
vlWc/eXx2AgBglpm4uoyjAGug6QE3CQFIdT2dlOHhzlos+ufB3LAx1X7DSJJzYBL0M0ah0ViolOk
b1yeE3fanftS6UJf7eT4QKUjHu6FFcFzfsmBYBLR9HbJzYGhQNmq9252CR/HrYspHVcLpjIDMJGi
uHpv3fUn8ULDqNCZC67Dlyv/rWKhd2a2FzcRhKF7pTfdw6Lwo/1vN5IDuNww9IwxOury/d6x/Nqp
c+vgnzkUwX+LNB7Lv7I7HDSdh+ImFmifDmMsfELW43R5yV2E8PN3zph69DKwyXbSCpoN7m8AcAH/
WKtmHG5KFYg9BF65tUWkHdPKBNqk3L54Ci3ObP8oTLXNMVj0hVBSe89su8m0ZWNhhTcFRBGt0e2n
mYze9S+klkAl4pFF6UxabG/igwExTzMehUUQWaSDQz4ZfkGNb5m1qYmHqeXZ6oMFKjca8Z4iMX9R
G8pgHW9B3Hhl6bB/WivdMdo8uzPIh2NGGUyeSnZ0pfYBwVh8jcXDYCOX3rw5T5+LIU6f2fuPC6hp
uuum0qNGSH3NMYDmhvcYiYuudo6zeUNiR5FKJhgqiqnvgbwiXSxlDaW+w2aBxGuCxUcodnAHyhPG
/4zCkekvXwzbxfkm9fzkIaQ7AzPnKGbS/Wk3M95oFS87SUfjMX+pJanyZV/pJUNdBOkfma9Z8zW0
jbymY33Aa9tQW2Hfwzv1621Ufodlnlkcj2t8UU+9w5A4p3PKV5/5/pOhU9JSxPGWs2Cvx4Xpaytt
m2wrbdr+vk8dN6BuV9iS5o8otGdJtsQUysCoPyEgQTtrTRuZeYj9uuIH2+YQ67u+APcgaFnOsD6z
QZZnoqfcN49Nq46fW7LmIPiTLwFsIuhgBDPaZGCQwidYnbW1pETkJ9zZCzasfI/f1EwfC5ajoB3p
pOMpVOnIvLBu34CDfrSI8rFOFnUXLat6xytBjyFPAXRXDB7bPRIlMSEb2KQuSm+T580rvau50IS+
eT70gmDhfhvm8olqSqjxzFDTuLAsdhiSbTMhJx3xj/koUrUbNX5uV9DnqPRUup9xk7tELDbZPCtQ
H3dIF1hwwPV1yIGXKSEEk9FBzoRQEg6Bk1aFhnexcWNbZ8G1JjTp9k3HSqDxD3CLN6Yy/CwPw1N+
pJxzUaWSZZX040Vj5gtf5f6M/GBy3G4YNY2PwFe0x6mwbEasSX8bzJprJk1Z4G0EEDBbxvkQT9Y/
QlNEQepuzIUp5imfphHjXiNXkOYaXNeNuDBGf+5q0iKGKalF8p5RlaSiMIHCO4VBTZBOdOAa9H5G
Pswat/qv6te/Pwozk5tOU2sgJLGOv7HM4kB9M2D7gWzE5Oi7rcHwzpnYeIS/wwCTKP6/kl48dTQp
b5JAT2SCF0jpV/36eah7P5F9+6vluktSJABfLZLYKf0yAyun1N99bOkZR/8duJzMWetfZoo1lsCK
JgmIkn/ogSb4ZTC+bqP0+Gk8Su9oeUZzqNI0XkqTpecGlii4pcUnFxioIFTKSVq/G9gFwYE80LVQ
g0OK0gG7A0KSHpWA9tS2b58xUu04h/9s9WnocQ9+dM76LjMu5tafxZ4f0U9alQpatCqZEh8+7clm
f4pjYf/q+T04X/0OHhkE8jRGn0Q6uwcR4sWFgPe/JjlTWm42ZyR8pkboCYfvOS2KiC4wJUfq21RV
yiZRiAnBXVgLLIdPWMsuVdqdq40P8g0dp6AtwP/pItyrlib+B1OdRg6IGoQgH0iiie2cel0ueOu4
IpJXWjRCQNmxhyqsWOAXkGrboNls45iMCqHK1/rdckKoeWn5gjEbTazfqUai/ZryV+DJbVqEIsoC
C/hFNAxB9Gs+vuI70vPdWeAxw+1CVqtYqTqBzfSEuK96bEG1YpUwJ/jMziVtCy6fKdakJjuu8YQb
zF1BkgENf83QEVVMpK/QevG5lQiH6rAQMZPSLNeMFeASSsLsWxhg0EA0nseshcNQ8856fKzd6Cji
GNiqespP4ibpmjqpGZaAalnNv8ZDb+j8X3gPYpbXHUAZZmQjT44YI981PANY2kZy3NHVjMEZYQet
pvdpImmte35luHJLqZX1rFNlGKAhxQviUbY6BVjy4+5i3QHFRk3TuFubYZDrMa2yTwNVaCF/O0OO
zdkkMd32TubSZzFTrISGUKVNnq1rUbML3l0PUTeDuDQHG8cQ0ygrD3Wv827GZp+dOJHP1IkzSQNU
mvV0PQo2S6yZk8jjyrX9qgk+NDHbCIRrHs3HJcYJ1BopcviUc6ouBF0NpsBAKSaPHLuxGswKrhtX
Qu0wlHnBwdSrjt5T8qeu5ksoTDZMaSxWM8GFlCEwwXKqrR0GNYsLSLFxvOZ/y/D/b80QU8GqI2fz
j4VZI2n9pVQgEcSOXu9uKFxFmOFYgu7dEP1Ly2gn3yYoOczxS+fskQSCjVzAzs+HG54nk+QYKAFw
La3gkTcLhLegjErHzrq0xfXgXcBWn6SAgrurjusJflHEtJ8fpYtGtlPIV1qhf0AUFF8dpuq9lsdy
O7shlDI3cN4JQJYD3XFJgH70geqiQ1dPNs1P7OJZSaTkL9qSnQ4HmG94j+ECnDJ2qxvdJVs9UOVu
FmNA7jTcIctjq71C8Cro+kPs8+GgdRwBs4A0sjouQZUIr8T6m21WPm6oP4INo2TkqT0g8QEhj9VH
WwGHzy4oE0IhHPSIjatA2jg3V8DJbyld7tSEnIolnhyf0v5+dqOZWwbzfTOFfcDeZhDMjINz9xzu
yyNoFOMzuSUqQFCS9ybBBR3qahCKNm8j/EVY5P/5LFrKp2Op/wZhHibSF7x4jzdIs7gNdw7yMpGS
4aqPmTsCI36VZ+mSXVbKR7pwPF9ottkbv8OSb35xtaOcTjJjhr3glIiFqnp49NypCCZPlaCQ4P2B
3UO40guXxaEjJ+klY9blqRrGMR2zP5kiicg8avXYJEXDtZ6I3wDyTw7gY8x+Hw7B+Ct2hvUCp66q
QV8DPSPApcR69ru5cM3s/3B33Tkl4MD8phtlgK2y1eYuUc8AAzEfxACS5tWD4spoWqBKevs3P2Tz
ygvnriR50eR2k894GI4C6fSeB7pe20rZogyGR/MmELLf0mgZ1aJy583jWKB8UYhdZMEDIhsHWgG+
mPyus7kSAZr9MdoKOEyPmTIad5jamQu9VsmkKmbUtrP4BX6r+LhaclUyrlAgaYNFBYHsgJJp9uP0
MDIxSgvHF5YRmEp8bQmsFmqQj+xa8oOQ+itPyZYpLf7iTGUIc40x80o7x0JlYZDamV5f/Z6rl3BP
Wl9145LN81ASYp9MBL4iNfrhxZlkOQzM3MGtQw94AfuDGQNReJ9hg+Mi9y2k5hXZ2j6KOAZsgCJL
h8Kll5tTxYvarH/21H1dtcJfzqZs4PNw67LrEAkvQBwcaqRNLaS9jsm+4ktnFE4ioB0cxx6t6Cfy
X9+I6Nj/udT1ZK/FD6VG/YxL2Y+VA3JIFBwm3p86RUrtqPXGgg2hs6+O1Cm5Su7sOMuehXlg1Enl
rN5EK4j0Xnk76dRNJQGYNhn05lGt0dj5QV8pptOOtRQmhgcZRe08Ubsa0PX0aX3eYQ60DvS1AH9F
UUtpVWUcaBGJizie3S5SGZla2vt4GFQP94+PKdOkE5FETg+Ldx5C6X5ZkHI0+cgtzIBA/wTNlJ36
XGru7vGyoigSQ5n98hzm5nWDIaZ9b1BdlJoT5lNW2ffL2ryirjgY3C5DcJYxcXYTtq8tcTJp6Cra
OylKIo/H54w5L55LbjkSpa9jiwSFEYOj3KFMbZv/LBMmiYDYHxuoM3bqG4zgoxbXAPlkmhfLZ1RI
tGo1r48lrqSN6w2K4vtIGlVlTO2f0Dn5VxH9A+9vw13n+yWXVM27UZ8U0sJ0hskTl0YFp7yAHaaT
+9g5nDSls4F44h1zsVa4E8AC2cBG3Euh687Dr0jKKxZHbG9KxQZonRYTQ22YiU/bl1V1E0nsEn+l
FcOS9qtG0zTDYyV93nf7B1ipz5eawloJUiBhmdx4yOqtNc3zWV3veEhUh10pt3gr9JHtKx+Hd9NI
P4N7EnLsURnJ9hrgNFBtOPjxg8Io0zN0l5c0teCmyehaCN8JtfIOLLveGeoI1Vn9gJBU3fpuT2pL
0M3wbol98e7iuZwn32GHdgcryBHpJwKExNcBCveJn6S4N9oLD+FyboRdDlkaKAz0u6rVR0P/Cd7A
vq0kf5+7YAW2IbAbVXf2ag9ctDhsTQf94ymmJCqhNii2HxIuYKCj83iN9AV96m1zHdI0vk/jrpsg
1OA3+LYJUOXo9GmvQBOcWIfow6ygVHl3gm8LKaK/qFMVw35PgDeNIXggOh3Y6Pg+tPTzNk11I7vx
RGbUYlOUe7mxk5KY7K1XoEZ62LBZD0nx/jPgJLQxW+3bTZXm9fqMqeAHjkUgHv/cP6y+vYTd3JP6
Fm9Z7a9nHGFPYnM3d2PguhmCpZb24oGUK1Z3slGbDCjGC/K4kmRAQb3EZiROS2rYQ+Nm2bjoIN22
m98Psk8UP+tF7fUW4FxgA7fWzkdCaiVVHbdG4AAwUDZae/A6RzO+tvM52AwH0LYmjdXyGibXY9xd
fsjE+7RL7z4SN39+gKRKbdcByz3qKwuIyKeXD1sDICULeSQdRZ3SXHPb+HZftSg3nGtJt8q03Dmh
XvZsEeUgrz3XxGSu9ODRPqFKSKQBmhj5UorqL1ZabMtNLim+8rKiSO4Tzdox3vck25cQT3V1oDtP
g0pXyYhRms0aOxegkSubgmwKl+r7NblL55ZACzFNjL2RSmbPA53wCpYQkcmnX75DLwdJLqD9Srpc
DGZs6qrLLG85qGHls39o0imvfCK61O4WTVojsK7PdnvUutT1JOESLwRJMu7ZPBWMjRmpvSWJKpRu
96wbCCAz/4fC1clohHEOBezAVXjaOvvCNd+uSsCyRueb4BqtzYZDAwbKDNrWLAJ689blf95AiPHW
HH2KPq7Ho0kAv/Tbmx60woJCoedh2vHC2ufJ1xRPivsOSbi+Spd1spSOXHc3h9G3IZposXMO1BgL
azc6hUETek+gvAqS/VsoSiBsK0NbYJi+Tk1M/Dxb8t/fTeQzq/Ny53S4wgT2qjkcH5pn4UZf4q1e
ahFoOx09X8kPRv7LrKnXflJVpega8+8m3yo3n9C4VhgWrKrI7QyWu3amyJ43CGI00MDnrtuDXzCr
tvazSpP8+4/YmrzzGJu8kGfJfK1SxE5+1Uu6inS5jQGMGq2EBQCoHuSC4I/R+Wpyu0Hi6HGAkHWY
39N50uV1uXhnEdsUvcnQvV4lLPD0kef/nZbTrOKvAGLVkVsz20sAlTityrkymNU+9iy1zmOZDlQ2
/R2b/iIJLIxi7yY5Gq06QxvPbh1uyUdRjiEObkDX6zp2DWBkGKoDeFSOAYVrvxZDRUkiIW0k45IX
6wQpH43O7IYMtUFC5o+lH+fPOE+SnBWKYvSRmuDoJ9HYdJV8MsmFFh5zPfQ0tDgkpsoG//cb3agA
CSFJTLcxH4rW2HVOMN/5saJGZ7WSNR6Qkil+xexpN/jVvnhSFlokZnjJcaJmlWqWKuvXnzcTdEqi
yHYQS0q7wOUI57B1ig6y3lbMNv7Kf8CSgjXiU6Lt8wb4BvWQS0v92Pozp2r1NU1K41wCdT/Uqfgl
NBZpQxMoIyCpCxbDZRC3rJLJh7n70XnonZ9onRAnylJIxsKuCHy1pv0x4fxSB1VCzY2KUvDsDiw+
os+S3HJyrliAXZMWLeKt9Fo3UnLR+QzaL8uoHPSU+6U9jooFMCVDx2/w1zKa0WDeu53D3uDED8Ag
UWDuq0X/ylwSe8oiJxJu8obE8vChVZvq/BnsfLeLihsSbLlOsAdDAz1ahziLTtq34PGztlSUuO6j
ritjFacIj1F/gDScKa7OKt1um4ZkATkBwMk7Vx35/XjePHZnEQzEDGjbSJ8Pfk5ycpQ/1ESvSDhT
PMED6uU0J7bB7ox4Nh73WVEHYVFeJW2YW0ItEUXmumimI5nJwa4Gk2PF6oLrrVrvDt2rQiHRk2UR
o2VI+jP4zNPvgmOIbFzzOCIwANxlitYOxhVRx6QoN6RXheVFIlusHmC10rq/su2EKtsD37JAh68r
q7C7U7uYhwfbpPkeVxmQw30/TeKtCIlBNMBgp4xmA5WbrVh2o4OHBHeh5Vfs0VQj/1I20i5lrThy
2MZ6SpEBrdgi1hNs3CUfVXvViPUVXHGhgNXJ5Qs5kUENs1owo8AbzcA43vhSmuMsosmscpxVLYaX
pFkoQMSGtBl2NsAQKzDkIfiql20yQQTjoX0/CC1cuSnfF3+TmKFNlFcZ5yHqUdZPaIrk1e6e04nf
Z0C9b53Lbv6ncmQuvOCPpA/qfxvRwHIbcVC2IRLXlGAOGXGC6ppn0rfmEn2GQ5ByJaUe/1fmyw0p
L24BZvjN7c2cEEp4IRFdQ8Jloh3N/GbJLpVD/WyozWHonRKQCA3+kMagzECXjJlVuUHQOQhkyysX
W6HGSLThyUY8RNdD8c0wSIvQxce1RU3a1XXTVRMxfTWjKT/Jy6KPYYcsziPYOMVh/WCYTX+s6dRd
xNBCxPaaEROeUXoNDDVAWmveSgxMnzNAtnMm/lwsIQRmii0mqQj7TodxA0LHFSXqN2fNuxb/MxzP
x/pknbHiOl7YI7MevEWFPmPyO9hUezIsqoXtv0uclLOCYThO/KRPkg/xcxTPb/CfTEI8F7zJ2hrL
78tMPbSl3A6a5a9jEQiI+KEy58cutIKY8M6661AT+L4hdRZ4tItXAFq+AvcF5G6uugMQ9ERKPW5o
Ru/tutZeKxefOovbQJGHBHDrA1BUziRAciaQt94qhiRYm6ecxzaEdidWIYlEUd+U4alX/hdfW/5U
sDvlBlGdH7kvJKFmzOt94Ri/lrMUF4jSm3i16XBxuXsjEt2UZ7IJWb2ovrm6VRgvzOTrYvs99bjL
IjHirB2s4zvrCIjxrCAQMp2f2ieotSnEi/Prwvh7anL4G7T7dsfN9h3NOtfdloLtn28CXZx0t31Q
PjQu4ownFuCXqWGob19IYIphBRI89E3ig0+xzL4aXRIspJXJuHv0P1tlgwogLLaQsqMX/6guhG8Z
AgZvnZvS+WgfFcD8uaQzYM9FTLBFUWD0BSSrTo8hpp7vSE59uLu/Tk7G3+ZcO1CNgG5FejbVyeEu
kUwt6I6ZHPwaQ+CxFvp/XGGopQWWe0httnAU4Wx4vwlccsewOPG9oVYHqMBeeUe5ju6c32g+EhzM
XwlBm+kx2JprD7xCoVP6KV6KlYUd1JO+F0VdCS7PD+WA83EGu2qTY78jL4SM0/wvTTWdWWrN3kzR
cGnwkKb01Vrik4mo/A6Y1gAewtVYgSnDrp7ojB4XpL1Lb6xsk85/0QkIIOMhC9JCZq6ydE/2g3/x
/ry736ueGRm643GJo+Dpr0qFIO99DATzzt6PMpL6YYYbXL1hYxzwLOhw/m2vn7JsqmtfI+bKtNyk
KYj9us4tzWUspjX8qdXascRsOHtrNkydGsixHcdGRqlJjO0ezgkgK0EsU7BnIn/12PO6/unI4QRy
xj7fB6RbNonLPKLwxeTNKO7v7f4RDjkvYAZ4WHbRj7JM6G/ygeKFsfO4IiwZ/75UKbcgxXFbMS2Y
sm2JcW48uFFFcPk8b028/tWL5B5trSJfA6eF2oHCW955vjBgyxFLnyzSTmPHhHEh8kVownhl3K3B
L7JHBhgBNIHMUeyu2MyWjRbu+iyAC8QvazL/thGp3YrOuw6z0GgJpt8DfjK74VhlYZIVhZK0ZorH
L7so9sL6kto8eShUtPMmrm0wIB3P9tSNbjBn/+boVvGYILRDO44tLJ6djT/PKHkvBWmf01OY+AWI
pQlarQ/W9dpZ2cHRSvXzqkXkSOnikHJU5wySOgW3rAhTB/112igyHg/CR9vvd/U87++mYJKqSBeW
sI7bjZ8LMC6JzNr7CpYNGPxkJ9aPoAfg7BoDWrJCYinsUYpW+OyWbFYpsP12+DHyBK5fXPzzArAO
Cf7kf8JCo+g1IKI6TDY2G2/deO+rLf8xB9ibxOJQ+1T9yfm2a3rD6v4dizhtQqidat/K/CsjMtQX
19yD0Zy11gyxdyZuJ6gangvqzz6na/MIoRBbcK7O1j98qvJnYi/t0CcD/bekmHSG/TXgezQT5/vS
NgnRWIVX6JQV+YUw1hiZpotI3p/jywhag0mmDfqTFVmIkBsuUexd7dg7UeCTVikE/w2I1JoF98a3
FKrrU3Mm2P2YeXt73HYVbqo/PTYx0pL+S8kw9MG0INDHbDVBgV/PpvORO6I5aMYXNvW18335FWV+
eMY4Eq447L6JzAkocE6dhn+rWXR+i5UcWNWEIf0eORULEBi/ou6ms5T1kQfb5pmRmAbeUJPe76Dd
scPwlD5lQq636eRGQyythoEOYSDFPqA7plwlz0Vv0ZiuSx2LDz2uFfKZIMzzvCJBwsCkrUsGNHNV
x9UcMRAaDFWBDfaey94fFAQnkre/Fv/8+Ge4ifhlPTmd0KBuFHYD8K+npaZPJNHxorx9Wmxpl3Yi
tQOKjnlShEGFgJKgrkcEHIS0bm+HP7G8hVUzmdDVLYfS3pCDE+vq/5kfIqXefKFhsNh6bbR/7De3
1jTfiDnCixzfkQzL3xf9eIp7UehahXjViPi7jnlFwEw4sdH8cm15KfP8Al55/RWD+VHv+Gspu1UK
u89Tsl7OkonPpyuBnCP+bDJWIjBX8oufEsRN96IRBjS4ZhSOrKWAypgftoIIG9dY71YKuRRyxLg0
aMPIS+gZFaHyWXrPbN37tEKAYqURg5QK75QVYg+qAVEVrSGhZY5NurPQlymbhoY72fSfdJYEK0hR
Quulr+hM9SGilYUGFUhCb8UgTOxzBFUn3u8P/5OcU8K+pDTFNb7quvHn+TfYdL7jdV9aM052obFC
jay8xlWeTYsr1O30ugNtoDDupfa3gPkNi4PtRbFhR5Mkbmm/FkTmRqZt3xfL0xLyXzGDDha3Xmvm
d9duRcN67ijPvQISGD5VQv8PlNqhThvq2ebzvhquvdhB6ewZkkp0fhEsYWSG+ysdaBgJUdesR6+s
anNJn5YVhpQsXULn1/KBHffwnunktKejsk2OdWYbep9lf7+CVxtOMxtej+w49cJJOetp/4t+SU19
PmH8+nZuWPBJ9GlcHkE8nioi49uTVxSbL3jZhIhdE1hqED0DJIx4qXf57oqbMG0Or/4LqaUQZFS7
11xzQP6npI60FZBDSQ44L51nXcndhvmfhDoiI02zDD4AkNPnt7haiRbdoolCJwm1Q/8QXra+HLXV
p+NIjv4Z0XK82LWQfWPjdy5/+kt9n70QNVV/F11SNxl2SbxMBTcomMQWdkWgRDjZkA/n+ul0QcOc
Kd0lJkkDrO6ckg3f/2Za7t4UZLSSVgJ7cW9H/WFH4q9yFA8XVyyiz8t+PkSvNlQq4MxzYHmaLsII
xa8JiOlge+qh7SC/rNuh0CFip64bF3Radf/MSB+JTCM8QoR8dlGb235brCrz1P/R4kQvcNNC+0nJ
FTpT3JzXGh7Kjyl63mEckzZZV7inowQLXqOFpt/SdnZsTxDFykuAC/O20VXbuADtukt+ujGu7gfb
EI5UvC8hqb9LIOCpYuD+SDMQfnpiJx/1WRPvusEf2wa0qaukFATCt6CVK4TnvyIkOxmDL6mZXpxb
j8ShBANWjdB6uYyx5crKO5DJ6hJOxswdMb6zoecX29p2xv3n9ANtiMrxKU7tjLUrNAq6DI7k2E7P
FIDT3HBbaV3DVxevb31wGi/30lOW/WsTW7adBZ1Nbqod2iR8ypmNKQZ427oRP6IHWZNivGGYa+5T
Kavgsmv4WPOchaGyoF+Q+LhcL/jXGHKc4YhGO/roJiONeSVHPX2Sl/yRVzlp/AKjqT74764XJK0y
M2ACOycXKZdF4AeZ25P8Xo11/hVfuPaVtAPeekK4ocDSrdUDYo03wHu8OLHumRlX0CWhvoCLnTik
CEkazdzfgaczgUVZm7i3M5WwSqMIQ4Fn8cvdHKz8cDNSwLCXMiLAf+1LLjfFtWTxZoUzzcasvhHM
/DFHLURmfJK+l2LQUzlyMHHXyTMPswkdTfx1vxUZASJl71LKsPP1oKicO7O0NyAVKYDlZANAlHMk
JL8f4m/XVsjB69oqM3X/dtuf46AlYo+kZReq8jA1orT5vYujRqZ4dZ/FS+464oLhfGTbMOu/uThY
PrQGUhK9wCPVTDUFWzkwNmXm8KZs7aa6xu7QE6eI1jM9A9SdsOOMjEp9LsDW6zgO0n5clDMKkTMe
La8MYhlD4FPjIPCUaih/k2dqfX/p5P21erJZNJBH68xHqanm6oha6mTFz/51pH+rEZWzysDElTZ5
Wc3LMtfaew9S3vqIRw/TT/zf7aZObUBdSDFKJJ4w1F7FtRy/cih4tqBgMD0ttQ/z1SubunYPo1eF
RkqF8CpWlVXvRdysb+S6uCk3oC+uhjen5A+KtvMPKl1BNekp3f/yyfqO42vXqZEJSoP3LQJfImJv
x3ycfIEQYy1GsgNhAksAvPiEW5tqckgwvm2VNppQXy0yvr98ScERS4jfYvU9r94viQ9IAq9CLsTm
9EGvZehKGi/ak9fsy7PyCjoPKHPzhsPPrYMaUKYlfxXjq0ZbtjvGFD5lR3P5RkRqnvMHkTYGlaGO
LsWWc8X+2tcv6GQPzz+cKkM1PUISQPixkk26EN6EdpHC/4Nyk5K5Pfha39J0Re8pgu8cMQFCWLFz
haOexpaq7o+BxkY6j0JwG/76I+IoyeVujkh4cpWsM4pn+yj/JIQgzG010/7FGBVJG4Iam0danIyS
uBYY6RY96tTtw5+5LWb5aQzuagYTAKgc9ldjDmBI6M5l6LsALkHo44HZno5ZhZxG8YSy29hSZuDq
00IWU4K9ejD2hUNTCfMLTe6AZkR+zudN+HFJntxaE/gxpv5IrF/lcJcdsRjoaXKElSlktlxoKivr
6mlbsDLlIocWpccdgq9ZNdw/uHFbmGMKk8pmS5THEzKsHDQVufizx0zZL+TzhQA9ROBMWwLmjPTk
QTJHU2fsomc5KezV++FWq/ggfCIgkfEHJ5moWaAIrFnBIvVwRdu1obNXCNvhC7HLtqymIimMC25b
2EQLClnUY4uekXycr3pe1vZUL19GDDdv7V/85MWsjTq6XTxsw1i9eWJ39sZCyzj7haclEJ5YN7EB
wAPlSQVVwipYRPLd+6GJQYYJdnXVIgpKPl2g4HVYCmCg+SRDgLVBOj6MW3ZzZWUzj8/gCWxq8lJv
NP+LtVMxlqItgbWc3K4heydRe13W9f1q3xQRRdlRF9Q9xYSPA4ZErW2IXTDY3nSwQh5fiMxcfLbo
b+bM5MSnvNzBGohP5jg/LoOMdvvPfYnW3L984lvNmcahhW7JTQzBfjruWZk/0rOoZPwGP9aHQdbR
5wGuu6YnDQokJv5ctqE16fADlPRiv6u1axoSk8Vu75f477WNKRc2j4QJZPYQVmywjgwnAOIr1ye+
xNwGPPY1vyOVAusw/SP5KSgr5EMI/8Hzk0mtuNaXUgAdyWgzDf70ucgSozlnIG2Bzd0ruXxDMgP4
BF9+cZVjTC9HDAWPZlM8aFGo0rObXNZO2b5xI6ICbR1ig4LSOkiRFXoII0JjA1AdIxhEysg6PlWw
zddZ3KhBy5HrOH/8qRv69W+P3qDQpfbiMyiOTIowV9CS+dy50kPm06KJXAVkA5mKZeCSAHQQNDq7
cmruLHlgkOr6Pd52nIy+1HXvtt/Bt4UwSiFfoCVINh/PlaDm3nPitHjzzIaSyHf7sQNgJoZJwhNO
/OW7z7QfYt/31GEWyLhCXG3HCkJthRvzZ1svH3EdTNupBxkbqA01TGsXy+o7p0fQ7SadoKh7MBPz
nM5sinhFw6jWzi1sJH/LGEG19KQN6zp2ObFl9p2lbHBW6qutKWQVka+mxAE6Pil6dKwuqN6ysk/B
ZXOIJ7OBMMpHY6CjBdQdLWEwTJjjXkC+GFgJqdVwGMQEN8rJVaeAnHWqBe9r+9hBkB8Cdh/6TW0S
qrw+vk+/ztpSNaswfvpI7r6X5zC/pDM50mXqc+lbeE9//hsaEZzD+Jb5Q8akJ/VQbvKP3sMhLive
k5Y8lmWNv5Su9Gvf01izqgNMeLXQwh/S3vwMq4pv9XB9Cz9P+yWTq0ShYzoZ4ttKkZMz/ceNVN2w
axTOQH871ukaU03jv1hhVzNRZ5osce+/HqUguPlKqOeVlgJRzV05pT4ZaVpgbCCmgQNFTO2a4cy5
kkVRDYMv6X5JwebzPWElwHo5P5OLFwgG/BpSfbYgnAyPFHxikN7OBEpRpqCjXzZ5ZSLykiHdEOat
MBhsVPUl8ayltep9Tn14BGRi5eIezGG9pD1uxojUiiAwd27B8k64F90+vkXISVrf8Uih0WMDrPJ/
d45a7scKgcWR802NB0x4K1AHpR4ZqfTS5PIwj6WImk/Mg/v0mcja2fXgfcCKO0tsNNKHOC8KWGM4
xr/rqwTa5NrDNpKEbGRfeFuO09xYxeqWiFGcnoPedKqlrBdK+3Bi+wI2+QISWZfWr1WtX5TdD3Lh
Aixe3nBY8PZtr54ntbpSRKUQK5RcM1RE2x0qf/iqgFUYIyWkhOCv4v2GaiGBQaDvdn79lXUnQL5I
H3CGgQGKWI6pJ2gdaiG2VNDO6Dc1s1bT4UW7EDRUfHU9TzNDKWr5TqlcOPcZOLeUFdqsBOz5+3PU
rfSfMyMLDRIRhKjaMi7R+SJZONbcWP2gWXFs3vcZVw53Xptb1+4YN2eb7n+EP9XbamHZGZhcYiEA
fIyJ6cjAlSnAl0sLWVRJZnT36kNkBVg9vQ/2JImII2iLZcuUMN2FylQ0IJpp0OhGV9zsCRiX31F2
zD1nYBeE6MmPxFjXVWljQ27xdjgxRKMR3HBw2QKoBHA2U0739xSjLG89XqKHtnngDLhjHRItKClk
eINogaHNz6aSTEy+5IFJQiWyXxMQvLv30uKWFQRcHcfT4YaG/PIAW2M4uV4XlV1jCU9tn+4L64lq
wKWVM9k5x9pdv6qHMTA9Fw3Dsan14kIK8nqAW3dOfX9GLhZ7LQgyRfmKxPOJwpmaGa0z52Ld4i30
CnPVu6W/mR8YGlzlMFCXJtThrZFAbBlDNR+GYnWqhCuON7L3crjAmxkNqJUrg/EF5OSLnwixNO9i
bdiNi5hHKKloiYCbPh7sGNbeywZ2nenHKjlx3b2IoHCeJPN4rPmYQ8Z+fV/1wdK/fj1LRktffNU/
tZ1LwDD2EGSfhjwLKgm4ELUzHy7uSu35iNAFCdM2h7ukJ76hbyvVHf5T/TrAWpg69nUG4jFnmGi6
XahHXCRnCMF/M8j3bwdPy5P57Z/XBNTTA9MvBm4aRaASVjNIxZhlYeacjfbe+Wy+oChlobT+3OuB
rkoi8IYijUFsxITkXyuXrqoomvcS2hqSBGu7fxPaWqMcQ36rY5SN+CrtljMQQCaD8QGyqkvZwZ+b
rJuW69LDqSvbcJmg+bRB+0BewSSYKsGXejN1RNHfWVgp/gzCN3be0jtcD2wC/fED1YpChje8yQpm
8Vgv5KBJkP1CR05wZoWU41K7OysKVYXuQDDXKJNuuOWjF6GE+pJOSzP5TJ7zmmrMuuXyabMJA5sw
0cFXYgX14SLfkackWPll95sT7tn6lmju0tC1SOdSdJ2HVgU3Stz9TCzuEVIuDxxah1XJx4YTq60Y
xMM4xKkaYNNHqFbOzwn4R9kRF8xQv71xYJb5sJ/tAtXBNTogrAnFjPWZw0Y0bOyelS/GgJ0qlKbv
wMd43O7h0psJSIFOiyzPAwfjpEBzxhUQYVkg8CQM5+LI+0MomwtyCQSHrba+RhHqghDw4K8lZs6S
IMm+syCTDS9FkwVBvZGHjkBf7pru9FOsWWT3GEKzAMOSVp+TgiU/v4deAD4gL+yfKDCq7KA6qSBH
COuonZnxG9cASoEraDyBE7298wK+kexI3il4eZOKJTNd62AKbYddk610E4YJcIh/wOjKYGr0NOXy
YDbD9GGqSfUav05v2WHH9+XHVovMzrHYaSjyqmFJG5jg0cnoAnD8ARc0ThnetytIfR+39hswGI5v
FULCOOwXAofOP6MKC+wLejWEa3OvoiE72qS1r9hd6FhxoqJo7tS/8bX2RhAJWyc844kmEFjCx9hO
4Ay7V7jbuZWNIvH1X9qiChGdZ6Q7Atj7ySSm4XscfacBbkvrygAln9mCOZidErLmp1yv8VT5QKT3
fvXDmiapIlKb+/sd6fttPGOFfuK10ZYHysqjYwQYkn6UkHLB5X9SHwcBHI12JE+pWekF0Tr5VhvI
mXiYMBZ4aWBoHIzg0IQzU7g91J7o+9CiZfw1h7xMGQRJlb2TJ/aLbcwIAUdlbG83GFz09uGNNUzP
GJrRJXlNqcKoBIALXiTh6mToPjRBDlAKgsbbN65bR9BD8P0HBtQeHJU9yfWA5U23sFJon7lQSEWq
5jaOXtIoTQtd5w4vO4+z/7d3OOSZJtqPk8mhxZjRLBemKrUv10wSxmIIfrYGXYDkyafJyzpEP4Hp
bqFHlYTpeY+pq9gk0nRIDduirBuIOkQ5wsAp1WwW5EW25YWq+sj//zz2ZoGL8LLfNpRNgsAPiqvm
CH+lxNnxRbPIiuMeSiDvjcP31BtY9WnBBvtfE4501ltVMRvkr9GRPJJnbARnW24yE1BVvVPkbH6B
7aOBiAaInD3TBpVcI9P4Rz7oAzPNHkPWp1wDTZAMYN+FVMWFY9sH9kFsSwaIg/jgZ02YnluAZlOr
FTBHG9+nu0eazl1wWL917IOgEkOzKNbRfubD3y1sLawOprs4CGH42oPjUPJmyz8KK2BEqZxPyMrU
casX2oiSMG2opBQ3QLWfJkWAiy3qmC9OBFtNiuLf0KVSNZQ1fnfT6r5tFuHHSxltETzgZeNf8Rn9
n3vHFI4R8d5cUGrL+OY9cjKsWYJVhgmFWYrFLOeyIVMSXP4gXld7g84EVinAx2P114qrJ/9RbIj0
k2dn0mWP5hx8XOuaeyPRsFdrRNwMQz52JM3hqebS+dquRlLWychYScaXGC6hjnKG/qyHQX2PClUk
ag5swjcrjN0smeSv8dqcd4lKhf6ijZ7ea7cNtftIxFVG74DbNc675Np9ihaNy1UZGdfN4t1MXw5+
vQzsVnLYQbNXppzt8ssTEudbbWMozNUJOVLOB4lfQc4rEt7BAe/C5VG8UhytOaeLQaGkHDlMO6dd
YURYGQKSRnYdg/XlXCNnOJiUrfKLJ27kDeUZWy7ick9V23LHSf0lPloFCP5irQzAlxex+oGJ59gv
Q8KPxmeDhU731OyugG3+h9RucG6o3LDw6twTKOBJWxMMpj7Wy8NV7Allz8NnbfxlnuGhGHVCrTzm
ZcBkMGknToFPw/KbIplJPqsTZXKy+REXRd+NMf9LtkjcpEZ9vts2lsu6G4CrxYkkEBJYhjch6qCp
63p0SrMVlF+4EoVYYWRhjTIKBdsHsNOsgvkkQID3YFLziZ6VfPsBrft8ATuWIJrd6PCvwT8y1MIV
ohISt9uEP7kIktp2hi8KZv1DbZK8M44O/6oSGDanai8Ygmn7c+0jCcWvaSINAXlUOnY6V50qUKeY
fdDE6daWIWZoqEkLcv6Jm5tDzACYPPCLr+FMdQhuUdRL5lbJ0zytdaOPz68wvcFDPJdCAwV/2ggy
7YtvhB9HMUwfyacA1ZEXpW4cMgClrQDi8kO+t6QCd6ngw7aXR7+ECW4zXOxNENwQBcmuI42qRmHh
PEDatrGlLiSnN4vCkKRfQxFSQ7JWaLlyfr9cMYw7HqIfp8uSSwG/vsbqkJsB3I9r7SQHxFzdtbkB
JDE8UgclzXQTb5aN1HILBJ73Pgq0rkrXTVFRDQYTwdF8uFRwFiw3vKrqS8KnWJmQZXrtpHpXb8mM
vGWzPAJxKdMRX6DNtWkGw2D852wYGaAZY4oZAGZ6lZwCQkVr/OnxebhLFZyiNSI/+n4KhtGGPBDX
cm1omDyNDmEdRrNeoD2IsQHTGxMOBfEMAVjUvS7G3/bNHOq/7UgdnjULnqd42pCzM5bVC+sgykHw
8SV3q8U8hq1sf6I7Sw1UE83c9QvIp0jfeboirb+DfI7Ep6yoswC+n2k+xtqRe6A7KBIe6Ub5qItO
GPW1z1Bmjs2Xa2Z+o3aORPUthh3XRw8eQLEbbSycnQmznMS74h7pA+LBQFhNCTnv8T/Lq9tENK9J
WKx4Pg43YpRbA9fiB+ATalSe/xLf+PWwGA8mmLTwNWK2CKjwzh6CACtZr3S9/RnxTR8BMDETAU3i
f9HdU5X0MsPMvrnY3NdQRmmh2uxFdyZGicKwQK7xjGlBWnwy6Ot0p4LnbCPaaB6Ves1S3dVy1DOh
9AhUAUla+AdSJmFFbKZtTF7MAMEgV4gQXYFK/2nWljybEOp20qY14KYfH1Bqppz8reeO0kzHHRv9
wJl+apb3M9kd80TEcWa6DgOPQXQi/WLlgn73X9ytPz4a37Y6mXzSYw1Ndt0GGr58NHCx4wHAQZiD
IY4NVport2Dp8xbAo/vzoNYuirSb8O4y5PZzAGvXBr4Ra4e8yyVbBqDNqbO4VZbZP/T3xWs3Guof
CkAlfbokni/KGHpyynaabLmHEliRu7FbYmfbZJQ9Xum24/fLpQ28RibbvJDTgZeHRz0t4h2kSvD8
b4+clvlreH4/cHLVPsSS6gykl5lFeD4Qn4cFbBv3lgMNoTWmrQTuF/Yoao9fMioe3ROcT43s0pym
o3GcUyezoxkPNpiUPSY0KAbVthimWbBhNQPcC1qUKogZsR0f7AdyYgejaSyphU4fijbZYByScCfa
rxOL910dCz8VfDQ0tNGg2PjCk4FYalaBioKmI9S2HvGtPw43fNiSNcpH42Y1Hxn8AAxqazwtDpsz
GnT+YOB0Dn+pHnoBYclcrCC3NHm7ACITuIl+Yjqxet5iHsr2NEiEZ69XSJc25NwnVFHX8tDoCZrJ
K8+S3npUXWNjJXezLxr8mDsVOu8GWSKL9M5ygcB7zbqG4oTjTzPvWwOfJZIof/n1UQUUUx20qgfq
Y2eqVDd/lqw5HEFoDW1xGD4N5vDHGM0Rjz9lthC3AIF6VOg6LQDhMtMW2huEzBZj/PsOu8KXR57c
njhiV8aY0JLh53fbPdp2YLwD081e+tRRrrCyKBOQNjfmEuf4Goud4lDbf9JAwK1dTU7KEh834Q4E
MoqKeAWP1nrClGuDxd7hrTMQBCncaWgNq1rY0VvluDovrJtZNp9MD/kNRdJOLnz7JM7EbnCXm7s7
rPWQF31tvOWRz6jqjIYrg1xeybTx+K0EYFcFuG5kqHuXKiLhBQkKSbC+RYxPvoKf530QeABe2Jph
SsnquuN/oFjWlqYiRFlcx3Vh0B2d7JbXuN7oryQOzZxQSX3y7s1bPMAp+Ahe4JRsmGd4hEinsRew
9jWDMnynXS7vaobL4kVFcHGdzRfWbC88o4VSL12R1rS1juS0zgZXP2Iykzp3w3ozC62+57S2oxNi
XpJbUKIbYfWuKBjCU1GdMtUMsKQVbMsSvcS9J4m+bMvbb308obFe5mtzOY82zpvKcpSlI153o3Ke
Hy2AmVyqVvrH38agbC0Hl1p7phCUEinXGUSYmAAcZBrBshun4412pzSrHf6Wy0aH5k4t7CUVKZC5
BscF0lY4wSUo8Uc8NG+3XBJTkom92PAaYhAK6V7wQNzTXZi7dQgg630/1wVhiegH/qaCU4uueuE4
Af1wvpoRSna4PFMbyDmDruXGKyoPaev5q89MjocQXMOwXIIekIVxt1pTzng5Ja5RauH6+OITIcwj
Z+v0mgu23eBc0VbAG1k5BYT9BXY5xC4A/U0GF4oBdpN58poCKhSAsMj1sp14yCJD3DgxSidJBCwD
UbiPWCdUCZzaP+Opuoy9COaY4OLIsG3COyqNIjRXT5eY1BhuYKDPcf9yQ6XagKePwHeyuxOc22Nn
CW/wKsgZEyZGbqw9RUfe8lN8F4YDQwr+fpdcCIQ7YrqXZqdmFgfO7pA6PS7B8zbO/cJLkZ2IJ6Js
wyH+v56aklFGsCqwEE1JMsN2MvuG5ahj7nUil6HtZD7zv+NipvrWBv7opBgwQkeL8hagCH1WNR9D
HIZ4aPA+ZzEMgEHqzUZUc6ZZFPF17YqHDx/9Gogm8ezInC2qGCXseEeI+rQl3kbKLUkdziXyWMtz
NXECG1Apuz2Y7OU57quoAgLZX1eFJjWSkXrrhRb1X6D3hmAMW2xTjcdVtDohYqrD+cBEB3R53IEd
RTxHXBZ49Ttf12ETMIfERrPdMHLT0pOpd46//060Vf8L9zxNduGxkpyHHuDFGErxMeg/kydD3D7O
XTymI53ejHzgncRVMRR7QaeHVkj4wx7k6vw8tZBC7paWZ6363lrONy3AhcL9cJX3dGhk5ITYJ5UI
76ulhmlvHMxz3FsINB0eVAjKG/+iCRBn68xHRXbTBug2N7rPpIkqBPRq/dMDDXNK6D2DamMM8mcB
Jh/AcoeP3buvdXjWu7GHw8vNV5HlmKIze5QsOYTHwu3cYiqXXZ/5ZdksmSHZksmsj9LWHI1ZMUOh
Sj+DhELTH8wnu8uYN2dRq6tyWxGWGAr8DP0jHbQmoq1cuLqA7iJxJ2MAEc87gHfy/2HYP8P2D/b8
vYN97rFVB96ZFQLNgxR54xFwFmN3tg/5cRojSn7Klx8q+4z9pgSCwJsmkS8LyCOHf8Gh5e5jGArC
d/bQLaDK/uPDTsvoB+ftRvSI6pzFl9V5iLhIT6D9bDdeYbZ19O2JODI+vX9sk8BufGV6SBjJLnzr
/YVzaO12UQzfzS8IsjiTFBYO5V1midWmiIgmtMIq9kphR8F8hgaKBWx8Ps0wyz0T3XMaMQb0xE2L
SCKmYYe/ohfE8pbp4G8nnAcZAXXUa98x5vXSyVfcFy7EpdtS9M4gh0mUkcHQoPVJy+BQMBqOZRq2
dmtdLclVpINVcqRfdP4yZXog1XfZcE/RtgcoRvRzeBKIiP0tDaWP4XX/gw/OGpxzOqhfY/qQFsip
hlT7qEMFXV02N2mbqpDo/a7gfiP0xLoKCR27yuwiDPC0xgkVakeIxGY2iJT9K6GW6Wm7ltpkig+a
WTLaAaHqUfex6N8ldy5mhnFzJ89IaaUZ104YS+FSAEvLqwBvB3F2sunjSxHBDuK0hUrRHjwv9uC0
6SWvE/sEKmF+N4jbiWwD/5ic7DVPRolwyZTCatYCvnoTKSD9HNJ7XQbgd006u7kQg97aPQE0Xxr5
uy4UJudUEOHZxgVThitBjo9699ayBWxKu+dWg8TQLTUmRwNwu0ack1iueAj87jQNbgpRKMgiaPJo
g2lXj4jHPsbMjccvs8IiVzlL6ZONnehM305hBfRPdrGY7oSK/3Or3tKGhkJ1HQsYIxAqxdHOtHhq
ZUdgJx7H4eHx/G1wv1ng1nDJwDvOBgDarkahGsyyG3mopZs3z3ssF0/dtZJa5fSQD85j1m5/JPNc
9pyuJ8d86OaChqZZDE46MGtPOnOUVpUGa4ElFoXvgvXUXtH/Ciqa0AMFW5MdTdHVIfYKOEpjHUhW
E0dGE/Sk4XkTX5lw1ExO3a8OtwXqUxT0Syoikwg0XucZbi8pIFWbYrjEJXVIRJVreYaY+20dysnj
yplj9jOHPUTZN32b2e6faPSX1b88eYb13nJtuIAQtZSFcsmgpplZIElyGJSSEKHsn4Bpk0HH7KJk
2CEcWZBB8fwRlahUbJcHLSxiN0e4Qg84Fqi1m0Ur851zVbAiFIH1oJiuE9E33vKLu99VPsOTbFtJ
jthv05hBJLlL5wVFT6rTK6n2SH6MFmBy1mrcG8YwgC3DoywP001hJuSMXP5Cigq0DTCivBZiYktp
okf/3aEZzo7888u2AJMLpMvFzFFcyz7E3dSWNbbzWnokeZT0su0OrRnoIbyh6A+nrM7mxGn+zOyh
dPiP53GLaODmtSwuUM/18tom5ESrhe1Xpjfn/TfK2Aqf452vCJ6KpExmnbBKk4GxxbGpTB7QaMbf
Jrs1rTA/5fUrqzP6OfExkUNKWImjwQV0hBq/fyslzz9AHm9SXJWGv33sMrHEOaKH1dcvm+hXnFH7
RVSzb2HNqxyFGFOhmGE8+AbMozssMbt1ni/u5+41y5kF5OQCJFHomcOsZhe2vmOtxsjPq15Amvr9
3q4IOrsXZzYbWUaCKAuojKLT/mNiqrm3zdETqDWIa1azZMvLGvv9ZvR+ghUIUkSOXIzbB34w+uMc
+CXQ8n4XMhwo66iw+/AldMGyeQvWBkPvjEcwFMjjWlx0mIMESF3FhNnCrVrHRLXFrO3jB4jDSlEP
BL8Dj2mlvlqOmrmsDSMz8R1sqwhvNbSRFcJOlCB9t1mz0pepwx02F5+k40UZSqquoPtAaE4fC+mS
5mS+IbaMV73SJOMXrePqbjUr8Z/83rlZyYRD0E+wkvqk3AjUlkk5wdltySGAORmIbSCy/J9DIaZe
U/r53azKeQKR3JuET8vUsFEAioSfD9ru6kjiA3WVrFdUIU38tZaqEshjpFEz5KnpcAPGvGy4pDOF
ShffUGqHO5PDCk1MRdWyFkdwx+t+26fwyEMYzv6HlK+AJd1MMW21xiFsaZVwihhqaM162XrXwPZh
b7MuynTj8anVe02SP84CaGk8PQbgy1JrerKSUObNGrohx5x9rJ8gjP9vnCDhx+jIiL/R4VfEowfC
Kw50qpLgCV1cGo92RRw/fHHfA4dAZBnPRrievYd10KOMMdw5G53ObRZBxREppkzjcPbFEXGTkigQ
0vEratpszH3iaKFaHtB09VLpcHo3BVBV1Am2NN3sXX4zRYb0XqCeiz3oiaUpYFkS05a61Kz+bSci
BWKw6BAZAYwMYaKK6MbP55atRuxKZ1mY4e8bxqbdNMN+SdzIEcwAS456619ytG/IBQPhA6VlI1fG
2YxZxiBjokhy6rZjjqyViEOgGavL77sZ3ysJaXwJ0BPivguJp5IGhaQ1f+CbIfcFY9GGJ3nbNE0y
MrLU1WHrRzN3FTYVocT5AxqHFFK6Mme+FETv14gGEUTMc8kK4/yyMnJWhKbmI3dzGwWAvT7wBafD
7l2116lB4Q5nAfYH+bd0p+q4sn3nnhhVHnEjUW1XS7tYv5SUVPAoE0jFBYWnFDHNzaPmdK2ac+wR
Cl71Kvcb2tnliRrWlAebIoPYTv0lpEZ1dKnkb4XNoaypKNmJLSu7ZOwo3tY8fZn5Qx/WoW+VvO5U
u0XmP6/ZpxDD+70opkBYuUSy/kVtqMKKclf9AsMxS61c6UWxJBfPLgNN9Txq7xJPI4BHwIJePDlA
lAvB9XZyxkHuXng7H/VSo5nnGdZxslQLrogVyXQq/q9KOqCGpSPjQ4a8/4sULmGth7XkHlEQu1Sb
6ra2K/Z0Mhkhl/blzJyjTuu7tyFw26MhGfQAUacTIPyTRrGNEVRiWfvazFztKtkEODFSwkzVA4AY
BNfDmY1geR3i1wbOGbhVn3pN8BSFsGShb0PKyBxmQ0NC7YAo4byf3qmy+R0hXN9zXn0yS/hvWxJv
Xla+Uql5Fe/yg2VU1s267gDDBS/GaZooRCGq0n9hjFLIfySN9wf/DKybrVKsyr1eFr+Ay/JK35A+
jEjI3EaA8JKlsuh6N2O9XlBQIX4A3VopEea6vgEhFSERO1JAIS/SAiDjLql+2sjj81l6QvY4fU3G
8mhzrQ0fmJz+A7SpFaN5CSuFY5o+k5CTpN60sniKJpq+oD351rkmugATpeX0FoYqYlOr3b3zQ6NJ
gpkhh783I33DxQFGRvOTgLxKYC6B9rW6fJDnTPqYwJGGpko/ucy3rRmZ3W+yid+YTIkQGdpozWD2
OC0kTy/NIZIHzie6ErgQHou19Jsdl7t+MFUgDtxnaZYTtR1mi/nC63LUmDYT5TDw2NMohIgwH2GQ
oVAv5Q7L1tni9kAQybCfjruCMBvIaSUmRiigs1oW+UpjCdwnpPOKAfxDUodcy7JUwjYwdMKsLTD5
kMi+p6sMrEvrAEs2rqzENsuuChhoeDK4hCQQ1OY8WKsmvSBjJkqW6q/73tXxaJshv3T2OIJW1x3N
+6e2zKG+d6ymwoP8Mn8k3UPdjUDem8dwqpx8zg99SxrXiLiqytRK5eaDF5xsBeeG/ivZizhtIbCw
46XdnKJ3bvRHG2yvXfbPMXY3qiCnZg8YrrHGTqzXOzDNPNPcqZHgWmfQU7XSckCjnMGUY8HaTKby
0OlGXuCwveUMRg702nkMa5IAhKBJMgoVWSN6ARIAKt25H95IYGclgQNuuW6QleMKCWtGQsupDTZT
IVr6GS9bo4YcZTLs6QfdzMeJSFNx0wINE4lGI6jHRoCbfMyLMQjggtn0OLyHtQ3mpiDudCdNrW3Y
T/JQHAD3JEuoAhVgQhKXWLCQSLeIp9zxJAJUNJqTZvJO6NCNcSpikHpzDyc42zwmtp8RIarCtXiZ
BTadT7okkCGU4Ofcec9ejwJQk0kt0hah2dM9yiwF6OVLyV9Hx+624ubEwl5ah8Dzkucgs8x89PRB
CbYlIo1l5wl1wurIHeOph5EYSmnwOux/0zCAAKKFiIBS3C0NO8ruOs5AuJlZ0Okef1qLRbakW5Pu
VAiiPhtM7EYo3uQwOnOjDZuG/qzlj+/Sb8ebxJzdLp44cZ8hCAKTKCravP/okA1Og4KeCD2VHI84
5mA2db71msmz2+8mB+YynBvayvYHQCqdjRpI7+NMf3f6Ka0W+mG43f1/m/Af3533c0KpZBo0Xl6l
Fxl1+F3bT6Ke+lj5UNSBCW6q3nZ4XWQphh+nMiU65ue/oV0d9Gipt8ekVqj9unZkda1mgxgWNXWF
Z8CvcQvT/Mft9oTF/KKZ/Q7lOGUNvzcN2osgAYgV0FXEmVD/QuaJQGWTYv1W0gs97m4/owMe6oyP
029wghUn/8EkyJGH7fcXOv+xu3tAwkKROn5+EnbxseAZHL7jnUl1yOeFtbrE0G3ag+9Nnr+NqdJ+
Zl80h/FDI4WrSOnW4d/IgQ7VRyRmUk6gppjdU4bcnBfJZPKgTwaVrCG4kmvC8Wi9iEV7YbQADZYU
zJzJ1Oq4GA9Jkym+yYWYVeYe1T7bD14IZ0OjbDdV8Jjx9u6nM8VtkQ+g/o1Sdx5NdJVfxn3ktjtx
pxoJl7LzqigqlHsADoyw4Rq1Mn0bydFBBdnTKFvHraF+8NWak5JllB2aYruPtuPqOtxV+/O4GtEY
VPLk+d4GW4nogB+krj4g67BSgGYe7G97iapc65vUsE0HL9HOpEJNsyqsdEC4wVaOvnNITyitjvuY
7YIplqBMwk736ym2pqb0FIAQwjdZqSwGF4LrA1qmCS5ZNjYEVFPJ7/R1vLqbjmH9XAkAFCsSq+C1
zIy77Uw/etwDoP/qJFnPDEuFrifa19+M3lr0jqBe/8IQgOwDPWgpybMFi9Nt2+Z/iSwmvSZqAZCq
IGj4tS8DRJR9QNpjFG2L6ljCM7VknoFVS1U095C51ERD48J5RCgFBAkXVWzC4zdBOMHSqU9lXqIY
ypusVDvBHmIy+2xVcU1uZ7vz5wAQ0dI2qAfjMlcWKU4c9wBZzcAvxUnVGIziWOucfYGczpEmBLuX
Y6Vt7ou2AG/pQq0YFlqte5gw2Bm3iGwbCFNKId5JfJT1X8AQxNsrZvZtQIr+cEPiyrAmfyx5nTYR
FZIEtPz41ZxakkgguGVzOH1In0Ch5AekQAhc8H4sRV/M/C4mxrnf4gZKwuimf6Zn/qAXbjvA7S+c
u9bVt9WcOCsUUnPGC49DUWTny1Vm3w3XJ0kUwYPy6O7yu39vqg9TsGE79d+CCY31/LBRFegfb3OM
pnoesTVQ2gI+ADgoIZ3G5H/YG2S5+RkZtmSBf79T1Ig2wNrxHPyV3GhICCpCu2Lwi92FakbO5Fut
qoQA/8F0FFvTZ7q9MjtueV3d5NBiehwOfVvOI6aeGYuDhFWhcagNtoVxdkc6f59K/HTvs8WuZQ72
y/Lr5VzbmQuZoUAq3EH8FnKzFfjB+BUGoRBGM99xcCJsQAGD0g/KgT1JSQMARlIy3kI4Cnf9RKkz
FK6wcrSSy9nf1/OZEBQovs8z36+w034HFWVpYw5P/ZJtDMdHqsCerO1fov3HH//tAd1Qk5q3iqMT
CWXxujYpLDoGV95xxCyrKQEVTzuiKSBdD4r/cSQ8OiacQCmMngS6PTQzV34ZRbJYu7rN5SVEUiFV
OCOgu66esNxKSDYr5IaIdWBKUgRDlcnRjTiA152QEwPOIgNJbY26lF4tEM8Bp9GzJdlHyyrt4fG0
jp5UxFZ27ZMFB2ugGc/tYNwTQ6SM4UrUNnM/JwvTCkQKggk6m7DaLXjEcAY5MkIah2YB+dpgq+Wq
GMOEdfDCtR42po0X9aFfLqgXdqwvgz+T/0J01Jj/IlSn8vURUTDk9nIp+42Rqv8PFTlsY/4kAGSX
PxRBDmIrDoKuH9Ef5x6AOgyBER/0VcjLF7pvWamcl0X7qFfQTQBUE9JUpsDC2bCcKCBdXNYe9nVb
ZykIltsX2QRRzvqkeYuBU9jmVeWhu7zt6l5jkT37fOgT7h33jvOlwaIt5zyeQfTV6kYGo0NIMZY7
fKWXKQdTTpPb/pi2qQUvXlJ9PeArjgOphbxrn8JhgLPrMLWj73IGCIuI3lt1dWKT78Z6kLe7OCtc
1XPrJHMC92L0bEa4hNT+ZNvq5XS7Dc26FNOVcct/ZBbLkRNvJrsWM7ZUIriJdsneDcv2i8Q+PCLh
D7tBnKvLnAM2jtsXfGl+l0gmr8Eq0vaEnXsaNutmZDR+lO7Nx2Dy/fUL7s5UzqT4gA9tnzv4Zfmj
JWyguHfFxb6KmK8Pk3JKu8X6VEA45IyTyw/xug8kj5Fx8YLG6udbPyje4XelbjcxS9/eLrIj+/yf
8xooRM0LTs7rhT6X0Px8EgWzNlmneduKDgRGlVwEegqyhzTB17TWZROT5GdAro2Ld8u7H/HU5Vha
h7NwflbANqxoPlpbJyUcdbrMf5H5TPW82bbpvSgT2Zq76q/ER8hCiIVmR72SYbVT47bE2mP/dnmb
e6YGRLPJk6JVTkaqiNt+ygmWt+aTfsWcRumYz+FME1VoExlNaKDqEnft0Rc0EpQqah+uyp75CRWv
5lZX+reLCCDqBEKTTQPQIf3C5UhNcDyR79rrbKxjbipwiRu5NoyEO1k6wjHRc5VU9xNXV1qaX0WX
FbtrhoqHsWgI+yh4KOvdk2MsslWKjEqZp1+JJomXwztJn9M/rrDWZVxc7XbH1klrI7pFwsr8i9L6
28BFcJoBUDIk39ey3RAeZhbfdf5q00RbvBy92T81Di90UJzDhO23LfI+kwPX5kXGdHOUOjkdtzK3
Co+Mu6bRwXUjbQEzUU4gsilZFRCLu2Hb0kd4dt4BPV3j/avDGO2+P7klBUYTKkB+TAAUVoawaTw3
1zNAq1kecdbOgAtF9/weD6T8HcmdUwQp3iP0NjyCZZeE0krljUwf30KtXZVKJhXxgSdqVyxFPodq
Hy1ns2/isTtUlpyTdjT1+QLVEjlEvmb+w9miJUsxzv6d1YubgQsf6IrvauRMsJ7ctC2z0HPo7nsE
Lf6dc4HqZRGcd7k2vm2bE1otYNMmdx8y7Yl8A+IfB7OpZKmKQj3QsrH5fST7d0ykPJC0/peSI9d1
zCERJcUhWRsmNfu1RWDLIPluS5LVLXc9hjKo0wYY5Z8hOKwN+EyWjFMWI+Ci5UwtyD6x4UN51yE1
+i1irejBU475i+TKSs0b11krnUN3CEpE+RpmzezLRnEangrhTcdoCBvMyqriI5ptoUt+s3dyCFOK
uNfzAzEggDjmis5DTe9zNLmF0bzfTJqesUdc2Ok0GMyQiL74eYLqtfBLS2YekIyYPjLOhO4mviPG
JqF6rq/deuXJIhz9NmIwWDSj3enBGmaPnWXFSpyPGcyDGWqcs/+a1GnEJDH722onF45jAUXonUQV
RFVRs3scX8WOl06ZceUcVAlpCb30BTC0XreOvXqD69FO2aEeyIMO0TtCxIIqsBGQ493ngZHczQo5
tkY4gZsp0h/989+/2vT35hstRYPo7MHP+OWOZrrdlW1BXJXDJXVNlR4uFooUSQ+3RYAtJD0Bps/i
hWrbe6G7uNL0GPGIKmPeyvIcQVWZIvdCtrbCvNnOYxxexn8mfkyyrDI8+GqTSmLLDa+dHdNYc5nr
tMBpbqoXzurakH5/XHc0TyOffbbceagmSdZSznSPxtd/n59SAPVGlMB+2m4fIoCWRyDzSDGapAvb
/HwTXt6rJeDULyeeRKiXrKkIwLZwbzbZc2r+f1c2uMMkE9Tw2Lqbl4XcnjwL9g/vmIxVzYjsLeva
PTeV/7/N1wfZDZjbeG2673WHRjEbRxKv07i0fDyuH2IHXSOIu0+KzD3xZeMv/+iYPtkUxag344ZR
cuok7MaQdQr2VbURMxM88/i1tD3t4ojk1Ggut0CqJN/WUDPKPAWldfxx7BLJle4IN+QCz3ccJJZl
tkCX5ji8Wsg0X8tvCGXO6yJY6o/Pm8qFNg4/y4lw6TTwG1u9FBdTArXZ10FcNl1/7WPMLJQO6kBK
5NvCSYsYE6PFRa7UtQBvfPC69uiF4CayMYsDO42ofunXVgN3g7HBjoXf7lup/sBZfaOUcyZef8pt
l23pxEPnDW0CjDwGG1eW9OAfkCRbPcgsEsCuuFE2bZLdTGBKzQpEtdcESyTnFXprwJVrbJYAL2UQ
GzltMEncvyTTWw0h0+vqj9oVmDfclWDSLKxQfztVVoEw11dzT/qxYxg85tvAxVJiirxnhR1LhXVH
A3emO/5xdcdga1JWin/u+wOna2olcXCOae51UJIKtYnL0DHdoXYS+dRygjR5nT1JF2rpFS9tl7K3
ugN5rgRL+/aZpuseURSpGg0+npscxvedqZ1wxOClr+Wb0MBUyMDJrltHEKe3UARTtq7jee5IMbsp
VCJQ1gSnwBUUIshvANIH8ROa0+Ou/vcFUhQj1Oh+UnBEQyxekoWk8Iz5vA1AcN08kcfYK0oqK+Lz
wfFTPYGXrQSXruVfaSQy/okTFmBFnUEane6KtvMhOw9G5LwJ5nZD1LIP/1r+J82eZVjDlvhoQ4P4
DaE7T/adxT+49ULXoWsN10/YqiuJiJZDxK7nOj5VxztTYSh4pezfYEf2iw0+AQyQDi0R910wARNU
tkmIXoEXazvo1fAZrwOXbnyEvSJNcu+mgHoro3JXTayHCDI2C6ApBMNuso2aBVZTZ9Y8mY9el7fp
+yGGSE+1D7Tiz5Jvx1uuFkPTR/Fjej4jJR9H8Iryt+RufT22n+2kutWgMaVTQdDqGVjwmJU8ODg4
TRBjrnspLkjLkysMPoHRxFEc1uBhSeoEW6WFe6To6i4Augujlby/K35pMWke2PzQd3WkJ9oh9pMJ
+hTcQQ8gVBP9R99Zdav78wCyhUkJu9r2yzkXV3ta7wqvA6rP6XGIEQJFngSkxThkfBsTkJcZc5a9
tM+CCuc9KOADY3eZvE7Afi960/nBWzXyo2iSKastsLMOLdT35/WtbYDc8t1bMg+F51tHexECvfK5
nuwPAF0HjBIvcFwO8tqGRSpduxAnuh0+RuNiRCrbWYwI5dcKXp9+Kvm9M86r/vtjOZmlZ9iLDVlw
1Wecs4kyEW2Trx2xIdym/sskjnKvuZ1eiinbYgf1FKzCRkZREahTOo1u+yUadjBJZ3FKzS3MTB0h
ZADZMyiyNLVZXZbG5uDM+l99qd89A/eYAY4np3Nh+KTqt69HKkZ5EplDUcpWEb421F7D9WuZkw+k
czIiKrRRXh5ODBCyeAclsc3V4OGLYwVj/R8SRG2E4GDLsQ9xHk/LzJPN7KYJh0ZhqpOhqpzMhTer
nVOetha5y1mrKmjHgRVVZOXZGWFkl436dpydVoC3qSZhvyxLRvin/Y4gucZnZtfNtpiu30B4lBMR
k9jc42LMAFM1ndl9Y65z2NAQLP5vcCYNNiAJxF7uX6ZkWz6EN7i/+Kuw57GyFaKO0mOlH/lTmTjG
R3XdI5KYfr8nnFjda0++JxARuG6t5FxaG1UhAbQ8i5ujGK3fqDahq8ahJBgaX3k+lOdBHy4Cp9ko
SgXFmR82yn5LZTyTfFdl59Udk8I99h6FFtJAZhSYIx4YCX5rVMWValufckOIOcrqyv45e1lf6reV
ojeGZGqdMQctV5eHQVYy44owS7KMI/ONLvf5xS+gHSOCjhX6MUKOEiVu0rV66Fa+COo+75eBVA0Z
k9KH+ieVwC9DaGwGqJPpdMwV+qElJHaKpwP3hT5Jkq634ImW0tF9VbrL/ioskrx1N6hSchNaoLDi
S/KZt3PrpnRONyXHKoM/YUGALlvugbsOuUw6UNRZnfN9pgEq1A1ntjhzHdhUcT95yEhO2ixKeRRj
0IvX1+Dyc7RinrGxIvmoNBiuPWclOi+FDrXqtdMEeLdXIx7SVuplwwyEeZH7s3FVnE2EFAureVS4
zimsKdVyWx+mZQHA7TQ4rBK49qTuXTVUiqmr8tr8jJRrqJf3A3RRi1I1cTtmtXCJb8uatLM7oHAB
3mnpJWLAqqGYuPu/p1bq+gHYaGQyXcHp2uvVxJt9wESQ3MeWhkVexPEbDq2omXF5gG/dpPvDUrsH
Lgy0tFiaQNFD63Z+1l8hb4NkNyJPE8xEaATpA8ITRJZx6mbx52R25TRusBMHX/vXRZjgE++Mu0UJ
cHB+RQ31mIuTKBqRvgVeA31M/b7MgiJ9zuHDUM8rdbslaM2hkrAtUYOIHXV6nq5CcWXA41/bCw/j
yOtLgs/vUHuZz2zLIJGTpsv7FtvRUcp759Y1u8RLJRZZqw2EzTRUXE41B5c1F8DGH63sJk3KMH0a
2ShTggsZt8Sg20Tlpm2tVRGSIRrTakjo9ckIrQqygwxVyugFWAVyRoCrPnEEGUCJ/1bvdUsTIyGf
PBIZbrtP1r0FMD9D49osWNdvSd8vblNyDcnyXRVBQe9xzU5r9D1rjCkYavfjiU7m8hiLCDoUU5tO
sxWybk/iAwERMkIH71rvMuAlgdKOzwFITFxu1GZt67wpamHd7OxPYuZnfNNoHfblq0VESmyPBGjJ
kh6VDwW9h7mCigH0R6tKJFJMGTvSdGQQgg/uomyweqIQNmIo0zulfsc3VJ4q1PlHrrSzgPS043qK
owgfYrhQLxK2QpduH2dd+wcUg+SdCdV2k9k0/CoFCYT5z/gVYgqe9ZW1gUVw1E3wa1z/9F9mH+4h
t1pLfrEdH24B6zZGXm3n0sniAsifFOhiDcCE2YrG60Sd7Ne90SwwpwmgKV6qr9C44ZW7EaFZkRnk
2n0ka+oJWQl4h41vDKkwJFDleZsLebMgSHNALST9SdTeLKYud7MecxSreXdWpC56UDbRyzYmXvn/
fSwqkb0DvcMMt62dx7qA63SVuc4LT1BT/6XjeFBBaL5mfizP6KTClLBJesb9UxmdK+HewNkfiZXT
/nyD4E9/b6tjoSakHi9n6CRb8auC5YQQIa6FnPCjNcf7MuaIGNYnCZwS3HFwuSdsEGHQLqilqRT0
4CvEujJR12zSnr54gUgRjmPppfv12iIH96Ozylw0xsNP1bgxneCzBtIR0WlUHh1Q7tmPvcOBEboz
vmX65Nn24M5VSd/xIkJcMijYrNrquobDs0i0xlujwEwBUIjkPkjrLxjqub3uXX5hh568ezEuf+v3
1nb2UNCWb9laq5YQC2+aClUsCA+ljzIW4D9bkdsVJoCnUHmBDL18X21WZqK0mcWvs6Dz+phqfl79
ePnjXN1LyAaxuI0G96CMSqrhrtw7F/EiPNG4/5R33W74S56+rcSY0q+OxsegooKn9PD1Ma4pcvD4
k7i4s09VI7e4BUSzaEe36QICnWwXuLRC6hsPjk0Pb9yl5Mkhp1ttGDZXToVKDBPgWq8fCm24b1XS
aP40FvId8XdDi7NcfLPu3dcwSLBKyrl9u1NE/TZ9hrc8GuRpyIWDcHAE1SYPZzTmb6dxEH2JtCdE
ZC4/bd6Y3y+xraASfzpe2jT8BW133AtQ/oWfCoPCXtez8nje/cO+JqQmYnjuYbVaDPNsBXq5yxT1
fgnZpjZxo4u0g2ulzlpZ8498F9DgFcWdk5K/lqu9DKyIAx0lSUsmofUol/eFpOXk7TlxD1Tqehzn
pX30PgaapnY8gMxk+wAKCyurtWE/1TemAUkFpY5v6Vlyhk07alomZUGXE2aKjO3/bY7xym1+XeZx
1JURSzYE0zo+DxTSH6NWcfNh7jDKacO5pWg5iwoUFYUNYZZlg7/yuyiO2zMGbbZJGoE3Re9WPomX
qZv5HaaIpn1AKOdZ0RL9idjo30m8xjl80MjRXmKKPSEYlzPUHz7Em7PB4a2r6XKwry72uB4kAB4Z
pNS88pqSerTvMObzf4gR4ZPaRlJqswxAXD3M03QCmvzAa/WM9o6qiwu/FK8ZA5rKV8lFMBdRBSAv
iVkiZRVtPCbhr9rD4h9hUEkdNz6DlkQvFBkhRJ9WdepdMOhyP8NetgfYEcBp7hoJ/epoOQzmlMfY
p2NX0vDde+QrRJk5ub2HpIdF0zJfK4p5/PugvdmnEYS0zFQUT/4z4PIatG/T9ZiVudWNG20dG24g
fplQ8QITLl4MZPYfAUkN0EYEkiRBhiZxT3tP8RMtB5EM9r14ofmUSfzJggkaVB65vcGzInoyCRyf
XWOEhCde6MZyeJGw9hGTk9/pNE6vdw9BJkUB7xQac2ezBI1fNQJAc5KeAZVWYhZW2dXPG0fphnRp
r2gpo4/WIO4JZU3Rrj1pIeKVj3UohVnldzPd5e1gBMp7bpqzLYxMcFC19H5ItykPbA9VvEWsm4xH
PcNn34serhf+zD6ZW2heErJDFd72CpFoLPkSsqO8Vv5H82LkVQuTeC3liDTmSPV0p8h4nLf7uhTK
U5iO/07jSXvGBRnU9/DZii/5pMD53SGiDoTUTHbfnfi/zUwdmJE7ddppiOvhyfZZik+v0C0Y5tub
Wjooez8rJNKw8ceIqioKipFAvrbKA1xH0K2f5f0LZIixbcxrbHXQzDMrwWfNgh4C0dWaZOjni9SJ
1E9yU4zf9CizdP2odHfZJxeWERx/qvAOourU/eVqs0icp0hJ1oVGOW+5hW91F24hxygznI4+Sma9
i7rnu6eyDATkoSVIGp18MIsiZCQON6YHDm1dyGHiNNvVzoFAEH043wjxh46SPixdJMvmByOkPGnB
b7QFDyI3+I1ylZTpN2/R2Up2NQ7n3v3qGxlcbXDkRRnQASfHcem2pqpNHDtHcS1vBWs4PevQopDl
fr1Y1diZl26oejJnTbLlQJD1dHoQaI/uxKzh6cHgLNEw7ANPbAdtT987WJNGtoKVqgWxOB6ekDB9
vxzLB+Oon1vN1LDn5MRIvJLLTTgYIyJqaweyrc2xAwdZPHLElgHkeN+bowVh23EkpSjLf9W+alg+
Yypl6kimKF75cPFMgSOFR8rjiLAg6C7a/UcDUgAsbEc6btPr8+m7RHBCQy1FSV/8dmuY+WqOH+wk
g72nTMX5LXs5ce18gg9HHntOy+pgzX6OcBhtzlXbuJHL8cXeWt2gAkDEfX7yIezfawxl9iYXwCxN
6kQcRkbIn/dRqPuZ0qyYoNw4uPr69VjokVizp/y3A4j6PyM4n1BivnUP+XMgmzASJekE9DFRiYDt
Jom4XTf6QYkWCgREsEvKqRjP0KkRokHHmU27ohGQpdfcIMRrY0OCJMdCHTAQMRIEi6Ngh4bovZrB
Wz9hbNFk3BkK7cksElCYiSiZY+TmXkQuLtZi+mBpM4LrnOhbLPa67TZxw1wE3Dl62z+bFkjeE4l8
k5ipnFvZF4iKe8AoDwyonjqImyynE8OAUzaTmg+8RMESGqX8qWZT8uBcDvB7QkuWTC8ycifKzs4U
h7upvaIOS7ZslhWWC4S6Rwbd/alXzmrRgjGQcu2RIaN5NAotYczEmydfrUJRpAdusu060UUubWxY
mz0SMb4fQkwnbg4EheIozpic9sCw6IHRPDoFPSscBzl5CcI1teP+hkco+63FSKqonZNULTaRqS6O
SjNDgTpIrNDieQexC39D3K7mrFg0XAA1ytw5cYNOYXp/42543VXFwPM91ItrMs3Btr+d5am7waeq
dkwkJU5j94pcGhWua//9N18h1xFERjtepHWEDc/4w7rGMP9LtHKv2KYkDEvVosJ+5HYtjsZNZqnH
htlPJCTywEg+ptq7JTf4pNP7Rkg8kIRSpo0VrT+Nf5xr/IVn/C3MCUT6XcRaIW62+RRmDz7UGvMm
4b/OAWJBQdlKmMMpSTSjG4OomAkFK8C31UIWUfKpOlCTznPB0SJdCo7NBR96BIn4JOMhi38kpGM/
QSo9a8cMutSzaJPt5b1BIp6FB2UVOcce8QWiBycon1mCgxmIg24Wsf14q8VrKur5L/+0Tlax2cZL
vKeh5ciczqUfRwQIHrQJ5EEwSIhUaLEKs+Xl1/uJNEb6CpUV7jLWudd7f6bHfXM04A4fwviMFK7t
kO1sOn4w54dc18HqB2g7hPX1ipZ6LlRKN30KxSxphdSqIBBf0Gfa5hHJ1Ph/hbPw4QNq0HHtScCM
wj+hBUxShq73hEcwF9aLrzvysD9lHFapI0OJVr/k0MZjKQR9P2q5AuSt0++SFigth5OTobeI2SlD
bUI39NrMKfJNfSahjr5t+RXoHRvDIXD/VXenPvSEHwnBUyKEwxPIx9Rz+9zFDY6bP9LQaf/3NcB0
77up5gB7howcYJx4LALpmQeMf7iLVx/yE236Z66fKOx3b9dkBp7DS+74vOcIf9Yke2gVLFM3KWu+
FiFlPfsWnWXlY78QU7Mzo8ag5NwrK79PRIwoekHBA5iVNsCDcuxbaFtCyn7cjW4YuQDW7iS9U04O
8W89OtY5hpjw9lbgFiIQfCWYd9e7G0JHTNd3WXLjWvGF9HJUeJG26TZ5GBYu26QaopnuNuGBU6P7
GRW4aveJDxMdhNwapcravJnu6KQ8IU+W81QqRA36DI7WdqnWk/0tty3gXghsQU1QWOysX+aRIZer
o3B5RbruA2tYaEGt5OatTTp6XNm1E1i5GYa02OJz6Rts+B9ixsy+k+xeBVDQrM/t09pgkX+0NSqb
xxwSaHWFjj4lXbHf6pjbPzp1Dl+EjVkbDKFmE920nvQgUvImvBz+roYrxxhmGfQCj2DbotYgEIYf
CyZ9vBzThlXV7Y4JmPUr8/3A65gVoLoT/NwX0X44q0Ei3dDSeUDz0iq7IXichmolAI7mFf4HSX3D
UCkHwbGi8b1OTehOcgMvhNCQGzuErIHHyGEEj+/pJPBWIxx4NXi4a5C/bpjKgUaoUnsmjKBnc4LA
SXW4+en5Wqh+HEC7R2JWlWJAMP+gvwT7L8WIiGOgLy/YBH5HsYgikpBxFxfqV18qJ2QUEHEf0ruV
qTTffyhn+zRQZNyxu7V3WRYarSfzVX+WkZwGV47riNvXC//bXzCX7BE8q21kC8YhRMtN4FXV1zgd
sX4vLSglL3NDf5BXTIhH8zhBtlVhRunfL1xvomWgujfrY7Ndxa8RFLWXC+bItSVfcPqeQ2mYCSU8
RufbSJEqDCXNTYl/m98kkPlf2bPJnN6IenxTquq4sglM8k7K0OdTY9OwwB1O0VOpJhQMNtrPZdiq
D9/arMpkQYacG4qZ/DG2my0EdtIlTt9FLVXqkourazoZSbr6/XnoxImlZLZjVD9Sl6HuFC/taU5y
zTfQktJNNn5T/vtOC2hEoSwdtNlk2SfJKd3AXeRF3JTkq/wPjIblNy3bEdIT/UPfAdWxscjE6r0E
M7sysG7wLlREt9uR0j/gzU3EhkTsdBZ82JIKkLB4m20tf4uT4LWwCObCw5CRH88lFIKm4W1gyXwY
+FVsYpa4W9Gmep/TiMu+DM4Uq+2N+Ujk5pKdmfSeBgOXWtGdG6g53/M1Q6XNIWoqP1VvNrzcn5M3
q9ghUeGkgCeCVeXjootX+xLtsmh0DdvuQUsfWz5tbJtApetNpzgi8elf2KkTnQvE4jL/8ErVRYNd
c1U+Q8gzsgrIomVT7UGlv0j0OQjQuDz8nTau/23oB4DjmzTpA3TDwAFRK6J7jeEayqCv5Cv7vC1G
ns4CvkMYbkpDQooesXHwn6AvHjdYmbEvvVy9U/sAdTNQRhG1XpYnHpjMGcZcRjOyrq4bxGUHTYwZ
S79QhaMC6F66QWHlhn/ZjX9pZFNNep4OhQ8bkElnZ7o56AElCmFQajaJDnNRfLPRzKQohgu37x/o
5tpMss9a5WOsQK6kRcCb8FmaIlstySSS6NZxyjPt8wbxu68LvDMqIKjY8dfgHevWA1GtMAlnwehR
TBh/IA4NExi0Hau5OwfhOc2jkisz84WXSJ/9M9nWFSGVFFB77i9qfekqXhEDzNGsUa+NiVU11qb+
qLqFysgPGQ0uSbo2my6oqv1fnxiJuEDUC9FxEw27cTrGCBPxxZtAPDSRK6CD8Yt200iZalZ1YbDG
vBKi/+ExYvTxY41MSyaLaGiY1rTYe0mHnf+4w2CHiei9VEbKVu2ZvKaaYkepV/JOtTt+U2SYh6tT
2USjy+PVESHn17pmbho8Kj7nbjLcx7rLRYyR3Nx6D9GZ+Rw/KSQFw3StR+6L1PtfQDJfCBGwfj5b
MGWsxocXXSbFJAgNDBqwQg+1gQCnGRJTr6wYkLz42r+V+RaC+W+KDGHq4CDiG6TGst5e/4JfUUUV
40ngF8STr04qRJTxQqpL/dFXh2YjoNOnJzYnX4umD84dZzLFQF227A7NT0jopDh/JoJ6cHrdmKO6
Jyxjnon6nzMKZmcvYfKfEllwaDN29ZgTbNZzZmwJPzzLHPW7E9dUS4JHk5XSJbVJi3KUfxrx+f3q
T6+nfeEOuhGulisCyV12lk/H/WQ9HpID/nHNo3b2YfNX0r4Fj65+a4g7BLWcklSrDiuLUzn6dZG1
LalYq+mycnLO4QVciDSyrSdAC6/GOykC/DiGpkSrFnZG24dG54qqml7YtDiGvUhEaED+ajZCIJQ6
hzwK7mjw7yy4jTKabJMkUbOqH4IewyndM1maxIYdrLKMAcg/2z0J9tmZyBEwFNGkMO6KyW8l+dAy
8w1v1blWF9ZE3vM7RF0O7+LG3T6FWP5J+jRwRaNUjOtZsfKwlOCz4JdFozcfMgAzhqbrXfSgSyED
6xV4XnKh/z6JFcyG7iuAjcxFoO09iuhYL1i6qWIi1IM/JTjY27Iy+FzCKshiVKMHTzyroaTiS29p
IJYV2fwotgHBhkc5bzW2q8bRRrYT7tpAXX69QU1lBzPcYs4Tj49g8CiYNZOb5g0jhUM0fGvOcJVX
/Lcx8jGXpirDSswIQEakDCYBAzJcj9LKAQ53Li9lQz1sp9oXbUjbkWAbLLOFKMF05u5iHa64UdnJ
ab6acaIwVx5HrKuI2cegCZuXyhKevVUc/z6kCZZ5wbfo0ozKm6hpCLBAWAAiQxJ51kmw10m5PVtl
zjYaz8Wc1bvBK9BOl3nNLOwyBk4XfcC5KtIugdVgcJ9S98zA4Ds5N27Tm2xeVTWGomnmAt+IXxSN
9pM1iRupl8XmYNwI4hmmeNHPgGAo5exWE6xHPaQBgWrgxTobrLzSrpb0AjZTdyooLaU6D4NOpmeh
VBrAls1k+S+cK1hw0XnTfBjubE0W2pU2BRM6O8SsiDhhZM8aSGKxbXIn+yamTGXtT3dvjQHk+2dw
ryU96M8RGMrtWFlC3+QKGuyXtcAN8ysmRFkZZ7jM8K4LZvyYYoLobjNrkCfgCOpNLnOqK2x4MJaT
2u2JdyAe2MZbbx7eP732i89JDveG7FIvlvH37WocaDq0VBjQP+nN4ECklE84rXtYyUHD4dE0nOG+
423ws9I8Hu7/qg8J2F/p0TFuAk7dYwjxdI/Rwpruq8dQWLLNVIu9zff+qLWr9r30iJtPdzhva2Bt
cLS/bVp5klqtmOXlILwb23XBzMnNlYGn7OtihLCSdyiSJ1wrCU9g9HyxoDXreGSfDHy5UiqvLqEi
rF/auFvg7Mg5nOyHM1E2vm/n5SOvaFzVLpeO2ezS7jlvjjvFMfwKKfPmRRf0CjZqUJ2r2Zo3niEL
oP0AI5LOYGsSwcMnmH2ecJjj9QldLx9WKPS1lIdK6JYAYGRg5bJy/qMBWqLW05hRZK/CgcD82zkG
y3GUj2zMrniVqc5OdTndYcXbLSZPOsSXuEeyxg26rL1U+EMcZjC+e/ic7v5Yjeg5wgZmeruL25aw
9cP4fz8K98bTuPY3GtIm2qs+vMUXDyVfCN27Q+xQ0PkZwOqWAeBqgOI+Pci1NR+RyEVeTJ4YD2II
9zYfRGmiGxlzKg4+BjN4t/Im/y3Y6yA2MMVhVWm4R9d8i0CkeUrsXSsPtirGimmBIjWl4v1hMfuT
U2Rflia8vd+wZdgdnM2F8jjLBb3sn9Wt2BEG3+4qFFD6hhr9qcFYmVp590JX4XQTsudyzy/n3RyU
j1d0Weebu7orojw/fStLhLL0v1CairUHDH7IpR1xCAX0pMcrpc25LFoeUj+IbXErLobC3jMYSux1
hqah66Vd+yj/gHvqXMUumlTorp7cgEv3999TjkqGRGH2kcuV6F/ie2u10zneE1EnnGbFeomQgDmf
03dKLUt9J8HLvTQ9ydORFe+HYMPnH5YIYoWbukrHr61tLT15juDHdqTJlAhRwWSfDlD8LNH6CZPL
HHersQzQBwRJBQTnyk/0DnQFhZXmQXHri/InmwX/9H7La6ufH6rl7phEUMJirYDCJGYHvPQFgjBU
iRRaGXuhNmDOb+u8XshlTLk0aTY/2kEQFBql9UmhppDZR7SZXTdD+QTmLEwaKdWZ3mZflRbz8gQo
/lwsGq+LO3vxXs/kaEy7vZ7ep0auBJ55GJh5HIUOSutlUbfaGN+g3wHknwjOfyThzlVOwIE0c+9u
7SMf9rZVaTULO1xUWzG4dzuI9L0mg6JVSEOEunIXW57452B0qW4t45E4C2rDgSfTgT/Co0Q3qHTA
oJiUmRfEUSS/2oQwCSAJ9gmiGGlYC296t+V3zp6TfKHWoqMa+QsB/SgN3GFu0y0v6TA6WakA/kus
EfXHHg1X5X3c9omtJhSLYyrL3krokNtEq28Z6sjp9jUIVp6huMa/8NuSaXGBZZzFEtLosHETCeUs
KK50hjkqTTUJc0YwxCV9NDqg4WyklRCgEhvfD4EU0rqU0v8twG4s9SW4IPbYRcRyYMJMH9OkaOjf
GONgcuEzoiOuLndX0PfJ03uKUSoJdYxZspC5NE96iRP8alqeSBmkZR+I3NvMMD8qVKist5s2wewI
mGA9STwa6pmvEb/UnJb4OpjJ9g8DhA61PrflE0OF6fDhJqx0eM0NX2r6ydqv4tJQ1iPMSUdEMLfz
qflltgrBkY1QwVfqWB38JG+QAkblKDCGmiKbWrOT94dw6NJZCsvYgJEN6X0VGkHiCEptpcPqr16p
Wk0Dnc2OU8MO/Rfp5TDsUEgXKTVQhTlRdVOmG5vaX2iyzVi1kL9jTde2b53gwQGxVC6aiWWEe21q
SePS+f1iYL2+1JS3HEVgFGthHER1IDQ9syUYuAlezcdasJOiVMLikg48k6lljVGlz/L5jaH4Wlo7
Km9zafpd39UHdS0fVbCMeFW16Tae7kJnlcg5R3/jmtCuXzHPTd2sYnIv7zCNir/g5BERYPW5zIEx
Z9iDamb1Jo0Zsyn1KPfTqEzrV4VVQdvqXvyL+qMmzHnz7opZMphL2idW1x1rJi+cQzngqzlTTA9U
HPo5G+qUH69sGZyOc9BDnKbdyybe8t6rtBcXMtVcRA0Yg7PB6wiFVcJxc2HlkT751gMOS6VGseJv
3dFcRQUTPQNRUJI7RoPrrG6bav8F+i8o7xih+IZnfv9EbORVqf4ZVQ1FTREJBt66kq4ExfdpiUoS
spXrWwl305axUg8YxTeeMUcgbesD4gQdjSqTDB+l210y2TOKAwvPJsqS4aBffUcBZcOVUCM317DO
8U2PdBSMKkvGjTF9/7VlovEyKrQyN5x3I8OJcp7nB2DwsZKm4tLz/e1rXPPdsb/NF7x8onD1TwQL
q3Gr8HOyTmWavEkF1lEdjLQ47UG88Bt/Xhgf9yrkP2pB9V5hKF8cMlcB/RLQ2Qtz8Vr6ZsrlX8Qm
Ac427mbv7udIB4b6J5mXIPew3hQbB4ZTq0zIB8frnzidfcfefE0TcjIsuaZSmsFjZcz70ney/egi
5tVd+leZCLJ7MLT9w+DiCDw3lehT4gKSs6zLOBPOwcNfus4USya5wBofZXtTLb/kBPykrGTVLiKu
lU3pJHLNqsOogEftMVGutKL9eq9+Y7MgigzGJa/V6+dfaCN03a9sRNX9d6390JEIKKK8Csda4yi/
ujpnDHUoW3gIt4Wx1f8KyMQ/iP623ZCvqNxVgboNv0cFP7B7LKu/56ZGi4+4hUXd0e1ikE974RWX
m8zVKCicUrvHI+HTlPO4DA2qBuAchnSuarQpfWsCoMZ1S+iSDI2Cs1pjaJsw2UVbT+NFUTReD3zQ
CgcGfUTkwAMfCBeGYuEIb3XjuDVkojJOC84IkhAIH4Qr1iUAXKW0ZNLtNOsS8y3gtTCQzkUPJItv
os2P7u85P1oZjfGogTUvjOtknWmOxIP9H3hCl9bkeZHw77cwIZNBfwGC5KFzXlJnAdIka3xXwpy8
3Y7Eb7PqJB2AApAaVf0y/sKpGx3zT5WoxQGrfI2BrWdgAs+AMuOBG+MLx9HQu/vemS98uZyL1U/n
MjUnUYKXEB9aEc7dksVjWtP+ejNSpzL5T6wdlxnENhgkYFK20/3OMQD9S07J35r3qXIMagCZtyty
iujbI3LBSy2yWrHSnm0oATK1gUmaVUPnEWheDi3VyfznxBuJCit6gNO5V7aJA5j4IITUDYvZEfCn
6lgBhdbdkcP5/YYroFczEL99SgUptTNYTloegIk1LRHsphsEe4wcyuR0CcAOB9482M/N+oobPmC2
/4X2ArFnpZCoODNtEI04noh8OIKcMk/GoOzaitzM1xYc3s190q8D5yunOrx3d9spN3klUar3ppcX
MLgyhC8AqVUTTATup9i9GF4iwHdPYXOLWi/0pIKSn7822ztS8bCW4aEG4TlNOIOezDIbQkdAzR0f
anO5yeKjWmZWfsf/pAcXGyaTLGcEalZG4lmUGtXCsubTq3xm9q27FxFieK88ntuSnij2CohlVK0Z
qyZ+oqp8HdlBeqRLZPDYAufmJdBI/i4JigzwnEP4RE5CqspvKpo52q0T3ks2SgWnqAB2U6GQAkAt
cYqyPf29JCcicQRZ+QeLARDeMISktUPuDMWJNakspOw7/qBHSrfI4V4lTPdNmQ36YBUkby1IfHwL
iW8LMHdcYXEjS41FGrfNKj/Cyw5XlSIOs2k0ZdZdhMWXpXHHSxXjU2C4R9/Nxqbn+Wo2U1Ow9yIX
b9Y/+DYyXEwet3BbAsfZN0Av+OonJ4xLhMeJiWUWNpPToFjkDjDogjiR343lvW2PMl1i5Y6SBgBV
bELAfLvmxAXp0HGj5eeNcrDYM6s1ODUD93bCeigUmRUA3fE8zc4FKu6qkUEG2HspAById1whtXMz
J63PzwwjkUSSYr/cR/ZzesgY+T+i6XYQJMHSIOSmOr8hPextK4LCw8wcvWPGKUsEeuE21ZaYBS7/
lW1Jd8aT1Y2dkt1OUHr9cVZp2QPsCPHrhe0IDCKUHk4MlW7c0cB+VnTjsh/D8cpB7nu6+gYo4m2D
XZsikiHY2UdZjp87mgfacYQvltt9joJmjVAGSrWGeK2BhKo3OfwSD4IXS5cwJvofyI1eac23suPF
aIPtJ/gwkeme6kH+LM+/rizO7gUomeeLU2Lz2lAjeI4OEZRRWUPdwLezLpFJLKNkQTlO5rFWQ9Fw
bugkfSrzzSRVCBLCx+cKxkzCrt1TlTYyu0fhL/xzBCyZf0JfRRDU6JMcED9/+1ddAgGABtzqlafC
UnFkWDYbHGzdiClNgtWxgwU8OwJhR7Y+0Eyov9QzcuY6/G4IOr0e8Ki9wKzrw19/DFzhXkSlH3mY
OCToWNfzWJeFJOD8MhTGuvTG/XfXp/CLKiXj/R9pOrZ/FEkTU0D+azapijuaGuCXIkNmqPukPJw4
gLmKrPgKoICVEgFRXTVdclRVyK5/h61rEjheAP5+RwwXsyUqNn97JFXXlzkgBAuZ3KACRo5rdiu8
taZaq3/F48s0DL3wr5nX82UUxSseuPul3ViGGpJUo4eocU+o3GNmiAhtuliR0oMAx728TzHCbD4z
LNYIXggyK2DGothCnBUkfsRVLnSno5TX7mLmrcM3uY3g7X5oaVfwvUNpmoC871BxsbDB5bP5YsqL
VS9ntC0x7iZkmVTHTaiIM34cov+DGlS63bVCWufMLbKG1u/F1uaaAzV2fxBOVaAK8NQymdCpzycc
YF0anU7HLYcLOIfWm9M6dR8Ng6CTp9I7qd4X9pQWzNvgNqly566ruC0ST6sdxG4m+c5NMRpX7xOH
rn18HCEQ3x/9Kjj8jdd06Wq1ri+yOmxUrHEmIoAKljQ4wnH3Rk6koznhovzD0N/r++CDydKwabis
ZQIFjYPE0kd4iHbN9CqCqJabWyNVqqMg/qBsmDU14EZn4rULlyY4AWkCayWyDx3kQypgMdoJA1HH
caaWvK/4m7jnX+8BfPM9YCPvZG4XOTfveMl4/gsR2pXuTMttuxuRfVzhwlSUBd8by7yitiU6oPAX
0HTRxm/09qN2hFKffmstv7EXgLtqmDlwngvq7oVwaZjtZg8khTjseX7JDQYPu4RTPzes/rneZKab
tznykUCrcVulblF4irJBw+eALAvQLUR29KQbaaRwZbYQLh0s288IHM9lcRn5DgSHVhjZ/w9yW9P2
T8MBY/vvdklFAb8lWIc4CiuKPFSFqS2l78GMKnc9Y61jCAdh4O+76UCNKght0tCZaXsPUizAsD75
+Zn44goZggNFrv7BWuEAmtGOzjIZth6I3UrVKohb7N4ZvuXtFGOTWQJlcpcIS69+diR9DFD9pFqE
7eKWeFnJ3mU27Id1ldD+bV7TYrzo/RjpuEaSPLTgz+W8/wXfsyemCHHbPDPaTIwMoXeZ6uPvDgO1
wH4dUT+5KtVhRaYfAz64EsDU9Jc6Bmbv6q8aCDi1oC8Ed4Wkq/jAW70tBDDnafchgyEoUb9bHqeE
zSIruhFW1uBri3qh4MZQ7EyHvBOVMIT0wWDAwGCGnvpwIgnkRcCdZMgqAK8WiAdw4AL+bXWnNr9F
Vn/KEgyRfiOCVwymSQXcVC4xMeODlW5FX81HDeLsJ8sczIE6/zKDI3lFJ8jxnfg1lFkoOijAq+Me
DKej3D/YMhq66724lq0JVzY+TsmwQTHKYp9ZTCMTS3iXKVb1XLV0dzoKaLwhskKOmP7lgHIzDKpz
0XKhMggjcn5IXc4qQmlg79V/0APf3Sc8DM6pf5EuflrgXcBLei57ljJyrKnBS1yAjm9MTi1rD23g
QsZTV64iJg2pAzgxCwdfKb4U8sWddu9khl+edKONYxTd1QFQ2ZebyAwNMv5D1Vooqu+/73tgGTFW
2jMjvvLvzyg5OHy6p9OfUJyAoSHUJr3w9akz5/3scVH04QeysFURqnL10hVaNxLVINkGk0+pCgyM
R9Ps9XOQGqfawxdUw7eKbogPFjMzsej/N+/n+kt1Ug9Q4JQNzOwYuINcoJYSd4gD+yjoW1XN8wJn
djttRQ81hYropTVGWNRmmVs49MqAOVSIGp8bgJdSQzg58aI81bMRP3cBxVbdJkyB7Y/lUq+Br+Ur
eFPp/F27+PjwGJ/Z/S4T3eLsYVdiPDd4/Wi3tyqGkuW2N+M0zbKdS8kEVBat1bxKRN9lIsdUtXkV
DrOmK9nMvIYczF6olcq6WH2Ezo2WBuiaEkkhPC9f1YCBRkUisq8RuItV9Pt1gsK6THAz3I6F4xvZ
TiPZU44NoVv0U1rPcno8TpBR7027MIPXEF4EfShaHqlrsfl9zR+UXSwSk/it1UT4zryzeSJFAxYW
caLWB/76ycUTaECvFpc+Xcr7P2kNGq+V6XRTE7tDWP15/gSIgsjUoW57Iu0937N3T/dYjJZ+blJi
C2ec/KMqPyoQY+fWSHNzf5aU2RZiuXX/eGXfIa3uexc4NbWHWvZHj+g5HZeSnqSYjB5N5r2HVJj/
ur9/5/lsDVRET6B06zZDMO9jtYAzSQscmLbqhvn/DC8W9xFYEk865BBfnrd0UEOuV3V1IOGAyb47
DjExd9TIz4KbGJWZahFqCwQYR4nIIgS0FFztQNDWb9CrasByjrXU6oPl0tkY2QwE81peKHBheYd0
J0dtguo8gm1ci02WkwOmSieJI+nR70vzor9kkMYnivORWVZtg1tcPBj3R6qHPfDtlDc39XKaYHt+
qfMqujd4TwCOQ1Q0GCSuBVdnc3xcr+4+eEycPmcPAfia43/PF7V6LrM7HL474YDnDk/rxQKzsLKi
byi7a2yQXByahke3C9FCSAFgvpnojk5Qi/LrlQNrs6es4euIl0bwAd2aSfotSh85kh2srnsvdHyS
gDcmkr28na8bTKfVE3eJ+PmSVTh5ev0VgGIcBkoSwcwnaGa2qCv+0JTgP2QWQ3SwadWLF8h1mlpf
/CSeLeluNfqnAouhyW81/O35EzjCaaoV/AMDrMMVy7ci6Fto+Ux7eMjyKlW5sInSycWFSuF2OWhn
dSRMUbGNR4YIRisL6QWbWWIenF8KN2p2JU7DBe0+wJ5nJO4L29feP2+0AWyhFDnU7VX4U8hgjVYG
m2BGgaJE7UJdqfg5TdcVeDlbeUCqta/PbxnGe6mX2xBnE0qiUqkJao4gwmCDN2q7A7zRU9hsBzru
a6wP5voZIjYGd6rfQkH6yPkFSRc3BGBq+4GJdXY4eeeaFRV2jMH1XPM+tJQ2xTSr9UlpyR73f6DX
gY+B+dEVOj8jqGuR2hhB4Ov2cqFN2XsvHwHqiFPnkSwW2a1L/RXjqTbzv7J39fjxPevEGzlZ2GPQ
wP7R7qDGC04dUKIBt/uunUe2hL2vRgRrQXy+86NW1AoFRfEaV6oCQuKNvYTt4T9sOwyLfPkp4YA+
G95WEWhd0QRJhIfWMB2UGNqdq7tzER9C+FfKbiOcflqFKIz0dhRP3tLBLqqM1+YoX96lJxWdFjEX
6CXq7/kCwuczucl9gaTlUxA9WJSRSyqH2nAMLKd2wwoulrAUAY+M3xIRdez8SIKLQKuBPItkhvJJ
mZMQ3MtTFoDf5y8N/MQBvDiuBCMBZSYKeFgCpGVHh0G5p695RKoVw/WEZQ1LyAgdqTAIdZP1cqBR
VWWlse7EN3THsFusmSF4HN3A/D4SZ1FfUuMSG4vwJ1vHU2zt4ZvyggAQTOKlEkhCNVGKK01PWHJK
lon4KgA/tJMuKXmgyrGHZD8Dl3k6VTIztd7VegDczKazZdYoK/lRrmqViG7Zq4AnnjhSbUWGjTsC
M2CFLQHXYceG7+smIeoNBS2JgUK3j+J3GeFufqCoo/aGXpwqeMQvd0XB8P6CxGx+5UaN9WRaXqms
6hojJnIdCq/bzoEBZDyO5qnnpEpCeqITBFpzYZfFG9ONBcRdFCJ4Jkwpp612e3lTIFyqx41aRCWG
X/swGBS3/nSFcwDKmCDFJ4H1K5qvr3DuTANv1HCN6qvfTIjfi2dQpfuqZpqM/X2VgGCKEc+va4gA
0d2FWjyRRVvToe94oAHWQ+6EKafCjo6KJ0fgtz1UspMyl2VhujfAxNrhGda4xu/eEwgo+iOZ9y7K
PjizYQhbu17XFZ9vCGoeM4wTtCbuQUK7CeMsaDGXezDdKad6jnII+D2+cTa6idQBbVMD0HRi2V4+
qn9LtnMbjMUpklyMf+81tidvUpIecwBDV87V8GCeWGMybFrF3adZuVnSw3PEiacrwiSMcJVnw6pL
aYkbqzNaPaPqanhHkzmJOIEfSWhX4BuOc/qJVSOGZ9qQmrABOfd7ETj5rh+osGwkKSAzLUjy+s7X
S0bndrl01J8ehEqAXeU+vohD7AsG1euCtymXF7RzT945nySUTNvx4VFvOiZTAfqazH7wYvH5lkwV
lNRN0vjPhf+drR9UaeinxOYaZ4wNrzew+GNn/3pZjYN164Ez2TK2LuhZWrprQZIf8+FWWjUmRwT7
PAoVFyBdOvFhlawTCnJ9jvqVeTn69AylMl0gmsIsChmF30U5lSQcf0HHcgTsVYfSmVpDdrYBwdnl
QzCalzx8xlNX9ACnLnxih9FuPtYrRiYAgFVz0qdSGR1yjlIuFEaY0Ki1nc3YxdtldjcCUXvKNHFu
RsLwpTgRFUVCUlbkPNv6tpLpXJyuMUvto0lx7j/vrdUUWaUzL95fh5L9JypYkZRgWJlCqvDyVyTb
xR6luSyVohRx4PsYNgVDIUqIE74vl3TNF0V/T+CrPVDdDrNAw6I3LXR57Ng/BHCB/HdTBkH7/1ci
oysRrMkJdZhRT7YLH4UgzMFd6BV3Fo81PIXT3PxrFdITCUUY4AIzGQCL5KHqDFO9fyflFhpIST8r
R0ELljLPFnGM7q2REHlGFITHA26j2e5IugsW1cz4bSfwGUq31R36w5lmMiBSwCBai8AM+qRnfj8Y
O2iH40U76CGAijagbSh225gI1JKfc93bpi7GsWSKZw30ObRvKKSbaLoXoDzpam+X2ZQLwHXQnEr7
GNsQzwGNAddv1vVHzLvYwuFQvW96PlveZpD4ml752pKof9EGsqGU/MMkTzfqAGl8Oj+fCVYGUJmc
oaOT3JjBOAb1ETaiEtrNUC4QQBV4RYZdlneEgOr8dg4Is0/8sYzfvsTGxP0fdWqc+J0HmfkMBo1F
+ThYjvbvD4udItnS/HPhYvHlUEGq9nw594frYt4e8FkgUMnmA54WBsDgVchT6vHOfS/s5IBV1CvA
jzbOUuHapjVsUPND5NXLE8/7ZZHkZwVuFss14y8SHXL5cNqFnF938AFXrKCupciMdrpDfpqgS/nZ
G/3muF9zNN1bC4Ynv7XGfKFkGTMFtBVaf/2TtbrB4Kg6owfIwa4IQ8ajJMe5v1Gn1h5Ee0SUtw3d
tmP54zp6s3FCBXPWSX3R9djKJXw9wzDczHfk66HQBx+Z83t5FGV9EmIlv21JhyvBdmAmOgQxhZl8
R32c2FoDVL7oNtv0K5ISPPKs3gqOl1IvyTCaMMKrumEffiGnCGEmqXIemg0+/5p9J1dY81UzjaM4
2kCCf4iDSKrF5R8R6o9qEJYf/MQVHOmoJzzX1Rppd53pdJpLpILj9zLENvyRYmM+kEgbMlgXXY9K
yDMo9SOGGNzUqjVObMhuRWIBYab6QLh/z2AhtbHx8UcMvDiN3BkOWXZDf+e8VCOdHszFNqZJh0NW
UJf1B4iMgt8NlTnn2PMCbCBdHP/h45io8IAYeBNO9wihieaoExwaNAvBPOpGmgUs5JIqwP9MRs4i
JK+Lh0BGnHKlYk/ppVOPvGvgMpa0/ACpheKg/YE8yubLthcLTxvtpGXlpKa/Cs3nGQr/hD7msDUG
PQ1gaGj4wbvWYLnUS48BT4oBWBxFwsiJE/i6AEHTrT3sCJErmHS2V38xvGHMQ739w6bgETm00Rbk
5UO2VTjaAjNvKCxZswiEdbIROoZqjPrczpAZKzRAb/Lsj3jW87s9mxaHbchz/qxR5yGMAJcjXf2Q
alB9yaxP8PnLERM1eoptkosl4caLEpjBW+jBiWWyhqsua8dsJVHqJHuC2W3YSh0GrZJy8FUmCHrM
kXNbI8hhNzjBzLaZ3xngsfCYOAwKoVIfuIaSI+2SJoNISpWlCLXBn90RA+hqTV3a7rlGzdjxUb1R
peb3945RbSZsGSPiGf9D5jvJzHt7ZCbjIqsuW/8lPZLK/L+3SUQDuucl9YDWZsIWwpsie+1E1/+1
vRnl8mK9giOjr3VZRJOQufBpNO8uzBJ6AHsM/tXnVzM8LOEZPnIIykImDYaaTmW4NeO7ivxZmUX4
rD4PzvbJZlpY0zjDpo+kYRYYskrgAsCMcA+Y0aYA1dsfMuCFy4PXT7XPFHe5yVEFTCYwBYAJ6NOH
q3+YbWT396JNK2f7S/KMIM197BcE3b0J1o0WpZDk6hKJTF3waPZVPtUlbns+pcwnrGwGV04NFrqf
7e19qMf6J0f6K/iA3briCM6W6kvWaLvaTxmg/WnW62/twtvog5xdXrr0hsInCVdoXN6IVUC+JTm5
HPMZuyi2aJNioKCVt9LIG5qwFO/Y+hhxpYp5StxtAC60QMgLLOsSlm+gN0/cTh/IuswbEKAewT1y
IFoj8ssYLmBKwiAFwN9No1S/AtrRAtUl5Jh06CTMxUcW8Do3TwLshY5ZI9Oam0etMBhCZ2jYGUQQ
ChpaEnS8VnMcw/FvtieFXaT9qJrLQFG+1fBNnkkC+Kmlx0s4+uegKwaJ+flApd2lwy30JRLEGd+W
dmd+lnOkJRQxtqutCnQxCaioaadFTG8s7XYFcssTfe50eUlmVP7S8GwL+Fy65j1a5BNdw0F+2lZT
2L2YenD/eYCFCwaWI7EpFWw0rm0XdYB+mJrcI2QF9LfAxOHuBQa7gt9dgmjNqerRL8+gaLBYB7O3
bVc4Te49WnQZHDQQKmQ2TryqKipv74YzEl5Redswx0ofSWRrNRZsCtbh0icCHYPNRRv3sqjxlZC4
HB/lqWxowur8vD5lTteYMYf4C9VOeYTbfU1gW6E3WapTXNu5ESvFQahC11FpUsvjc5guMBG+YfQB
Qs7xEH+iRnyBld9QshnqFZdktnr1uPv0FyEmMfo1GQqmRTPSwj+XV4nV1NOnJMcxJz4cHqSXQADq
xSnYk0sjwZkS6i7meiseZHNIWF0TgTHnBMbYCYjbw/902UdRUTjSG4vIPatxJofWGZSSpFHelWyJ
W7DB4UBM38L9gtrDUgDHCTj2X49aIs9Guwf0B4wc6MQvwO2L1JWkAYzjoYnbtTNm3UjEYGeVhm5g
yG/0EPkcD86ZGXeA5Zi/7do8pqe4+8W8888Uq+1FTeghLSYTWnrhPI7WqBvbfqXL+zUPC3swzSJy
2xgnHIVSVKOdgN2Nm6sa2V3Sds+rMqxN4cYdb8nOtN5pqemC4qR0YJuYrD+1BvFkwRekf4m3eCJf
LaYFozMab3Mg+iOjxazszltxalp3fbBX6iCle/yvtdzF0FGKl4WSj8CxVW6/4/AQQ5hKx7DIPEm3
YSqPGUYeYOZZ2Yif5FkQlIZ3bVBcKfVQjrlZkKg6b4Its0jiVx+ACvFDZgEgU1VFek6LS27QgoBv
8GBfttv/o2Jjq2JhiLVpFxnEqgXfHe2Kmqmsr+CineqHEE+/fyCJuxW6y3qS6+HWDBLapgupAEE0
nlLxepnBMS9BOoP53/DZWvkAKUOPKbCYNw9qdrWyZVz0TsYHy2tTXsiKgOJhb3jz834iE7MQTg3k
UonesSe71CJMJONHmzoVT2nXalrGlnnaalct9h8GS6oOujHFekZG3CptPhw68aOUA+YHIO8g5pt2
xchY1yw2XeRRDoUP0IfbEnJIK2vzNkq9SrgLG48McJ8r/sKZ0h+rHSpMf1NUF79kV/9LorRC3zHE
zxqY41GTLA7YEZWaub2zhqKwb0bOH9pxIfM9iUJyosyP+MlfPT279jYfpH9w6O8/iMiEshk7f/KT
nnqPd3aKlZxD8zICdgBp1QaRUWqniAxL2iIH2sF7JHVb2f5yeloWsylqVPbQXYGo6wzQZqxWupmf
nXUzHRAZ7Dmwc8caqWXiIWMWeM4e27RZEGv+u/bdcMC3iP6F53v8+0/j57F8ovOCJJvwiIIZnaaT
kpQX/FZm/92b7y/reQDLDETcN9QiuZvDHoqeuSNkm+/lMY4I1AqDD5raIoqeTEmbObIuIrkyDHpN
mEiV5gPU3CnWF1ZxY7OOTLc04IfdOd8xna/QVP44du1prC6qpL3k6qOYoyUlH9l6bDXrJJRc9o39
rnlMVLfoIVDLTCb/1HhOsyvvI8Crb+Kzi4wB7eJrUhM05R9gS1/TnTWtiDvgrgK1ZnG74p4674lf
9jMN/ospclOnCQQWieOxVPANtDXCDHOEx1e5JtgHA1ELZkWs3/68IYGOrXHrTF7rk4rNPh26qFt7
PXOlR6i6GsoN9OtFvfXJL41bb8cipJkXzTiqKIl7ILDTfYydozGG8cRhQkfXlTjfekdNIiB0x8+M
Qw38VqhHP8Y8YEL1E/IXzoRLaRyWYYLjPR89ful2C4ygTax0yCb/79LgzesmyOMGpY0nsq4gIXVE
qSbh95/b6EyiWWzdpzx/IP2MmPL7+q1kdX74vBy9S0YTFwG+UIAjgluqk66O2HxYvpq/uMDT1UWc
LS8Eab63kQ656X9zTV7SgsSdPs1noxh1424WUzKV9tmVOW+nyLrF2l9TPxZamVedyz4HS9b5F4Pl
5a8fZ0YaPcbaN4QVb8xnZdyuelBLn1KY1IfbhygWt9vgmUkjFuvKYaWRpJRraaHaqR+/Qs3dXjWV
JNGYPfO46pwFWee3+7cEzZd4B5lF/8jd3JQf/6au7mV2jqp52u+xRFmztH39DZjUVat8x5XU3SQm
uW2/j/6l0XpdrNZPFsT3e9b0CT42nTVn4JbAW3R70E09+NGq0kbe8lugdGAxooFM4y2SFyxy4B6s
zSbto9FdCSKy4vhHlX7biKqPcFgwefP4pwqg3uZIomUlfFfPUktoHO0VeST/xau8aXomG+YJgtvU
N98xImuyuqTQ0Kbhn7N2XqFEe4J+aNFD4vWuf4xsFGE3jdqNg+UW8KVSX+JDczwyAHs1QVMKyrE+
THmrHAkU/mvcvs0td/HWPPb+X84V0/wG1YDKIDekLOwXvlqvkG7xJXTpcuVkfN9G8oPc8fELuzok
0n82681cNxx2Wa6sYdAYV6SYJlx7Aj5TpIs9MRRsBpVAoyni46TJARGtoCin+k5J8Mb1E0cHprGg
co/FvTM7s0hOlShT3XpmQDEvO8UdzqLiLDsmZAlPd6hLxjNIUj5VMbwT+UpsaGPlVge+jGH6poYm
G0b2GaHUPKv7oNAVu8FqV7FtK3V+f2Y6prp0BSS7nc6GtegbNASi2xD3Ak/1ZGpQsd3VoGcSxQlZ
mfaOEPxc/dwnzufpxCUwX7sZ/aNVyHrvYTE4+2U5DRvI3z1YguI+b9huICOi6Tgn2jHFQFVsYfUx
xRSIo1rNjyCRjSmouSHOuQiSnEbfCF6UXzznZDUCwPQG80MlFacIL4zwlp7wDGsSXSMb93/I1Oup
Ygu8TSKsXOnjhuYL8bqSpin9TWTEL5RGxd/9KFLoECczpEzNJjFNRE7hXcFFJPNa8CCnUkbFOw6p
mai5QfbOp0f2zIfwKVh7R97zVVpNfWjfif45rLBq8R3lfWuPuTG/D3SiJs3h12Et9TwJWoZBuNCk
Oe8ViE52bNCDrMLrKhKuXHMkR9EbnJ48uXRYV6MeX+O1h/GroJnvw7bxNvrLa1OY6H1osqZ7iD+u
KGk3ubZTTdnLvm/JjbDjhvW7jG41uVxqJjIa9PgyYUdhPbur1WSTil5g4BbXpxDzbCO3hC4eyGeO
+ZjKZaWZ5wFvop+6aJU8jSeJtV0cou8N1mCzNpJh+V5lDB+fKH57p51jmcKCsi1TEfxapXKwKW9l
BjM+OUJfR4FW3QBV7ZRqdxcRhWOrSlLDtfV3C7+mWUcgp+dXkkTeE6ugK+sHuXJ/u9XLFIBGlRec
13PF5ulM6PiVN5+Tl/m+CZkfFacxnvGwiwrsq46ZzY3VkpDrRAHNh3WqaC/bSRy3WLa18rs/P3dq
89zdIgydv++0l1J+x56ggbmwQzSYOXaSkqjrfJ1b0wV+pcUMY9KBjSVRWTLrF1rVA2KfLXn3iGmH
5/BSFGDjUccPtQmUiEb/y5hD6KKeNjWwrVGtO0BHPGTcoYwz+Bvbbt2iDzRjz0c+xUG6lXpup8V+
djg83dZzYX8esfi4ndN5DCLvpT0UlYrr5SgYQkJxciAbdC7H0v0fMGNoSybaLIH8lCmuFqS4Yi8p
N9wYAk9zWvSzT8itbicmOq0cXHcyp6nmKeL5fMfEd0Vf0ZzJBWSD/n55/oQoESsuo6rXbCGQNlUs
5C21U0AHvJjq8iA5QcdSuKqjrhO8T/IrxgtTah3J+qesq+aHA2L25gW6Ewel99CLMXFBIuP2oXVC
iREoRtm3aK/F3Hi3ZRNg9rRazZwFvMHFlyHk3mwAQJnBWILQkQHOCXjvAOazz8cTAt0DGw222FJd
+GskkXnBHah6pfu7y3csS19qeiqQLDWCLiR077NpXw81z0tjJuxy09jd2bqV5e4hftKFczF33Qrn
N5npLOSq4tIWsIR2+iv6ScRUCjDI9eNXPEWf2GOPkCS6QxXuZ/Y1cFa0Bsavaf5Z3ds7DeaDc56m
PYMvltz/86vKGxdc5DbJmYNFc28XE7AiTVFKZMBf1GG+t0jCg2agxycM3stLqUmus7kBGMKyi1ED
8RbjlX91z/XHJpD4LLhUI8M7mbb92TcYckxpkx0GcboS2Otx7hAKDyjs//zXJbgqHP5WmZFHuZe1
+SZzT9uIEH7Rs/kJiL3BAW/MRJNK5Hbo4NJ5LSVwU1DmtqruwaPlPdtSRATfXOyvY3Q/uQvag2h5
w5rr7SKpaRlpfpsdTHjs3JYidCz7/YXwtxX3pOm1jI4wJi1saEKH4Vv6zOZ1sDiO7HLIWXlV1T2k
nGcokHn6Y1zjHQ7xBJ4PejTM9ulFNowWiEstIYORcUBv4QBfjMq6kAFl6YLwKF2q+wE5j8cUI7op
1QHi1OGwWbo8ZfJaaXpDTFnQJpHxHFjBFXttO6V1RXGDlM+8OYLpgX33pFg/qCtuUcOLWxv/bltB
rh34pLNpCrMbLoOsGV66xlIHtfW2ZUN7wZPmlUXOoCgcJDUWA+8V+TT3J1vLfR5pqqCenA/e8pI8
blEoE99goB37VX6vdFBD0n/kFLSEKyQuPiOaLqRIdK505fdhXIKZz63izbPUft8z8d6IJIiROMR8
P0u4l/UnWJOu2vZM8ccnn9gMy4hLD2THnQ2H0JzW737/Yjzeu6ulPSjPHGqwQyK+0FB3okRVDoX4
r+wUEerApX6W6ohCOEi/8ZAmLOupAkYeVmxpxR4ZqmmpwgKY2GNoshUZ9zojtqXRvW4m+G/430eR
h0Ho+HYSjxHzWJaQK01hkQUZHrEYB4HlQx2EaueQqdsyCI2dEFm3UjV7zr7YN/G2WPliPCXJxlIq
2gvDTLeyIfA7PKwuUqfvo/KX5CuPMrh1wEVSUlSk/BHgJfaAGgMeHKX+GziE2G++o2vSAQ3U96on
S6eTjnIU5UbpbIIc5Y3JMV9OsjhhoE27U5B3P0tCNxd8TBpHzSnpKAL5EL6z8ioEVz5dKXNjRa2S
uTPhoITJBf02GZ5CO5Uu0ZtmHoCscYccd0vdEUj9vDQCLgtSLbs0HZ9rdC6mr5meUMXmpExumyu3
guxAteK4F3107/v6vBjugcZW9jn5gzAYEIy02rOqQs/v6xGRV+lsJxIO1wcEg1pLryZ4zicGeg7m
qVUN7KaPZvuunSr/0ohxJpyKXUYR6t51dHQUuqKm+xdUXpvcqjHNAQT2hik7IwqApABDDNYUUH4B
sQWchfaZz/G34mRqpJ2nyOnpw745QYIV9Qt6TfFtWdrj1hYiBk56D8VWjvN3t52RdZQhzxo27bOP
lj0VRhDwZhMmQoWrkOLWcpGcxdHw/JeHn6U2izs8/Y7eoa+kToVXLJ3iEWPnSaGiItn5xSx4AASJ
PRGJEnhEMJg+H7XgC6CkPkKqCqwgq1nDrtrAIs+/tQXMLnSCnW1PbSmsiw7F6haM5aaUwTTvpkX/
+GgZ55CFcqQMXRQfY3XCXMVFbXK36BxmYqzrM/UjqXA7q1QbwUWzHzQDliZFeJRAHLyHEX/bYIrY
/00hn05VlIf7gar49OgMAGDMMs88Fn2hJB2bL7/xwSS87EjAY8awqWuwKxuvAHgECtEZ+9HaGhfC
5IV5Wh07sBEXzjkGoO4eBxjRI+sqltBI5oAoLljGwLCQQcnzpjPTC7XDrtFMvX1D8193LOkTRQgK
kNLCHKoKxs3TsMEv2cRzimnk6kgEGFUd9sWQefb8PcCnKAoSVmdBaNgN6vAF/QZ1hHBnwT/ezKUj
D0XX8JZ30tTKjeGuvD8i5jDf3ofCncVnLGeHsGGXjDtK6R/y8A5OQ9+uOqgNUiloaMwb5eMiV94g
sCTFgDT0jtr80u52rQnnz0q/Hwea+3uwW+M7y2D5TtHo3vvijmdpjORNmyu5kBm7HBLlTxhNFeo1
Rryc4WFkmaR5BVjk3eBxTaNFVUGIy7LiGMXWUDSmhp7RNznpESCAxd+mZHL3QTy8HRE1RCYwVAeE
f7C0mI+sM8dMryKCI7l6Q/cZicXGEP+hFoQeLyLVfyTKpMb/gZDdFbs09wL55vM6u2z/qB56ifHY
CZ2Bm1o/hbAWtVhCFfgEJog/utuDlMXKPTRL6wrzQErP1S334WaGN737fKZLnIqvI9fC3Yttp8PN
TZ/Jn/bFDKzNPXjo9xsQQqDlMY5h8hhDN9L01ac29kgNfuZugyMG23bVUWUB6a9vGxrskSCqIGg/
1dxY9bM3BYDoTSAP4+5trxNj34iZU5YMlhmYVGvaZqUSO0MDvpjh6coTqlT6e4mcEGqXcWowxkt+
DCRRuSQApnFJtzeYf5aw7l0yFV++LopFaRxa6ZnkzWGoNjSydXuv5FfNBeioLChjaKesKS2HBvF8
swIzHgNSz6C2dXsL13Z0SAQYvIfq3aCSijLvo2A/rTScPtoIHzPDFTmkVO8IT4orc6+SdKI+488j
TTcdbx2Wo1DR2rb+qv2Vov+h3HcmuKvu4sqLZ2BdHt9WwG7qKqbI/I/y12RIbzQT1dbzNeLIyLim
mdHdIGuTaA2MZmHiph3IhHwBkfxD9oI7cWOrpcmfaTA5w9KvCND/4ROc1ly8OGYiVVf+Fz9B4uoc
tGBONYZl6hZnn4AAL5YuEsShO9ApLoq4SVce+SLerkH8An0D8QPSuZmzfnX8wDWRHb6BVClmrPkh
x5gmB0EqhZyMDUiVr33dr/OGtnNxDPReT2gIf8QVMOag0aZTjRO1dYKFddpS5p0IHmM733B1uBvy
H362+PfgH/6ha78/DbsRkgEqc7bgimiVehXXz9JihTLgwnxQdS0qe0qfx0IFJjiAXWoSZTAzH5kk
DsDyMRVXKrpDx5pef4B48uoEvrpvV+rwcw7DIGYAFUqBPK0FwUBMRANDYiLx040vv4nwe4AoY7gX
zTHqZuS5tcqhX1hbYLOVwGsde4QOktq6g0fzJb03vuTlk2vFl0UnNlGPbMgfK1P2EBbld5uoweuA
Hg6YxutTGjjMP+rm24dxpViMr7Pul7rDlAna/SP1SocqtAb221tj9g5dxOiFkeOl4QOjqdja7vDA
fr96AhuOs7lH1wfn+PXOjvxKS2B+aGTc8ACfrtmAJsGFVGXeTlAOcuoLTtLOLmWVtEymIm9mJKA4
OoQ5f354ZkOwtfnXxLtW+HxBrYiwCFfZ6B3xSJ3qB5/itT+8tnVUc0beE0MNuK2WqC+LdXWGZ13L
6CpMxcfMG4dw1KgIKm+bc3BMtfE3ycRqT5Evxe0ywoRkTFc9NRUjaiXXxrfZnTBEbVY7zLTmtjSY
d5pIss6xcc4KLFyfpNewpkjzpqUBx41DzbcX4ZZbayI5/K3Re/N/I/VVgGVh3OtvIxaHsKPp3V+r
UrOyXVX3BEYYjShZHAmLT1tZftHed8MKT6caghQfiGl4LcBo37EDoprXGrJpUiahGnSLGc6FcKkO
chMdTm3rUnzXfG14BEHkpu17XQ0+ggxqq/dwDFr9cb62hCOAunkQ0nH1BL89yV3fimaAdJTR0O3y
WLl14+3uYSOSzYNxQ1pFJzRc0QdPJg52pqS1fE+3YwW0TzbFWCFmGL4ysGKBjrSTReC0IiGLhlQ6
w1UZPao9iFGVPkYAhcwMbw+jQhx+HBSlfwXbcPBJLywHloHugOVhxLx3hW+Kl88QO2KYm0aw08HV
7wQgesb+di6jvjCmjGW81rKKoQpWFkPJJP03slkNHWTC1a73l+eNJCK8RvYwwK+4si1sUbV8OKm8
KYpJ4LkhejQgtz77KcJrz7ilSMl+/ddQ0Vw/qckAL/5uDyQ90EXcnBxpop9YwcMCWCYwXtf9BCpo
qagg6X2fg3zh2ls+la964H8Ze2hulFKo1Ge1N0mxnSlN+xgOG8UxSheTSb9XI3HgbXbuSrBBBkzh
t1CrVMLOnKSVEw33d6TGBtkH06wd6s5/Q50yV0mA8MxAMPREJl7mjDD2ZvqJNMgMLuhIhQlrzBiz
WDa2KVFkbG9Edy6Nf8HB2HggZUsPfIjdeDhvVfXEl8pY7SH5CvnjQ7dr0hKFuQquubsUf7Z4fKuN
lKhBMx7fufqx7vklnD68+MlxZ7JgICuLSWLQGxY9+peF4ycsVmcj5XDMDOHU/OFL6NSt/ZzFPLdx
0v/KyKnDBBmbKIS7KAsz+msW64P2/oVJMx+KquKRTAskEooqRJp2FO37v5fnlIXtlxzEyvwdLjPv
9up3SPaMfyUNQ7pmMZtONsPRTZpPgW9UDOdEJXXU9OBuRPkOCbnf/lm190VqhPl91b2MikUMoJB2
zBXxASt5kw4dV1CVMXy6R3xCY/Xes/D4Nas8IfYej8dxkBDxjQazCK2iloSkhHlu5dQnfsFPe6ua
L8cycU1swodOEhc8uBuuZGPvKKE/Slfz2I3NXhXVQ1BXw9gsDjlDbk/g5C9qQxohL9hirz2oX5X8
5J53g4UZA3WK6bi6woLYxNhazmbRs5mP3j6GHE2rGLq5M7M5WWe6xoiHKALejuG+53cKDGGD927n
fJOz+MdBrgf09eaLtBoyvCJR+1hCifhinRu2cUGqhZ5OVdJ2Kj1oCpclkdmhSkxY2g1fMHgJuH9R
BXp1urVbhqNiMkNrFdtcY1V7vlm3abDhBjgACrtRfFMDnJF6bU5gpIXNBkMSTqA/oa76R5p9Os2n
rj9Edy63Mk/Cu12DSbNyRLZx6TDPBpV48sMEKWuDMq7Yc81qlvXmAqy2LagDPKnh7K8UFXt4lh29
k2AZVjcYd4DWDpv/VkLEEhdlt+Q9pMdJjoQF4pC5gNhnUb85zmpdQMDqWEOyAGpS/qNZSVmuBhFU
Ra36Hwb/YxmW37V5J5bwfI0TxaLfbVCxL3fnKk2HU3+yc24I4Mfi5voZvHbOZzc8k0wtYZBkcdVl
1Hr1lf/bNn5auhsm8Zuda8u7QM5fNCK/kliJAewtDArplKl2qaJHYCRmLmW9lQwomi7w7Dv9O3H3
Yn5v+Eq1tw4EaBR/r15BGVxGJFTsuwT+tNN5pu7/R9kTTsiBxm40aXAZupxbQ9GI18+cq3Dmh8pv
CDAQawRGbiSLuS4qzBcMrAjHnXUxu7M9fh7b3ACl0GO59pYedBUDm3M1+WVMQ0X4BAv8H6fGU9Kp
yFcLKhpEaitK9AtoqBnqtEKuJ6QmfiUaI7vAF+KULUMfSSx80qzoZoBaAaf0NEqMPDHAxME7qbXz
OUQv8FSXRW2ZmCYtfsARKdhlY3apYua/4E4oXBHdoVDyYcfXgwNVv24mV2F/uzpB+ZCynHGS3U95
f5l7a1JTURGTbC8j2DuAmPuplxP+EOJYTtBNc9Z8IzW2eIkvG0daiW38OBg1LX3lJ2tZTUQI5mox
PLD+HJbqAWC+iWmEjscoxQL/bKglJS57M3/wBFC9TVyIzUocvyJE1rp8cOSruyqJ/WzvbpBiyEh4
AM4CqJacbVVy1jdtrUEdyFtuViRcfTDRlLgMIvBDlzZi7ZJD7YWhwcHXgY7+5h6/bMOiJwo4xoFb
SrEONa9nOQ39TNwKXfawfQJUUoj0RrlsOP4X/s45Id/QUleAy0ryz0aHSNrygHTu3XLvSD4khFP9
cHmYIaQLz15PILjCQ5bVZtbTNkAVMGKIWK2lpTW8I9EKRIXXZ8QklUA1Hv9kO5FSPUE+991ZZUt4
U3k/s3bwSBrKoRnTcl4AIOKmb4TNWJ7lVs3g5mpUvGrDJi5ZaoprvCRYbBHgtYvRg0FLDRdNGP+X
ZoI434wXrxoynEuw6qmHHfKEDGOATzotRSyVpNNXJwvysL1iJKxv8se6imx2WYnFMrPv6im4ZiiN
XM++5xmNGnLRNcH7oliKEKQ4WMMKmUzBRyRGKUC7waJnIEYfAk58LnwLp64rfeiTnCzmJHY4pjse
aJjAsF3O/B7fff4T+O5LZmJ/bq01eqWc9X2Oh36sDENQsUHqCgxCGkF8KgESUo7jxVFWlN8Bzhij
5OGp09/itJMdkHyQTQILezHYsTZqV1RY6n51GDzX7oAaSeMnFLU19GYKMMotYkUnkKeenlqxTYiD
c8tjjx4YZ5yaJKiVoI2aDlMVD27lOmA6jwmgobFCcptr89crw8XJh7nfXhPb45eyLV9d3KSxp8N7
BoOThKH01XCMamxtjxU3cZVMynJrzZOnMoNJk0ywH//yBwna5OUcwoy4iOT5ShddCqd+feOwn63e
hdQz9VV28KypoPyd8SCdVvrUP/mqpl4dTQ9JUMww0f0lC+21xYx/kNqkX2avJAlL7rag/d5YDHmZ
ygctyS51Vy2U2OV5d/i87Ya4mszyMd4q4+Dpj6q4z1cOAqSLItMIVGeOh39qdABVLaaV+mDKklM3
iFKuIvZdNhbusT6KkJ23ri71zgW57iLh1hQCiLNDV6G7fowOox/f10h0Sf5NyHFBKmYE6fZdCp6c
ZKsG/OQPueCMjrfbNPOdATQOnjcnik39jbLGOmRNgsD8T6UIhotbiKEtHWz6hWyNp6Bzem0S8Uf8
UxodhPh/vUayiNcYVrzdPZDiwWWVoUSM4BUJl1PxUeI+DLvxvk9Jw6M5iXVyDyChfRDknQV3GEOG
E6/eSsEcurLxhJxj3u87fIXU1qmsSh5ryqMKHSvomP8Z0kJKqVwdMjf98/nwlX63sphaRUg/Mgx6
iRp0RnJ6wko0GCxchi00qyNEgYj++hmHZof7n/OpuIyMQsTmqI/C9FPp/xpypZI+upRz6UDMow9I
kkxsI3oV7QqqOR+ijwxTnBrr1MLk9+iiLxYOlY2daXwfKo5T4QQIVu/WIbiRixSYFFWHt/Ii6C/j
Y1/+4OKI6KtxcccBX7jrg8Rfmb2oKDLZOXSVlts+LzQd2SZTnki46X5NkyxgVQZ/hw9S/pdC8PQC
D+huIPaFJ8FGDQYOEp/SnxruvxW+64diYdnhf3hKdVBXVnkCFh0B2FyEkaGuzTPG/gorPd72B7Ol
SV9noPYUrgkyxdrxosLkPBRommfPg/FnhUkKD6F0lHcUt+ZXO9R4NlNhn2W+4KEc/vosA/RFOphZ
sn2EOpHeGrM/+AgpWir0cGT6P68nT6iwwS9+Cz+yuB1LXXEPcDXXWd+dU37aX7W+g735y6FCpBa0
fAE21OBmn8M7+NQkoCUxRmzVpnqC/0MeOhZp1PTcfaok61YJVGCf3daRM4QJWW53xGA5QlxmK0HE
BIwbidCGvbYW2AIfxuxX7YbiQdbdu4/6OuCaF6bSjkxtIV0ei8HjBXARAHhsUnn/d1pBPt4j48AE
FxgmdsJvcfOd/5QU4R9gfiOdrl8E58idK2sMWgf4ApM9AhRLArBYE45FXMzYu+bzQqnJvFDapH0O
8OvVlQDPghdJt5NUNX2zyIE6j31vBFIbJHWKqs3nOiw+K5NkvfpDXnT6HyJnyDWBaPcHMZzW8V6O
cxl6bgbpu4b+8vK2bbat0Iab3GeBa4OpDahApj0ErU5BGNJUfTUSj+pB9lIT7KxK9HUqlIFoVBDk
7BDObPTKp1FBJyrs5GGxzR0CdXeIy+1QbeKgUUK2IvCbTreskeb4Qwqp6rTsiQ3k8cpWTdHiq/gn
lobDG2P+aPOUkIXiCvvwWQVRwyEVm1btaXZmex+ycvXVvzl7LrNEL65YtEaK5/dC7D7kICXLDbqG
rZgueuojHwXAN0SCKT2n1/5aj1txWfC4QKdQLjJkNiug2slHT80WFYYBCKNUK+OuwFhmDnSfm5LK
rdjPo5mz5GNN1hvCMS7U2Ya128e/2gGJuKAHYqR1Qc53L2DwUQFsHV7nIH0ZpMuc9a9IBawGOt0V
6u2gjzaqmkh8NOhiFHpUZ2OFx5/kz20INwtmleMr6aKIebhKFAr5iV+d/6sVGDHYU/pC7FGmZBm6
R6VuIU4Or7QJ6b7+UBB0x/klB9xunoFfbA9o572aBBPTehiJJgMOwLnBDXxMDy4t9UxMiZ5ktKg9
lM6G5ZkuP6K6d+S4KwpIQsKTTDj7eW8+QSegRKdAmrM6QxNWzkhCtL1/tQknS7p13QTlKAm7WTVp
/emPdPgQHJFhajBqerVKfEEQfgJFlSUoNYeG2ujczTtt5Af52/icqdr9zNeSA9R1Wi5jWhkQI7DB
MO2sAYKWPOLHb9y5/xNGpywWchSWOIUet7alauKVjoxToZ7YojiuYi7N5jc+M36nj1InD2NEuobG
AzRBH0o0tygL1dgsxVI0diEN8xm0NiwNPA2z6iAypTzg2RtvqmnWW9AHT0xtW7u3SJpOBjxOURnu
kXL9Mlc8DMiLprw9BCh/N9XZlq4JAx9CRvxRfI6QqvaITIiZqZLXcinUNyAXULBCQLfnDe0CP8F+
vSSKrg+jDO9C+GPqyc2DunAa8M8ZYukIAqZW6e4jiy9tYOWxAyVQy66kYhnWeMeJ6djmyQsxDJ2O
HS2bppyBz090aZP51Tx9VqoukLlnl3EIOYdh0kwyOhnnuC1goM/l3PSKKA0Db0ylqCLGNPuK97Oy
Fc3yzz6/wWTALETo5AUjEcDrGWzKngR/VuMuiR/win77lGm8XwdDgJW3dAlhxLN6O2n8i049GdIz
mz4e/wQwhW9Nouxz1qcV8Vj/1/xixN6KxZtdAAqf5/umMiicBXyp7R5Wcnw0RePimMVg0tw61mmX
8BwopBUkW8Mi8uRZvzDnungC9v1/8osE70OqEki3urk6GLDenQQtKtcDWWXLIk6rPv8EDBaSt8ZB
OVOYvRYFDx48gVMRz5lOzMY2IzMNUCWl9vm3Nl4ORzYGiNA5YilznY0imRV5GuM3XiV4/oAkfgNX
us19eY92igv7kbtFDIaR9mbIyfLPlPyagop0rx4qPJyuFfSbO40eUMrpsalOcIUekE21+MaeSBig
OU+RuErHEZ/A8jPRi7T/Zb/isNa4gnNX6EPdvlYgTPfN4RLB1JSqIZYve4A+XwioaQbvKHekzroY
WXp0iJyN018H5LNh6tRt4e1O90hJ2BG2IzYvkcyizwqMUwCC5GMn31a8gaksMPC77cO1+kVfzCkH
OkqvPjKrV53uFWTfHuk4QgI446Zn/oG3xr9yLBMEfjpncpRuc+yxOFSPAGvrk1Wr3H9q1LYZnGou
u8VZYnHWQEZ4G4LoR6e7fu77YogSSvdrqYJAPsyKC+Og0OvHx/VnNNYlAlKz4vek/3mR1ecewE2Y
RBBAELrbatryC/e4WPOiztlFdlL4Mr1W5+pA67aLgM9SlnLiFs1K6h+6en/jI1MwoqSfhM71He5V
oaeIO67AvkIR23sZ4BD1QDSiCiBFklcir9jnfylFyMzxT4foGIlPziC7T5yJ1xF07FsNrN/F3Fsh
6k8negGCIp8Fxhd4p5BuTAHLD6S5tmD51TXWGqaZrCBa/LTLJvYMJfZ7okSoleN82DZcdQf6di4q
GiOZbncRUAtun3RhcbyJBvFeqDAFVaVIIEGX2PVyKtpbWMxbUc/bImLAlfKzl6SbeLZi0ud4y06C
38F4T6gnW//7pgh1SPmayjeq+X3ou5ut0tEAJ8CPL4h/YRXsSltU6x2QOTdLjHzt1mTXiEc6n53Z
0xG0EALWwbhe7qckS4JcVusPot3W6WIgUQ9i5ez330RWRGJxSSk6pT3Na+09YMr1vTEwJCKaHtQk
GPtTLIFiLbEJsVZJrJ8AsfCfzx3z7XIpwNQ4Y73bgS2tqlz035Hfrei2mcAW8KRkL3Qx3JXG0jQh
1+wR0XxyR8gVlv3fL+YLDzjl2cREUmS199+gTgMl6zDw3kdd5ntYMT5BLby/8g48b4SyHanv+0/4
JZy6VPwrfn6yrhXAJLYImyDuGqJV6YSZwqhxOhRtfJtU85VTfHgtZfq6N9pnOn53WSVQRWsz99AW
XEDLq0ds3xKCeAT6Roqh6XJv3QYWo7u0RRdSqcro2ntjqCdREruZoPQY4u9oeAL95IsGAIpJejDe
MdQnmRM4KXNx7KxShgJ7OZtXr1PNqNyCf3tMKvb0eCv9+7mdoscNFKs1q+r1hIN0NzgZI3QkRjRb
MomoG2c68lNM+PTQwSFvIjFDEQtd+n57wtpKCFGCpeSrs96+YDjE9fHZoBfIWogs6JxmoITkACHm
8/5BHMsApJ2mBMyMmfq49zrsLBkqPuh1584wBLvj1I2Nnc/0GAm6ZhDCdXY4ESh1kuMhRlPbeT9G
krztGffPatjXkYsBGZA/4ZhFDqPcFosGfocIgEE24q7R+wblNvImyMu4hRTau7Cx3eDs5O3kCUks
jRQDFCeVfX3ZLoHa6nG5Mdh8ghsk4+iJZsPDnmMdcH9ESTTCSyw6EhpeICoCeFw0pFWqAVgZUvR8
881wg9IQPUqh+05YefMcnqEAFhfeYmpWUjkbwrM2x4XCnW4i77GNoEU85s4zI1dlSS72Ew/maTNP
UE+IhLkvQMQhTwCWLFVmt75c3y2Li4qiQyV+5Ju5pbYR5VaM0T6mm+K3vhDg/wqSJVBeKJogMXNv
wuMzI9MFU4sdtm3AeGgKW7U8eKCIDc2tFJtj91tUr1udbauBqIh/exVi2DF+fUy/dftWiX2MGgoC
vIA16sqF9hCkFJrLU/xhU2eCNnj6qEq4tjbLp/XnIrJlQvN/Y039A+4oYIKIZ7pQyaxkS/gbra5r
X321IgKnqIRvFVQMyiVg+AML30AyPxZmUmtnsTmPWWbYi5bzSTjd2SDwG7FRF9aJl2yVFAdHJzsH
kmGz+m9rfUoLOJG+SK+odoQ/CzJt9d3vaYctXZsatkzOHwrHEjGx/kGQGHjH7TX5bgPHTxU3iyI7
wpgtDVnuJM49SNWoITIlOV0JENqAe7MXVhj6MG1DlQg0Dlbcaxjh8JRIWMJcpfzjYYqihxZxsFg8
LxuVIZelrgKjIEKUGmeSmbtYJA5A1JTrn5Kg0zPqcKH4wdnlrvZsCLT5XXVaqeFZWbHsSAIyjkt2
qBHx84X+DDsLU9kbVTpA76ZAzbC0d1BVtAdsPCm/uwzCMiKrzE/D3qCvovU3NZIl/Mj6tD42ogpc
eSiGhKb+LihIi2qDyh02On26uUD4BMy08aNqRqR+bUdooyTAOthx+k4qbYu8EFAdPTC3oEP+l9gP
1qoQPR2g/tULiwRKslRNHQAmHpYS/YR4MP/G/skkWn7LQd5xgk/rb//G3bcuvdN4IDm68H7t8ntX
2D/TMz1ZasaW8AFFXytv0J7vLyQRJ9s+0/V8ax2WitaFmBgg5PbEKe3I+lJisSRURNhQlCgYnQg7
av0719qcfezeubQ3fJ3uOZQqbwFnfC8OJz7opmAaNc+RLV1ZJ7ANeD6bHtlxAAJn3FmRDG8lYREn
yFAckuWwKS6r4+HbVFYbtmpQfcC03Mm+Ox6sH8tke+F9mmSCe/6fsj79rUfcpuSqrm/UpmUFF8+Z
uUXlxFsy/80qO6tfGIkr5ubuxHLDgBG8pbujLrGTOSzm6bC27sE88Gi5C3mwiD/tEYMOt6yQw7Hy
Ywu/DsIDXMZnI65MWX6tDiGD+JFPWio66YvVmh71r4J714pivKS/6YOIKihF2aedPGfaQr2u9QgN
9y6zta9CUR2mJH4szNQt57EYucEQz3O/KzsXWFqz6/s0RVARqxRSXjMtitfr8SbVfzr/F1UL1LJz
q3RlpVNeeLb87w8vaQmBeJ5rwi/+htZosG4MbFoGreLKxkZ8Qt4682ZVajif6WlDZmEzGbd8Nka1
AFy2WULkW4fzbSSrcrzFZ+eMNOUgZHQQNJiuT/AbST/cV0I2eHYdHhZ7R0PzUivwD7MHlyyBQM6F
TR6QPNPNyojWEtD4UbF71AK0+z8shRbBnXl53gvHXTSXJBgD5TaCUGCHUsBgwztxLgWxUQQ3m8WL
804rp9d78TdyapIlqCQzN/7+mffcVQtxLYwjVrS9NgN9bOkT5HhmASC4qP5U0xTAo5fJm3FyP08y
OFGHueEguFu8nZZDahPL3oBXOZ7eKr+k/9jlYfQd7Y7DwOOIO6uA0YuMK6bBsN/LjsRj2gxxP+dJ
zhjZeBHjDJZcxL3K5l+pyWpn1hn08hdULET6HpyvhMLmkOPQGv+r9bVJZF4TsWu7tDuoefhSwzoE
rm/rnFqwsf0Fes9DMeI6MAy/Gk5tFjeUfzPYcf+WDBjWOFpA3yqtYZjWRUbmvu5K0yHxMLxvTIRq
brNWhbmCfGTaj906sD9ttnjLGyj1iM4zraRlo8StecDfZbe/t+2h6hentyKQGHebHp6PIC7B6pv0
nz9oYBjnoRNt2dwdrj1TS4orPtUlLjl3xs7gTvenBUrbrEBOzdHlbrBtjBeXh8IEbjFY8syKb/Ig
8WWTTdDjSLvzZXGEHTyp8RSsfUrfXgMcC3l64Xvb7DCk8XcDueK7qtEU2OeLEIR4pVJlAu2HvUxE
cwVajWB2ZQSqVHktOjSv9QeUiq5IHk7nHdQbRTw1u8qc0SsfFJBe7cVNrdfEx7SDqbs6FIpqtFvX
RiUiEu+iQoIONw1GpAU9gp5fHmKIr+KaJDNuUEtAb5SrD6oOMim8QsuKefnhTV8xzEVMyTSg0QeY
9X4FztUn3qddVpPtSTsmX9j/VCqI3ZYxa03ykXAtqYd4fMI0DbcVTNfC2bXIMdWJLF3TgMkIeDMc
em+HQryZizfmWLJJ6H9ErQIRMQj29g8t1iJRDDj8DkoEyoQnjdwdyRAAN45mVd9jzcWuqEvq5YJQ
otxthB1uZ9eOHz/KVvuzABrh3Pfi4bAtWQ09E3a03c4XOgQJpyQ/4tX2d/0Z+7pMaNTt4EbPV1Mo
EZE2NvMjki+q5RAXWTqnJdW04GrMVMWy0Sm70C7U+6yF6bEiK0LW7KOezJPEqcqqkEF5W1wP4dk5
dtoiDF5SMnRRcl1XDcmDrV8h8vZ065EMZsUqYUdJAhNfBB2FIXL8BSbAlNqWTEA54ci0Zeue2Xh4
zes7/HjVwV6RE0X57q4cQRi7gCGR7gKMdNP3OCUcLr+5QOCp+L13XcNZlGI8kyWnrqBpzfToSlqq
Yf8rWtld8jNQl5Hg15H3kaX8/b+QZJQswLxNp64IW5t6Rhm/FVGJqFpxtfghjHBQSLE6JAEGawY3
RV9+rGGPnvcggEsaFu2ztQmvF2E+b04MWdsXPZS9cqSTkVTUt5t5KkgWw2MeLLzFTbCT58MYC3ng
bg2NcOzrf/4bBDlhY+e7awPfVsJb0Vfu6QChNgWlVlJrNo/L7fJbLY2ybsq/aOSffZ4EmGVKu4bc
5kVEq1klpn8JsdlsD945TflOih+6oKeHcDdJjrDPOKkWWXbp5vBWtnKWL7cGy91FYJNqCfcpIgCW
7b7WZmq6dvrTaDFT7yc/uFLp2ZghIRDYi7jECbZ8VCaG9kbPLWIQrZdNRZAy9TLYx3A1hczr1kv4
W7i7tY4NMJ1CoOOlJpnsj5QB3tkUetGlt6L3GKyyjpsCgPhOC513cFu8byidhl4mViShKF50a6Nq
EmGfRt4apRbz/PAqbkJEhoEtBeN75h4/c9iAjHNk1rvo0CNoufYEYXG3vvtOHhyCQ1hY7DbxaueQ
Ws7Ts5kB2+srTCrfmeI3rLjKw9ZVFmu26lpLgD/KN3/JrZZANxX6JBZvA+nymJIvbtUmnyuuqMhP
WoL8bWqT6XF1bD+isGxtvaACwVBhZUg2wif2Bfilrj/HLM/y4jUVl6LJhCNGgIPIsy+V+oF97aWL
JFHfHIDuPaFHe04jDqaGswZfWWu/9QiewwvBHagD5KIV21V0Dbn6HWnbU/bGLpb6/q6hR65PsIlg
o6WV6EjiykFydinPQIGOcVXbQGEkNis7XYsSvdwPTq4lMCAyBcXPgYBDBcMBGA6iVhR0++p70UBg
Z02dP77Uj7l2UlWTNSli0ln9ahkzGEBF6smxI/AOE3JYcZZxEPLO2vJaPr0CF2t5OjdqdQu9Jwbe
o/mEvc432bIx997zAmcRqW/aJSc/7NwQgsueWCxNprif+Sr2gl0nJCygXDiAFcS9Bt4In+IAe9xS
mzNVYnqam9m46OgMjZ7XYdz+AaO1T0zMY2jiOVmZlAqXvLqO0u+w9DWSmJ/xibE0Zy2/d40KhLRY
ipZNBFvN0Nm2Als2HAsV9idbEJc0NKPpR6Qm0wmFBZR2T3i42MgExopUyk3BMDf4w85y2oxu7NI2
drL4+7EQOKB6SGU02Fm4Jr8IFk3iAYxB8kqTTWhq0V+fbDC0MeNwUxA/TnisOmAUaTBWogPNXWHi
tDrqdNtKLXfHhSS4nt/YwN+V8FlFejwlsOS2GskwX6hxPnxWyWjmNtfDnv4cH0ccmZZXwGmRUoV1
QvnUHLHfsbbQj7cHYn1AAogQkWI7a8Eu+9ZXjox4Ggh2B1aG0pEO/0euemjYGNauvrI/srfFHuMa
PC/YTEJFsCoL4nzxLAyV2gZv70EeRFHAAqV+HXZR+TcoMyNo4kQF37PsuQKakigvOovqOqFv/p/k
4s8sqRh019B8/K2H39JIDfNE7mx4M2BSTRl++QxjYhG4haqPzuXl/mMQyGhI7wKt9A3CvJs4S/5R
F6g1/yqeeHZTileAKTPLJ/4pwiNIJkT9ZREE39Q83LwTVU0iyhqg58323sePhioM+PvHnP9QQcIe
og9f+fF3gW8K4HtOAxQh2ttgVG5PZO7XwZzZEZbIZk2Ex2wLPvwcNZSocie1xhzB+hLX5dkeoMta
oC6eyr4kAeWzcB2yXuWYOUY9I16WH/rKepvywpIasTJKPZcjUapNEVEwkz+Q8eEMbJ/r7fqrlT7F
r7pGjFdycCXziwN8J2rfO2dqGLv5fTl1hKvltjT7EP/1T7k7mUG6uK6YRHkobAb9YsVtyqSlbT3z
W3tWkjhwS2zf9El4TiY/qUJGa3rd854Xdjwy1rYzWvDSWzNP8rgE+RD+qRrdrFjKerLHx+Zdh7tv
806OKrnCPQA3BPaDdG6eQNqL2z3/1uaeEEBPlWQsikR9Se83fe+EwyH5N7ut0yWhID3sslSOidaL
0W8mSoXBTL+OM3SBsHtWXkV1IE6CROKRAMkT4Hx4dnUggUvvQFJmxrFST8FQFFPs3+CIpc89BVtu
JVltAKA0dCIEdOoKq1XgRvhSry+WDSPAmAV+5MteBFFshK89l4g8kMUK57aWnmp5enQi8uLGzP0J
H55goAHfbr2nHhXXiFpbz2JRX402CCxtxoDNHUmxgDGXfKWj6ymdBq/fKFxfcvTjKZnagvQ83anU
gjZrqfbdmo3vbf/uYE44tbsAsp7kMzCA8ewiG21gm/Adhmn27hshtp5VcHEKiPa0qhpKS98KmS+N
kZuY07lN3qnsZP/98huTS1hx41qW7jmxgXp/t/RMlvyLF0cEFvIm+0PtA3iBg230FZWEQjdecsxW
dvO9FxAJBcFmMx/qEOdNH+oNGoY82phDeALZLrXAH7f7fKSZG13MPwWC2kKc4x0LO/YAWO9RGuRR
GeM19WzP5NLYGqUdWQoH5wO3rBiLsJ6lVxnN20cV4u3o/tq41B4y5I8cJnwrSpfQonmckBoGELAd
IammHTYWdignmhqjRgibm7nAI++WfF6mrWRF7SWxkrtzKwygN70X2YSZhQoAzpMxEoz0ltTanBTo
wk4W5bcTptrHeEoz4+leLN2yWXw78S4/GPEMgeRxHhLztyD9PndCaO3oHFnjm/vcLeXcO/ziwBmt
i3fkk48XV8uR02cIQ90lOlQ5OHULCq0and/Qe++xQ6fhF58nmI5HHFJXx/ex+yZ+YpaVuAE7mXZt
ed8bNoq+wYB0rlrIW/uGLU5pHY0NV7Ky7NfdfqnSiqNsn6Y0Rerm8ABeisZ/+yqCwRs8v53bFCPH
/emC0O+19n1BJN1b0FKM1f6YjtHoDjmHQmv1+pJeMFZzpKETvsMODYGtRzrEHeozFy6jwTm0aexq
jAfx4OM/c+fj3/0UQiLC5Jt3sPYwvTjKE2Aa7n1oCdAHKy2n64GUxKkG9jxfMxZ6Rl1i1BZPgjVp
qyXvPx5s52e1Mk+2wYpAyzhHPjSxsexM53Pq5f7Zry2PmIRNFhkAkN/pLeoPzjZjbJRk/VlHQbOa
Brs+vw0DS/qQMeXjH0Z+0X0VDXqkpyZZW8APwacyA0AqL7WfYzsxDg57wHA7F7JCa/ZAzLOxGEm3
tgEThgVR/+//TkpICH2jBEeS00yTxPj4Kh7Syiz1SyHoFJq/QMLeUssK9ZsM93fdqOTHe5FdlDMW
F4n80AGIxYQJct3Cz/FFnGfhwIwhoHdsIPNEZtRwibCz8IS9UTkS/X+M/+4dxUZ8I9NAXyEYtbxl
tsDcVg8+Ct1rsfnjP945IYDejPaXUxAXvtURQEcGmYsHj4xtpl9QjUf9RAf5IdDPZNDzQICqi4XE
XYvKO2L/mo7vTGe2acDdkEGFyEk9ZklCleFJMymxy9/Z672g41ZQ2vI1osIxfXYFQwmdcASIHyhC
bzy2WIC+sl+oScfZ3gS4d+ELeztYxBEcnhM5geShivKIZlNUD2tFGBVxC+1dCmKS898ckVLJBzPG
TmPFAU2VJ0wovezklsbDrtjsFQwygH9AYqQsMnFaPK0YdUY5J8bmitjo7deVRISzMCxulKXOav3U
y3/cJdtWcaBEdQjNZ+zqF80qYhQ4z+IYRqgQQg7hvqRAJvkMzHvHMgRU/Q+BfHIFSckjpJwfJM6Z
eXeluuB/kpaeqadA8rX0FwczF5+8xtl/tGd7LKXiRBFjycsNJ68BtTNU0qEsmcDkT2nNGlXVsKDw
QSCCNBqoFeO0YthMt3spHkrNJAuFDjQ0fELs+RAGewF5xv4Bzx4YyCE7ouhuA5wR4LwM6BeIF+Lt
xPSFU1ken5iAncXy3KKUJE/rDQAu5JFsgISYlR2Y4ZNBMaW702CyQEBo0SxDTDDIgivup0dgtkgw
Dpe5eCwiZQer9Tg/QxTSGT/3Cz9OAp0zc3fM33v2s9y5YtOsV7cDsXHmMic3Xy8LvuALulm59QlQ
iNUsHyW5h0C0sMt2fbRIUb1GLM4I1qYZzCmhJmh3woAhLUea08QKvP6EaIiWrDCArGTvV2dk733V
7E/hEgo7nLtjixKGmus8+Qq4W9SROem5piivq5wEBH2zWi/1GxTe2DKOz1fVq/WnmAnKV9ILeYgx
k/1PPpSuBi/sh6W3RLXSdXgXD0OKhraGyOJzmeSvlygIT7JTQNpPpDuA8cJIaexg5m8PwYw1jeMH
QY4iXnKElG55DSxk8UXp+zULX5m/G1wCTkLPrTZd+up3PNvBqrJ/7xBU5ozsCZLSaEGykQmFLPWq
NBR5V/KQFRdwPcx6RbMTEHm5/lVzHPd+x+/c2hVsWhqauK6iGWRn8IUU1m0hxmUL5knOL0xSaKDj
59E3eE24nH/0AnvIhiHaq+iC+1E2dAEvBLidMEMld3SsTJfFgizKBRNuUHlDAbAeSUf5dASKPZU4
CvWNRScUlL2fl4XCYBPh5O1y+aVS6JnxTkvamJjKpkPpPAMxJWRFqYKNJulcMsTY1YbjfE+a9y62
4g2rIHnasJHO0hldl8uDgkKPKYeYOPPX2V4g74fgfC+8NIaGJWfvGRkwSra7B0hRS1/8v5OzcFBv
IWNwmTPEzve+lRb6hXL5wbghngZXFjsqkYBs/BSA095i7rX7I8nwrIBuVh509yiYwUpmKal9jjx4
I6qeJ2tUJ8HU4VZZwn33WiY6vUwL5cy3zZHVyGxCSL3cYEUqubx9a+csW+Rte8zTNgdxhIiAVn6t
kpKnkH7FnDS8UxsfHFBstr37uzqDwM+EWYy3+KhaqG4th55nGps9x2K0Mok1U3U7JDYONvbIBkkg
I3dKajXGdp66nw8DWrKVnX1ZsxsnRamffiH1VjTp3MHRbJzLOalr1+rDOzi8o+qRRjCWX5/U9PHP
HMi60TrR4phSvtKpkeZtA3LlbyZt23AioXSblkq7vIUblvCLELyApvf90gTNvhyxsLRTwzmfsrAQ
U5enmXFjV8zC4rmOJ8XEmVd/Oc9323S2IEwTUzdYehfCpM4dmTAcTCc5QIEk1xj0K3luDM6fWFOL
d4KeWJCaCFyYiZi9zF6xxXiX3NnrIY3M4wyoA7iV8knvkvO1qsocE3pcEoHpDK5pTR2+keU7Ngir
qBD5EWl4+4VPaODnCfN2wkIDybDQh3CpdfvEKHp/sxZTEHqHktCj5ppuk7zSJzEZi3t0NHKJqKcy
82E146x2a8tcurLuhlALhm6Ri7DB/Pnc8f2VM6x1W/pfIBOznIWEttHM6PXhBWCLJ2CN3qTPeNnE
31f4l7uGxzeFF30vRzh52POVjQ/vKvU9yIjKvQpmveK+7JeF95bnOZdZbGw9d5N9HbDDNaHuBLCq
z8OEG33EC0/Odci2hlb5gnvf04gxorzO5f49ZkBEG4eYDEZ8dODHwgQ29GOO5texWrmFZF5xTQnZ
FGvQand9LtA1J2jnC4C3JpPm1Y0NqYyaN3pqDUuzQDtIfQbytq2O9gLYEH/JGGHqnSxS1IU8vWFP
a1mXGhVpTk2YvfVhTZGPbE/2OJ/b1TdwX3NjwWZ93Qy+JvCgU1PPQtA0OAwXooflxYQ9m9cdKulY
B49ZEVECQ9Tak31h4hbT5WZn1LCvQxyIUeJu8UBjOsxWDeLoSLrllUWSKrMKs3EaHoBct+aEGqr1
z9ZG579HBBRHWwXkCC8y9+Rd3RUADW02ccIqAkY+uz0UnIKCZDYQ5gayQh3+t0aUZIz+uv2W4DJS
0NYDo8sPFMEY7yb+0Nws5S6TESW4G1LNTcfGJlWfEVuIf7/2of3CdLLmXQiwBv/6RLptThluSIMg
la0TUeEgY4l+dOt1u8f6ZUj9l8zxqT6zRc9FsNy63XhWvUJV/vJgPXrjXs40zKnTBbYZdnBo+iSR
otdL5bYASYwKVQllE5tVrHMmKFxdMkKTvQNIg9myGGQCUoOiJkcSAEQiXo3mKZUKASucEAH+tr1x
Zlm7v6L9aerZCIgKRrJjKV1vUH9HMjfTQJNNtA3pQo1VDmORPgUs3ANmb7yVIa9h4gmfa0xPQUTT
ovLpdKv6kkWDmaj9nO3LMM1hsn7E8R6+0m/iqPQCdE+aRDSvCj2X5l+FMUaZoHKT3BItSzkBX6HP
zcTv4GMxRrwGk5WAfaWEspGhBUaIZhOTB2+7xi76OuYkLufKOpJqYfHTpnTtonRyclSZSnrb5ycS
Lj2WPADfHxKWyd0E0aMSqhK0/HqJ6C7G0ZCJ1G7U+3Z5aSQe/CbV06vlbbFLZbi0gy+4PPH5ZEaN
MbkPfbVVIFImJZe+KImcTOwjPpSUtvOdQllfTOiBEcOMcKqaeNC+y5novXp+BYQzKYKV0/18a+Wy
U7gdkXbQjzvDPc/VHvR1dP48pHXcz9C2xJpSCnUZRA+hN7noFcf7fVh2sZaexdJCMS8c8zfoPKCB
GgZ8aNnpVvqpxrxQnNQkRdXF9G2U8wcu9x6Svg3U4+uI661UJ6aRr+IpozAeAlooPQJmMnKLUkWy
pAwVohSEDV2lSCfZwji73gSSZjh69/u2u5MNLAMgS1ADNRbU/UQ0ISoZ/R12K2GJ05LYcu7k8PsO
PLxALQ9lM3gL06Dt8fr+AIEcb9W4RG6Tj54QvTE6sTOM40qLuiYVvrX1BEcwBp0+A3IL0OCPj8s0
OQMrexti7kiDIQGVp4r+uxpr+Ed0XXeN14QyFvrDZVzaEp6OeqrfYmdE1TIi1X79rY/Jm/Pri1gx
rwCsRa0XKdBeBLzGdbsDttDggijhQv4aVctMQjbQfU+cm3wLH9jZw4xQeqyKvw7VizXrHDgPHjEt
rmqGUtka50CwjNj0ySQ92j3pDJHK3qhM5ymg+/iVifqPVRnU6sdEr0lOOWiOsfyZ35GZ3+MFPwSf
gtStV7C4vZ+jEr+yFfu7QAGgZxog6HD81jop5SzykhwnFyqDsG9FwTCHZhaNrnwM1CXxlFiq2D23
NPfF2PbyNRcCAmssJfr/Bo/FYBOa/q+0oOXJMZTF4xzoN9NMLh5WUKIPb+CR3sZJ2OgHOP9Uempl
k0S992Jy0IknZ7kgT5qdWOVL43D/k3l2e7sYrAbS8J2664qmwAOILZyXGyjOgX2ndF1/YOFyVO9F
UbsoYBRZSiILyHmMXd5rui1IueU+y6fcP2zhoceO2JeJHy0WnbIXS7uGK0psXQhoiUNzvp0ggBlj
zMLp6KI4LN1oOrGTwnDYfRZfZZ7B/BWD3uYuxOZA6+Hk2ULzt4xHJUmcWMmQeUoqb7VTU29Y/yKP
TVczrILt/BDIc/LcpYIaSLFk1yJhKPfZar0O4yoYEC+XecFF7OSHujz1RmXhdpgG/+AlH2dGuRZ3
mgJB3dEaags8sL6XW0PCVzex4u8IuAOPmWIh2OxvpYx2WogEOecVw0hWm8jwDPhCL+QYSAIpxuEn
gGbD2OPXHwhwQud8MIa6tyF1DKTVLI4DSubwAtAMsIQ+mykkQf7sDJLhONZsx8FN9KY1b0fsO5Ef
UgRoiTNqFnzvwMCw9HLUc8eXrQvu/LutZ7rxU5pUi3qaNcmUmFEImWL6vj8nwhBDiVwyaVGYHC0R
PpjHeUU2IJ78bNEz2+TYMzBmfxMFkT1M8bPAZ+3OMp7K94q9CjEYuCbDLenwjt48wy0Bp8Pa1vAX
sMAttsnf1bFdwvR6c573icfsDlf1ZXuBHHHbMC3G2QjCi/+fQUHLkvjfX/Vfgcp2ANjWdAxDJc4K
cbmse5bSKhkceN34yLc7/VizlCcb5mFLD97v6TUmvalZU7Yr6LyiejbbZBKVaZTTEU1XUW6g/Mni
a4FW/xlsV63i4/uC3y8Occ1RHxgZ8mr4diOzmii7uEgB8Lh2OIylyzevLKh+i+90TnwuLipcecSs
Yrmie+mvkcpsYlPQJIz4Z5U0+vImlA4q7aDJ02Yi6+I2pyX+SFO8RR0CIpwhoYXWz1DqquffRK7/
z3VTsxzHMY3sZsckjilwVKz/MN/ehqEZouA4cW4HRoZlXBsJQPEDFf9S4R/kaWlNXNK964bHe/4J
wAqwbIUMotbBxQpumnW1Hr6kvUTU61mp+5VOt3CcElXbpUjTjgZxUacHMi+iNDBkJoVUsfb4/Ds1
XSDd4Pwa1Elg1+rwAEurTF0ZgDPYrH+qijdMqy58nqntyhJoz6+FzqY+Z+b7ftbLFzt9TSN4kJfg
6aArdDlp89Meh4E8i7FHT0ZqvIeDaZ/bsfbWLGLW2wTSTq1dXdUGYHaJCG3mK8rAVf40JFYIt/kx
RDq0K8dRsb4UTWrYexwxQ5FPBeUED+Vmz2h+Sky55SvW1Z/U/aBPwRGy9iUfnb7qCreWorL60ApQ
Jq/xtTOw66xWFS2Kl4KY8frkUvgYvlmf4TceF5Tr5W9gq7r5tgsfaNyJIqa4teHoyXjcZMNYZGRu
V0ogTL28rUeWvcRtraShEvdTt1scIvWRUBu0oUGE+x3kql4rtFl1KEfMeKvdPiSvsGuSSNBcpCD5
drxjZSHmBeU85+ba4NG9Kx8ZBHLP4FJDPnw4NST/uF9QwPDsXBhz4LezzTkI1Dmtyd3TWfJ5T4Z/
hneHJZJ4bBOVe/8FVgmx7HM5OrpggT+gvWjilDg9dGQ47/Bnqay7uTn6rf6lP/QZM/1BAcKM3UK3
yGTrsXJCB3yWRPeg2T6Ilu5KxIJzd5yZF5SedSLdJhNyrbQ4rr9EIzf7qyP2Lx+2E+AmIGjWVd+2
Ui0ydGZn4tSdA/51KwHkK2kzUlT/kPiosKQXHSeQzQinoqqNLWAwmUTl2IJmdc7/SSoja79rxzWc
wfEKu7PO50U1V93uCN+6cvKHJcut7mNH4sEk1GAq58l4U7h1drH3UT/BvsiKi1n9H4yu5FxMt6WP
Bm8oaBZgW7uWcae+34xJ31NuRA56DLzCl2vHfcufkzZpmbK9PnzYeSQq6iRT3n40huOajlg4XxuZ
pn8Xfu91fOyRh/AMpURkt0FM1p6znnYIJ/xARFYbqs6NSKGxZO5wIFtw3Wg1qYiJL66eRQgLBtSb
T4jkKDsfDugm9iQeWTRlhO+URGyDmsq43XkHuQvaX1oCbm3qvZHaSfeth/7dcILa9jJ4o90wfqwe
6SXDRgaqxjNK7oRGm2OA4juh9qSpbA5b3yRW6G2DgrLs62zk/mcCbF0Rli7IDBWNZLOaxVwCxE+C
e6d7LD3jAdDPAA5m48JdjdOOaGAS7yVQz8cVN1WDk2q/PCJw21Mb1lA/eAUJht/9a7mCHPH7Wc8t
SQcWJVnj01L9kPTkdvfhUJ7I7acZjDKSQYK9RriSHL+OMwTHV/koeX4ouxe00/gBY5tRf2v35Iug
J9+4C+cZ3Rx0uWienT1s832zkmespvyK4mYSx/dQ6G5Cy7NAvXV1GOlSj8G2ZPjMmpwADZmNXs4U
BowiUfPn+b3cU7St3JYPKCbgyfUjfoLI174DQTiAB0dPPc3a2Wy4KXNFF6PK0kkATEyi/qmtwY0/
ztn91EY0UdEzGGvy2+1Un+mYyFO6B4OIZ6mMD4tno/Q8ur96yBDcy3wYDP00VOZXoCYELE9lBfYV
wcGc/h2spUeIwdk/mM/ggOcAbC4dhl2cxQ53pjVxYZjqa7l65E8B+gcZbujJxycW1LVLH1CvDue8
w6EqB1RlcN23HCbBpM881xFNIZVoUqoNLKjMx2Oh2TiE34OFUy5C8wmFLegPmQ+YpnRieOeKA//N
UiGP9xhfoNoUSGe7onzRyc1aEw7sSSGHvQO7C9hFhyRRElw0mEcbPRuQ8rlgwineQTFPThpDRp8O
0G+fy3vsvH1B1Y4fu2MR+h1cbqO2XPf0Mf+HMJvhUnKycEKAo7snoDWuVwozALW4lFARoaBIKBNT
ex7khIpMkUIk9VJ6hlN99fSQ3lQ4vHFGDWBC/3CrF8y9qGqY1Rq74dnyUz306Lg3pArf8D+NyX7n
wrCazoZH/zBQ7JIWgQKUgmPWvBDcjHYO2tgtZqlxk7fj6SYCSD7yhQ197vysq/EKpLHq+vv0DrOc
CPuEERZBcnYRc3tUW8LLLZpfNRt87DYsguvIdwq1+XngE4GCbtwYMh9CsyQOcziMp7NLCoFsSRRx
vRIg8mgubE5Nh5bCIsebmbTxrPEakopKW+k9V7oCJjQdNPrvtDT/b2lrKQE1lIK8abyCePktZq9X
HaXmXoLE2tAkPo/CoZHQsVU1EaVFxulQdjHrKMMclizT59wa3xymbchh1+8zUi+yUripachhr4jT
FCGJ6m1YskvE4t6kmj9IOYeu8GBU19gZTnEzE7eZnekpmcvm04VSywy9o7qeaUVa6PqlFt/qgKhG
+1NEwExuNFYQ8esNuPbl+UX7radZ4vncRJpfauRKubWd/MKe+7+FlATxYWrGyoKSYojSzYoK0V4w
afHhOWv/iNJjcnwL4AA1Y33LXTJ65CHlWdBotP18ZAYH1eOyxzY0WYhe4W0pg+9ug5TWiDqQ+x4v
l98h3JJ3Bz4kEQaB6L7wqGbukH6OEqTyuvNtW2dHWcmieLhTnB+yKcBA6+457EhN8wNf4YEa+LtQ
fZ0lodJbEwQp7V+9+cHkxaOWwdkm5LWRFu5WmbjGyhyRU2qOtiJljaiCDu0nFDn2uNLSWiRJc7Fe
lSGjnvyjwy0M49ddAHBzWubPF9WkvLOkgwZvZvmT1SYSABpsQlr/Bqom1K1a16mnlyWpcoIDonLB
EpiJJ2p+3yJmlsYru02MBADwumHB8MeygfSpEVZBR8BYgtm3pr3sLQoLDmdL16GnzL7TiWgsK+OO
cKMC7R/pFU9pb5Q/3Izzt0lgJeiqskjptIrtf9I3ZYGFZMrC5kEND0MGmaYg1HO809h8XLH/XZ87
U9ROgEz3W+VISZ2WcrqAL2Fc0SNrlK5Yw93oHjloNN49EJ+yvMw5AQ4h8mzTaMLGXaemp/zJTCuv
BNGapBRMUlNArzpft95jFjcarPwaPquppWWK/PLYWxYD5UX+F0SIWAjyf953emPMSMQgzAT26KJi
+RNCuLMFacYeU+Zt+cZ18AiPalJQRzu03O/JHNwvEVQyV/U49loWnE2HdevkgoMftk9n4om9+yIR
OuFpJjgT4RIIyzr0//dE6b5ZP9GoPXK8PJljcKx/8bSWkXb6XgWwoU/GJQOiM4oWONgIql7MKqHR
ft5cJYDgkI/urT5RAmHH1xHiwpQj1aFpxoRvYq1BGXg3QLF5lHEGq/5pcJofzL9+QcHliK8sjyiH
fczHyKm1Jn+Ih/dHYcsEtAuK3sc81hVmeyaiIYuUuAbAIMZSGjO7csiAmDwrYZ75saTGc3CSAG18
QQJOOk0Vsy2HGWtaDPBOzqfqR17iNkeFYXf6DtMQx9upTmeF1IVeyJe19iyPHFU6jxj0Moo4hUQB
4IYL54dlsS30UlvmCH4Qwy4A/izWgKub6pRo9ykSN81sqfXSub1HzVxDRHxTVBGFI1lfG0nSuGOc
yyqp2rK211S4nLshg08Lm0ghsyI4hn/bff8DuJbrDok2YhfQoKs6yUhMzSCpREWPd3lkLKBc/q11
NkyPreRCoL2OeCHTdoLkHxgH2DXk0eguMIb5+ETaiiZWnhhSbiJsMT+FVMSFbJuHcNBUXM1C2Wet
zm841lAol4LQdl2L6j+PI7E35/u7ej3iiwIG/6FyJ8IpLGDDOjV9+HrRpleSEOLamOrOY3o4XRiV
IJsAMykhAJldjaikKb0hFCiO3r13k5lacBcn359EuchAl+bvSi70RIxPS4Gk4BMCsBNarhWwWo1m
2nlLjbte9zIOahcPBuOt+2d9DIe7nj8VkCkd5kXEKFtmmZcKjJ/HZ10iWtQutb/5517ujKMgdfta
XdUbZleeB9wu17r4OI/dZYJkEUtNIiDTesF+GBtVT0HxR+ZJwwIdoF2p7umlMdFSfEeTd+wLa6jT
qul5LAjChtCQLF7/+kLKhfQrGGxu8KWYKI8ZQatvnnXlZBIM4WSzE1i/bzLgfSlSW0fmrjDKcoPP
hakp3bHyUiNR/FQreOrpeUIAonyt/27MA2LIU/vEcVxksEO6BJKXgNu20hZ0ac56s8g0jygwwbkQ
m2FT68MhB+rPxWo6FTik03n7XJevsB9nMqRwoNGgS+OJoMJ0u0gwAKCMyYpIg1WZ0ZcCtd5CgDp4
Gxm1cKcfOKgmILeoEzkZSK0x0tESXyLRunQOvJ+LjauX5y+iyKfjSDz1puyqfyPFYUcIc1S/JDvv
Se0dlzH1C1iij1iJT/8LXEPauhS+uRlT3UCLiwDEvDn/4PZul8eeYGzWSTloX5AGbzmUAqpvO2CX
aHyQ9JomIsSQsu1XBXVthmZDeERZyyf1IYxi3g7Y+l6nLxsF8eHvv329IfkwrsK8MFlWZA0EQ2Ot
syfQIfpvGnDWvVLNmVc38NF/cFokcaGPH1PxX7U375QVW4oZbOT5kU1BbPO4EypSr+qBBMhdqrOc
DROLInsJiK3yIgkq8RAQBWISdGMYc5KmU2G3uQmIljxwzEP2bO+vn/tHqAAY30Zj0bhjyYI4n1Qm
BZ7i1BAg02dyG9q2CnaW0+gIUjHcFU1sLL1CF56u4tgkmAnXZ3WdfVbDL1W441h1jkqgkwHP4iFp
c5R4cbJv4XhrDYUrRKddHmtKSI4PaS3srpw2sD4a0K981XhnGyDkfGqa0QoX8tRF//n7lwHw/kV0
GseMttaI2ABsxUtJn4+THEm8tkVLw4agkgzkW3BuNjelDxPkah6eZty4yNU5ye0HclIpLt1XWgq1
1kmHgFhf9hoiztNMAdVDauc3aU0RXQw7xC4p26AaplWK+P/uUaNZhTGzeNRsERXv14L8CWI8fmTo
Uq+P5l2vXLFYmto4qWYle7KZbw0zew5btd3Y1JqoBDiVE8dmty8InvPFutTfA2za8+8OTv7QOF6w
yZ5AMJMnTGTsQA596T9M5pHFZmQARkGyNdV6tMpfePJSyJQRu1hBJi6HF+EK0X5oOytGQ2VraA9g
jeaYiU8w3mQRCpBW0vbAOpewyyXk22qM2Z0iHHPL+v/adg06o4V4ESPsdZipAT3a6jbwZe4kMk8B
PmapwUwt9V/xKl65wNGSehgiIAk9GMeVTT2YOlPvtj06TdMGqoLcklx7dm9qDC4tSyWlskrZQIUn
ZV4fUEKZ+1mzd7P3Bj44Q1Ymi3izIlKZORcfqaA6g13ybOGNhHn5sy2iOZXQgzRssaLlhvnDsIy7
1a0io5oX/6/ZHkUWKcrIqyGOTE9/0RwElSX5eqgoPZTal5jw+qn90ZkCw+H21WoekFtzIvEPd65Z
feW0G4TDM+JyAhTFNXyNfEFJiWCfNeS8cbPGvSqksLuJx8l6oaxmTiLtlwSOBYB3YUygUsFv1e4G
+xqDMYLnSkO39/55bXpB6koeROcNe5mS/bgzKGvDLfOdpOEhP2BOzmCVFbrrwVeFWqi2Qk7xurJ6
FwEjqN4WxY0XzsGVUiNptwla9x63JE6yz0hA4AT9GsBHYebsU3wanjonOUZBN7mAuP8Y7MZyEh61
wy16CDOVREas7QzjLYB7j3dEiDwWVFAwzCB3oz8aYd0QhcvbCT9j0X37I9n8kHphVWuLTwx2X5co
4OcQ0WjSTg1tjY0lQ7fIA6wh7TI2JBYhlnG3AG1YSmasWRHY6Oxmtl8j9j1Z5uHjg+v3m1G+I1jW
DlO7y+lHS2csR4a8FIf3TrA/ZOFB/r1TyiN6CM3oQqH68lqsGQcN09TQAESqQZ044wkfJccaWIBO
Zxz17IjYWd83WeWmFb16tf1+dX9ORJhJEQRtJoKlwHbY6IiZmzw2QVJGO9cki2Iw1itKmPQIZazA
M/etjS91GdER2TQrDgkmsgiwjHgUcsD8PPI7V1OPnU/0Ra++6V58r5mDwlR3oxnrEnmZiZjqWM5X
bvG7v7DDU/3l3/bXPoNQLlsYwzfERicsyXuuFiAz2273CuE609TQEjpt+HgAjLcgV0hzdLVBwkXD
g/gmFLrDvV5y1Tep2m7FM6WCZLLRJdgMnH553AfEKr4RXMSKn5kH8l+DwLitnWX6SBYecFpR5Vo6
cBPN4EABKXEWEeFmIvy4MLvfTcGMmpZGue6x4JlzYD3TWdOmON+s28mhBNgx8dAy73t+wXEKJFgv
9SXdAbUY6TWlUy5xKiWvdY897bxHsdbjZEXJxPwHttQcclhTvCGsVaLaN9qun8PROjBrNxECuIuv
f/4ionfI9bms7I1NCHrcDYH7VAhZKVG0JMHKsrPbNbwDKzXkjQ+z3RxlYvvQ+g6uEEse9uNhy9Lr
hS0CAe0BBwFDoM+ywGLhBfMS1UebDhTBKeB98THWTEJ8i6RHLvNyzokqMaxtd0J23FLbB0dWb7Hk
9/GMkXMZ+eft+IogPiFCuHqrHg3BVUPntpoB/v3iYwytkDSJ9GW51TVyww5dIKb6H/ABxD2FTbwB
p0Fh3AwhG3PZhfvNOa1htKCk/tCnIikQ+ixkFgqWqFRKdVWEhkN5TmWZofgowIMbAmp1xJN5pCg1
AXQj5UKOlx6BoYe6LKoeivRFKbkRP0rJlAAe4Axmqj5UipGWVTmPzEeX7FN8AvR3CYbmKZZlvF/p
m1/yfIxqHlwSOl5ILXnz94wcvLx5ILdibUb0buETh7JeXvtWCgkAWQpsDwn8ISIxE4NR+QHRacMe
sWxaP1zkEOaB6PTwhb8/Ge6Xf7047KPQa858KHcLGIui/5dNDpyJ3QehVCXY/s1YZguvlPNoZUSS
AmzCzpL04LIu1hQQXM5uogoERL9/n3A4CwX4cmYs/DWelUWDhb+9mMq/jb4c4WUVEEkKNrTTqRUN
pJIyXbMGeiHLJQfH3tTnca6RKj9A11I2OSbmQcL/fbEZW0nGQVRMI3E4mBVAQN4w6Rt/AziQdIrb
cqyn60Zcm+s91+6kLC7u+5q0/KYS4FjeW7QgbQxPmUiivmGAjB5QvF0TujOvN6uqHMSoYK48wxW7
MiBX2RYNLqGW/xKYpXorDsIOBtvPCLzcUfnppZGerKB4OJJIb+YMkRaFU7xTrtyS6ngplOYw9Tat
N2IZKL+DToWa3pZ7xxMg773J3J6sDm4Yb8LNUQJUoZ8u+lyeFe4g5QmJdPRudyrqAHLFxk0kzhlW
87lSbOwXmI8V7k86I9Oz+q2FcuC8YuX6C/MYAgITH+7bpnCpsJK5FKqC+x7ZsM/4W5yIO3m6cGyi
+Fiop8FCDkhyi5TCIypL2o6LmES+pVadn1vA9KGVyqMv0q9deR7WOvKyMYm8gIgkgv8TU3EEANBM
fGqDYu/AKZr5KPktj6pW0lgA7v2/0g+BbL7CbfCuatBn1NZqy540vmAH8A0PmZRI0w0ztx68Bda+
qI83QUfP659xddhBnxaeZjJk7aZVK3rtRlU/aW/wRnwb8ix7SUughArhOzRlYKqAvbWkf+iwbRgR
XMDLtyCJWBsifh+wjNWMwjg5YxX6uTqFBh+WEqXxxTOR2jIWg68KFhPEnf3bzbYdLOY5vA91Bb18
Mf+US9BPMGC8m7Nq5zF2rWDdwTfuXfQtHX5uWESdRbslsnXTs+1pFPP6Bi1kOvRh55zCkU9hDSAG
Ue3OdRNowfj3qXVvget773v4cvh5XYZX8b6STPxphO6ruNNqo5yZ+HC8dn8jdh3TZ07Hu15ooAXf
12TzjJQ8tUkT2kKMjNBUgHo732N3zbafAC+tPY9y9lOYV7NzqMLAfOuJhON7+MOADSS7rNXALHtO
MVRWRDjQ+PGzm6xZ2ToIiYX2vYRWPh7R9+zNyXsgI0u1wkhSjlTfyMJNfsKTmPMoR6pb1UGi185I
gNYkLKcf6dXoo0vJFATorT+yP/ZckwLuEFS07lDk54ylsDwFfv+rOhPTpyB4ga8gk7p2rJ+lx+lc
yAL3zu/yWVuLcrYOi6Ud+fj9x/Hc/njv7i8Bd0ougbM7M5SN6w5dxrArG+CjmarOLfQhHB8bevR2
HMfSUVr/dANZlm05+iWsCmjdd3tvcwjbcTP2vL8VmILx89wYBKAswCLjjjd0bwpohcGYUDdZZSQG
fiuGZ9iVK4rSBza3n401E+XqH+Go74rcKyjnH0xWY2IyYSiyY1oHJCygULzkO/Y0SoMxXcRQzqQx
AOoa62L0m205UojH30s9gWI0GhJNuYD41pLQvHAMB2XELlzZTwxD6DX1u0iM7cXe5Tf0GSOjP/1B
J2LnC3eEEEeNtVqgKSrVMwjnsPvjIPCBfr3QZL1UfN5a5RtN9FX5QTmVwxSRzGV8gltjbSyysUFu
ZqY41kFcPhLK++JquXdTZuXFSpFJxRQjFYTPJ1aww3FvHGsPIgDaSAFTn50fbtaE4+1EYZdMMw6F
vYlQABIdGQUloT2rWm4QaRNLbfENsaGjZLxddoQHtiGHvsPB3GGIvDi6RYLye7Ib/NQ/ycYHYll4
UWLMJP6m9uQb55H+MDE6C2dCpziW84xYlde6YEy2riiJlvbRn4gZZyVUvyaRhk0PzDzgakvf2kBF
XQOMJU/Nh1TUCHg0qCL2PaGJaX+MS9xLWbXd12hwbcfAjJMt/yEf0poK33LW/T9gAvREc0rWTP0w
nHHmYQJE8HC3p41fNZaWb7fQ1WVg4I1GQ7y8oaI/F1lkPi3xtamGnwukZDPYhiX9+darL+lRZcgK
pTfQXifhO9C5BxxxBA/Vmg/cItB/w2gzCQXTYi/b84MUix68V03igkYVptK2ukMrOiT0jqWJb60r
9Bl/KKnIgyxZW05zoj/y5xbN/0tgw+c1YaJ2DED1DWiFi04xYtCQOXe4y5zXKNHz71C+6RFGi/u4
0L3JAILcHaqc3t3jKurRanUmwYfdEvhvgBvF4oxQ7oGnloswfBnWSap04/1DnXepmWKkknqSyx3G
mnujJ6zUXfRY1oygICHdcJMqUQ7O5gVxnMYfZs0TjKUYaCEm0ESIv9YlCJCZKnzJof3TVXppLO0C
sKwd47WeAcuhYt6bGkygSEPTeAHgmqQZkA4II1zbidXus7zwEU93CfAQUBsDLSHpWmLze6g5AQLm
9iFSdpHQG18fF277oTGQD653Qt9KsmvamsVhlZHcqeN32EpNOVNKk0OEtmATG6pDLafFhcMrnGWO
7rzP98kShGDbUj9Q/HN5RiMGy8qFX5wT1YSBt8PX/oP3TBJP7bHGn9ewJWNds0hxslAsAPEMZ9hq
VdLphVUNxtUYecdDkuicTvDu0RvoFJTTvBNL/CK3ZUt3+AlQq4SvFdSg1JMxFPg2XvItaWySwrGA
sWvWBSzxTG8tCf8SD80AbJPnef7G4V3KZqJM6CeXkwcq3HXkcYZL45vgjaHp9tLJWI+lHwcniC4D
wfclIkiN+UuDocfc0g+4RNEO1ek4lgS7fC1HsTf0AnFHD6brBs6zAunNIOCEd0bQ7Yr/BZY1wAxn
A3kw8TcsoFLfRXkhiRfPrmO8Uen/ceepdNWHpaktW+Mh3RUKJ2J1Cxn1w2V7T5RT1IZRsf2YjC3U
/xBoZAlxbroK/fR6rHaggrAUvsYvD+I7Oj1heTOtVTAmGaQ+6zHmtuQbE/OmT9d0MSfKZFkFSees
TKVss78X/0mGOXnHRqp/S7P6GnWyU5K+NZvsWRxd2FdvEklH79MA8zSkgcAx1wCEyyMr9ZghC062
cZzS7Dygu0CnLtnK4KYeannl7DK4B2MQLcWIZ0WQfcS0JxarVsqrUvCHkkh8OH9W+SwU2++rghl+
BaivJfVVKF62b+GXt8lwatAlVMjtLqzFhWYOHCDCYjMh9xi/4+7uvcKAuZq34v7zKPBtnrdZgLin
hjErcWyD6FNl61Y73CZoNu6VjdwUdtjeHgtRvWbxXLO6+tFN4oLP9x49YZe9bH2H9k/b5llBTyNz
tN2EFBjxKhcp4y1nTY4mS/jm4pc1XYyyIVfwgYXnMgn/5/aonmfZYkcwP7MrAuGc6leGCnRYPr+B
Inw2kx1G5g5Kzma6OceQcM66G/zOUAbcOMetT+HSyZkbvsJ31lwYjU+8erbB9R6HOf/dtEtHsdyz
lSMZ79Vua2fqmVjcWNxKKxcH5CoGIuFQJYJvqq+7ucrXjnizgxBCwY899sIiNCZRMRo9fTxRi9Mu
dTqz2YSwQD4Yujz+l5i/cg+TD6XoBm+C03y9xjrEXMaerYlbdyXSEY2bikU1lGkKyreyiI5m7Ycp
yFl24bbsAPe109zULETNcTdpvoSEW0AXsI9HxuOkAAjzOBkssstiBH6Fa1gR/oNCP/209brp34kC
/O2AOtAN9dp5V/IGPJfUqSpsATcO4CmfDk+sTaijEeH91y6Hhb/c/D+AVkr0Q+ZCArdwzZKQsPNp
A2zUqLXRIEEcWHDXLVmCL/PoVoRmv+sDcL3YJD2+XCy267t93VE3N9ig9b4vULONMYQqOMpwKuQX
lU/Oj95djkSQqL/nO2j207teVy5ccRmLgx5IP+FmbqUJs7Tgl6cXo3BhUVS2SY3uFtoXL92U1WDF
0FeL+AR5Ngz9yhF62P8rYLwqFEK5ztL/opMY69gu+LQRUS9D0S/zqzZc/YVX0GVBHV13kJm/y148
2josrDIP1bcOyliwR5H25c/UhF7fZwJAR3Rjywy3izDEaO6vAsPU6ea/jjAGRC6C9kpSQsqXGnJd
X8rDq3kK9dTiMnVJa7ItLmNSDAHWdTZu+cmJEIcFG7iz8Evh785ttY7jTN//zqg5VOS6zHovlgjk
OnUQ2PdVcSBtF1JC5mmKeS5CHuSlxqooFmiaCRmV4QDHEiroC8f5ajFN93uXAFTTlmZL3GJOvKjN
5iCBIglLcWC5vdGjnVlq79kDGz85RbYVouoWjKAFLPOxcyK1qjcVEkjCE9c9cdyrqL09HEsAMDa1
Ur9NsAQCL0vuxcjs0kfIXQJ4E0CDU7bwU+ydGTNdFleZUHbULyLXJ11jtQBHxjVvSPBx61Lq5UIT
pb1oEd8/Ndykwt+fUwluyrC/82kPo1d22xreiifty5aZrkuaJT7tdnApP8jI/1Uw1AWthS9ikTsa
BPUw9nhrhI1chGDX2V7dXysvNFVDTpgr9kuOl0vWUrDVmR7CrZFAgmaeM2vc9DnxVU76+M1X9F2e
KJOEBFxwn6VP71/e0cbcR7mO/zatJS9uuIgrMFLUWkGAJ5vpu8KM8yHo9vsxps5HmBLI1/oxT6m7
oU6LwS77Mmkg/ZkHsngqYlJmNXxyIkZwt1xEtgX452Jl9nt2z1aPIvDTVZwT/XctAHpD88NNmtGB
NuWxkWo40lz09n587tdkDuMUmQ8QJMBa0aMehSgtkbA4AUUim9Ijx8EM46SZp3WEeFvFz6YMyRyn
0QdcJlcDnwDTElrt8+YoviwpfDGyF5yeYkkY04EkN7gYJj9Qo1UPWZt6WFRo60tgRLDwqr/135cj
W3UEwQfIB62xbXBj+prjsJM+qwlf85Cap7a7icdT35mfl3DgPXByPcHasBsOjLLfS2Q/O3Y9uAX0
62FFKvclQnX+uFiXB79hp2hascWNhtEvUKgLV0lLlJQ/ZM8ipYf1a7KCdg3e9PCprgozpmXYWnho
F34OOGCSI80jQOjlUT2ALZMZUUCsZYpQVnSVr/ZbPdv9fif9s+CPrib1pxDl4jYVKWmSLtX5Yaxj
+5W8EbyDlriblHIYqdwB+zHwOt1bCGP1TXTMGwylMoSPLZQECC6e4iNXv6h3gQFB2tSFP6d4XxCu
owFOOFlobdg8A/A92PVY+jKzRqVBvL2cuepeNNjWE0u3q9H1CnH0Egj7ZW55L9AUr+ClMAwANjIJ
wA9EYG4FWSPiyvRo25X8HaHhQNW2GbdvJAJDc3urfuHBFfftnK+MOynJUXzOWE9ewFRFw9wbyysP
oSVzyWHj4/HEWeHpkSxOK8u7PQmkvp5BRbCiXw6IkjiWrKYWOlSt4Np0wYegW2FfsLA6mZm3NMDJ
++X+dKTaGU1RsgS97TJDtzwbJbJZWbm8kF225trP6kjhhlLGskzFAZ1hQkUcN/klwvs1lpBk+G7z
95h6/t5NIdgOxv0WkIgfjzS++EPh6Tlh6BdIEgQl/7BY6i5GcoXIdaPSZNg4c7FoW9Wack38vruf
FG+OqW+/CBUw6cfIuApI0pPhdpBo5OP2UJk1I6YCd/PqF0f8oAoivRjmbvccpKDwfvFzg8GkMssq
D0XwHvOQCOnJHcfwPRE04KvQF46pfI1lUXsJ4fRoUIz5tpN31dNwyWfYzX2wUc0AWD6VG4U030uc
izoUhQ1ksKWIq2CTiDYANoDSZBzptwihZXcmguTTGmncfpvhr80360E4WFhyKvXEpq1+7LuK3FJJ
9i+nWyosT6BxYplP+RtPNeIfmrovqeBY4U9xpZxWjUK3bjbsHIdUpNJ592FmFqsH+yIkSdCd4qdU
ObthDZcS77eGaTJueCrzJYdSO9aCKLr4lAnmk3ArJYovwVV6OXmQfbrgsJVCIfDdCU1ShqpmlUY+
mTb+tAhBfu5TuMnwUmgPbMTgGGjR0KbmHLcqM+xO12tnrC+vn4tZZMnL92iDukCidqqBqHuiYXV8
hbEJGhr4gV9a3KMbsolKO8wczF5LJ2B1WNYLn2iJQbra3JZDCwFHrHmt+HJj5J1lc1jn8d1kHtNU
KMGh131ZW2uW+9a11WqHN2wxlaRO/rBt5xV7XJdyD9hFiA4a3sJ5rGI5Qzu8yZLIrDJSoXFsLsj4
1BZRuZ7mHQe0EFPtvs9Sw361liD28bN9TMW5MRm962WI1m7kfSXu/kkGH8YndxEanjHupxSu9V5R
0F4in6JKebjKEXwXGvX0XVykb1oI/9YZJMiTW42A05RVx/3eqQrx60LUTNy91FMnYqmmr9nIoSVk
RGvWmeR7EHX1iCSUJLPC2RAssj3v8a0B/WXQDWO6he6iv93wrY7Yuke13kQ+WmZ+b5SQbZ6OL8ZA
T0mrGA9o5zzqqYU5cHgnW5UjCMxzQm9VBEJlOqlPRU4tgniGdGECZig3F5fboUZyTNycjgDnMmL/
t5h2UJND+fKwNmVydJPhoBplcmkEJmaDp6Pc5KP91qKNkqdFi/ymq1Xk74z+09OSiFO9s7YqTbYt
UfuVmDKS1z7DMEpTdKOak/G9hgOGsB7LMKz7gP9t/WqCcg9RP5ScfAxmfoTbLExKfKXxZrzmDtJE
IQ0ofoBQ/cbr0Dz9VthB/+A5NOk7GbCqxv0yrDzNmgd65D72EGvB6WunMzmTLwge/+SqnaqJbYCd
maQ0cEyP+PlyHhrVoU/4vJWnxalnO9M6iGqyWSCvnLl69424yxRbW6sqfLXvp0fZmXUUHS4RPM3/
jcL8GxGvIeylpy+EoGumKkvEDKkf6OSCY4wla6mF8dD+I7OI/unujFAcp4ZKT4g7HWl3bLuyncXp
pQci01bAXarg25W5p0Iyadbx2zQclpzd+9TfraXBAZmjBhQ3N8Nmtq6R3eWnynVjAuE7E2TSF7VU
LQVThDlbrng5bdhRm8jLni6zXSEr5SeXtZP+7xCHx0ezRkGH1kKzQ0/zKZo9efIbg353FogsrPcp
6zh7f1fDgggKqRxQcli7cz1DKPH6i0hPcb4JnaEKTa1CBzMP79PeFtA5GzGjYH7Bkfhw7FAFKMuP
YKt0P94yhcpvJT27WjXyJJYPtHSJshXYEjzIsMdK5xx4zy5LuxuWJgkkXN5fbx75AjPfIDGofAu2
Z71aixJXblzEa54QtFRt7rQ5KKMEJ2ZoSXp3SzwOMUR5HfASwecEY0P4boptBKupA1Fa1kUhy1Ry
U2jOq+mPm4aT1qikJC8tCnBZ/7rMvevJYP37RQIoQeIfpX6kBLUKCkWFhTyo8z+s+M55YiK8JIJn
tHTHzDK7C49ri+vkXtSol+hvDFrOX0q4xm6YHAAeaLrNHTA69eLmVU6AJOebPfy0CdfkcN5YTw9Z
2uSexhsalV+GZWHzcJeBM07OnjH+8PU8q65HXPv6l/x/Y54ktIvxjzzYRe8fpwE6+OriTEmnLFVK
iNmskBGCPS7PMs8aNoWvsLPfxzrDvRstdm2h69Q2PMA2uHf4nz7wzgs2CXGWgsqUMYUsuRqRJFYQ
1AFF4vrxnugOPumbahYOBDKr0j0spEzIFeUAWZ5oT0/nlygpBEd3myy5L4k55cO58IrXeOLpJw89
5oCyAyf8PAieNh4OPIYxg6KxafnEJchBBHviCcdnkpKPiNiP7IGgW4MyJtBS5T2MR8RuLlyfsPpB
XoajK4bchDz13/JZ0fQsEWwQ9Pk1hs4nwe+zp1Aqcuy8C9v6z0RPTo7eWREcQtkIDzuDeLWGy3K7
Nhiod/NNwFNa+jGAtqkM0rmKq8IxwCXiDEgohxmaU1KXbZtLNbM5XpjvFmDfn8Uvq7nyFTprusZG
AcbqxQSgZ2t7snz73MPgHYvlAhFVTkVKVuXjgshd7Yxj101BIToPy5KJ2WBYPBa57os6xzBQ783Z
7hllvhnqF+XqQqPxoJu3WrSf22vnTBRMJ0islj7pQh2RQf47OPVO3akVf7U1RBHxdymX8va1VFSi
aYD979HUXoL3LJPwnHSrHl6V88/T3qXG3U2YtDPy27KDXZguMbANjwjsu1oHPIYwrE696CymXUTf
o/crSfSukjquMaRH3Eg9PGr2uJz9IGeiYMAUjPpVbmWouRabvBC+VelRNvJB3xTOsUiSDoIthLP+
svLcHjxZRKoded5bIb0SDG2q4eG4IMtCq3y25NOdwPNkfNa6d6+9YlKri/hmRLPq8wUrwOJGkj4c
idP72mNXNatwQn//i7902ynIrJNfgZ0OIP6bDC7P+27E6xoBw3QtTx61jHxVmNz3TbnwxVDpv3WY
MChu9B7XTZ8Ava9x71bTUtQ+u7yLWw4ESn7hyb7PyompoeowbvAMbo793g25XqDQl0b9Q3jUOcRr
UlfkbzdlBYLOAnFp2ZG1MSTHBbLkip9iRDLYAhqW9Ox1M2kriOsP99f+kGVpAwuP+VAFPUirUEjB
7fr17M/ZL3B90+68+1svxxWzPOz6N44keG7QACzPLKQsgnd+kCHIJQQDjLSNDMiEek3FTdsvi56/
bGZwrehMQf4QJYbrQ2TkZ7UApeMXyx/D8MnFJ/Eh5WVv6N649wZ6vTJM5im/I0WtHkKPvEir9C0a
wVw6j5+B4WbxrSN9Y4IfIS7txqOru2nK5hHYR4GeCCbK9pYSPb6b3843hU+jNTGQwVLViFXUKPFs
ItTeedTYQK7Hu+Kdd+xIglsq0UeIA+PvRB/Nq+4g/fYNkGfE7tT7KWznBSFdbIhtgN2G58ysjDaz
IWxdttjNRw3ghVaGY8HMKtAhZgPHHjE+QUYblY6ufGMfhoTdeGNpJujSnumbJchGDuH0kwSFnJVl
SzLEo4L+yX+qJLWpH8RnOi/iitdLXzUcV7lNdweGELEfkeA+SdJjtCsrkgeSwuvt+ZJoWYKsx+Pe
nF68YgrTFl9N9SgBa2M6QyzSIvMO7sSs8sNuB2G1D7fsMqgCsD/9pkVIoHHwvsxlyj/p/lo3xR6m
kQnnWXNyW77j9igWG7gbByZzSgediD+fgSwd3Ioqt+HvGaEAZZ6w1LLdML9aYvw3XWmn+3xdIaLA
VvydtERFKBExgnwD+EVrK87pE+YRRZg7bHudF9YBLnvu3IVwyCoDRLp6SZvLtbkED5IRoXu/cSpl
z9D6vdGTx0IK4YdWtYwFtjkgOINtZbDUqvmbJn4z+kgQtZhOK0y6CFtY3FumSRRA65d6H3tVdENJ
9NxeijbjU+F9XzQLwkYicSZCg6U+iT1XIzkuoUPqkJ2t4u48GQFJwjeEQ7zhzINgTuq+zaN08O+H
EFe7MKR+W5AF8wXEeSVKX54lIxqhlhPPImVYE23HNTgP3ynLTz220F6pgwcUEy35fi37N9sEDAsS
f9yxcBUoYKc/5Ca6RNjNq32eJpnpjnZqabOO6YHyQWwKqPCmP6ynv+UQjgGh1z4gSw865t+jUk4+
lQNZfWMKqHTCEa7lGpEQoAp9jwQiujW/rQ0xT2OvD9qNH2hpptcwzuY/qMvUmw0tglq4evSSj8wG
QpcAgufHIq5H7TLxXmJLXoX3vtboo2/fcpfjwShydYHgP0n0kjuaFVzvhBjsADKa/ci/fPNTQohV
zyQa+WulhXXI4wKFo10DNeTftGSiBwX6fp3f6wDJg9oqPMk0BWmExyPqnJFhqn7jupZ7yd/OmEcL
xf2nGydVkSXFBZFXn4lBSilM9LGrie+VIgQSVq8ZfMuIMP0+zM/na62IyF2s7C4czd4kbvDaXXPV
ZmMc+yPWGpkSPtjmodMe0K7CtCWOyZtySOIfzS+v+B4jiATXmbp/N4j/Al2p9nrmwCMkFFlphsRZ
tf9vyAn3088FuI32f6yNKKueYk1fhkDmE1XobUz/hpP8SMqL4ev05IY+MI/HFnUJ1qMCJp0Nzh+c
feN/BYTdr0+LMKVZfK/bbKvzr7UbgesSwWc2p46cCaMVkgvHmueSTU18wdJSsQwhK/r0eH1qbliU
jwUSjHeTh9JhM4wHHnGo4jlkmoz11TPQH4wf2I+CR4C6qfRd7FmQuRJuZHAOOgNGj8+ggNFHOKez
g+uurgnpY0NKl+06QlF/2uarMuOG73ipwTqhWT2LZJ8kBQtGm0xwqgi5GISQdWM0qVjLkf5mXP/w
8a6V1xYW9kMk6qpQLXm0SjWolip0w04aXzeOZ8KBtZN1GQqmj6Za/Z7fcOj/e+H5kHHjl/ddFn2/
Ky9E6eYEwaMoxP4Hdh5XFRvPXhL57u26hUyWAZ3bbBLWTJR8V8Mh32UH4PIa/z8uKF2Bcq/gkXZd
Y1Jyvrxm8XNM12G7AtNpfPaoth9T2TBeqQFstKa1mQltAklo2HT6lC0/nTZva3f9DISyLvtvGSx5
Lt4QYt6nwodFuQSHq9sKZ7EvHw5MfPNmjNeWhf55u1qC8kQQicHlkA7x/4V04+oxjBSIshqT1nsD
qwZTGd0YC+IZVZV//02bZ1N8/324UrYKxtRPQxBX1joE/VFkEvaFUw/cmolPzrf0LHcSkupzanb6
mZ7YQJqolh4TUvHOJF9ySDihfBxhuRjTeEap1lZ+0FLn/+QEyhqxN4tEMpAWZiAaZlmYw8S93bjr
CQmQ2prshfNemHtRMN1RjUmNZNO//TNE1RxpLSbVWjKmNkqBmEBi/aXNWBxBUJkIhdaK14dirT/N
6vMjNexUUsCe85C9bgGZ70LFw8nSayUW2tpZFAPvbipcc9opDxZMm2zLpZ7RvnCS1DOJ/8uphVOM
hVhtnnqcjw35FhpkGWVxH4icqTUS+9BJG6D7YDmylN5Ko0MrqAyxWn2woVY2330/LNrtVYVqAyDa
b8D1mKNm/kmLtOHE9/Pnbn8rvlD+bptGKTfqAs6WKYW9m8le8PAETMlsmIeJcW+HXTxMaYmGZlSV
NpkYG8mitbXhd9ehc0Vu9BnTWubLmDutko678zZCmr6Vv+sAjpFe594+06gmEWVTswzDCCvIJa5w
N+ms4w2CsWTD6KSNayv8votjjlc2YiaxhzQ2tGiW96jhMet0g2y4ZVks1g4jOYL/V1P4lcUtEwBM
Y6bdAwDHoly+N3Al6lEjB/KKj6lhexRgIghIXzvgo/F0ucZEQnS4dbV1Ie3LlUUdawUQ70FoMO5E
7PypSGce4wdN+4TlHy5pCx/WAiFfvVgpI+gZ3daygwaipVbYnETsSUvIdOoqHVddjA1ZHDCOtw0Q
oFj7cazCnNm230ab+yRqDNskMNl2E6oVZgqhRVFlPA8pSADbSipQULQ5Jxh5HcuaAn4CGLxTInt9
JU+lYkyD9ykkeGVzEHyXS+DKsRixiTN1xz/yhfeYSS1m4IM6cCEZ9ayEt+0Lbvibp0GHhODNLJKg
5ke7TKPBwXaWyMSvYnlUqVbLsYuqKOXuS5hO467nhti9V/3w0krPkFmEwTvLWxbvPrp9bayL6Q8K
t0L96iSC2iH+5cq2Rar7x1JeMg3/iPF1UThQXdGBeSXa5xkH91c79c6fkzpmYu/XczzRSlnBf1NK
iPVw10TMFm4rHDrCYcdiyiw8quDkU6ZWHS5Ys4/ZpQXwD7JWcBme6FW10a/jCo8TATJxMN5567XN
F9Bv3pfRjJf5MquqIhneYBSmUfDmGnBQF480YvoRQXn/F/h3kFuFRLCHJUbLsmajodKRXdb+7VIv
yGHH5KUUE3UqWnpUJdrOM0Zo2EUAkyAbD3kLXeUVrC45xPy51GAmmtoTJCQ1PYNjP7pl+z2wMjtu
QYglXw3wfpwQz5dnMYcKXRnNB8Av1rCrie4ap2dPEpnwpT0iOyN6h9CXn1lL+M5GZAYybprXJO79
A8l84RSe0KBLL58j3++eFmz7d37Ya88AJGhProWRmYbBws4jCxvkP+0ME8rMWvPqaAdlV5Rriq5c
HYRHOTSccCHQHC6/2uorIyYEyFm8zJBkn0sN30ETkN9hNURhg/oYSg9syowL4MSjwjIYjBptb8Ps
xkWOblLy/3X+Zc1vJhJ5v+JZGcMz5zTbsj+pIpyHAln+nbGTiZ/6VIBE9b30PiMRAyuvakqfirCM
fsazf1PcslNvupEWoOKw4Q3hRzwC73NnvIYuvSOrLW9Ls0iMnUr8SpPc2guL9ve+WhLkKd/ZjXuP
5r6T0U00d0lV3YYWfEy0gmk0FzxV9O1/bQvC471hJSvWYNvlinnUDd51cGM6sC7oTjscFJO/xJ6B
ld1k3mwb90PN6OjJRQWfQz8jTVQURQ/SNWBup8aIN/+3qCWz7/EJ9KPd8smYr6HoUOxHDHKmwSWg
VRgHnADampIZ1w2FV1QZZDgTfM+Pia9+duqGgchfasQg37u3hFb6IVMfYtVlKfbBfEI6dgimYCXb
2RW0gzRATYIkbvJqGsKkNpKK5WzVtKZeDxjj/6HgtDR6rLjjSjWu3yHq0OdpkF11g2JAadMWBrsG
jUvqnY6vWRpkUblCKC8+nYWw9S/4n+ujeJOaY7RxSyJXF61JBZ2L1LwMvjBd3D+f4feuX+nwr/zB
Rs3qVvVvhojVwNXT6rf1jQahLIHij+45AfRVn5lZFFDxBOfHTX4u7PUQB5cD2CdZrbca0ntDs8AI
QRobbwxZppqedZDKGUN0RXXg8/t9X5VmpKCWHc1h27p4hecEBQOEYJqGA+URU8uvUb4mu+eaRiWP
Os3QN4pR5i0A1+COTVEpwX/lVor4AzpqzZFkbLvEg9h0+cCsuVR4P+kK6YXxm8QUjfiemU37HEE5
aRoNY+DuU8LqvJxUR58SgUqz48aAizmdw+17pPqDiurojnFmYLkG4NxyHi2XbZOieX28b/oY9doT
kAqATG8OQjsgFF7yPYxDnojeNBTXWKkKWWy+cerkpe2Dts1DquukhgGuLXiBmIdJ60hSxDaR/APs
Lp01iDY2OaYrOOOmnCF7IEJufGHNgMFbEFFXQ9CeqHFQRRMbGw8D0/4oIs1DMVfiPT87YdvUwr1g
uI/p0adSGD1LNHomFrlfZrSoCwjQssVdTPFTd9FdkGfuInm49tvcyD+Q90oblOlnY4FprFosTg9m
cM3d2sZqi4N3DvSCZqthvymFlAvuwDEsKQUynsDxxnOykubEfZB0X9NsyGRVS0Lo8tmuLkhkX7/O
2Xne/MvanZX2jEUQeZkuU9Q5czLEIf5l6mgad/nassR6pyPpyYcNhgysafDhl/wBTMC1A6D+IASm
orcvBrtERkdAnyOV497Meg0xfhSd9i6B90hWVJHImxjUY3W7EZEA4OHO+B7Df/pJWCQD9SRiW3Sv
sPRwhpxSXQmx7HfwziGm6r5f073px/y/aPubFo2At07TWnlrHaO1UyCkm7kh53dNA0JDxJotUUfG
q1ejWaGf83Mlzz4v8xqD55iUQSPBZmuMtDeukZAz89ahrXMo5wvEBxJ1u8zHdnGPra2ZT19uLdlt
vy+EgF/ViZcCELTZj+htkCmcN6yfdOTxcS5+bPW1cwdI4xUDI7kJsL/I5Osd427wka7mCv/d//7l
tjdt9+mpyTzHulgTKR6ZkhQ3LN9mKBfrc8ACyKDZMXbfYxNsAMIPrhpUuePBJhrd70DyG3q7EgBp
zyt6fy9o164PvX+FuQH818LxHQ6sNthlyWtk2LfMw7vCW/DFSaQPrg+Jv2Iw66PCFIAboA0W/IZJ
uFZMU36vKZO0ftD6y8HkmEE+Mm5uBJ2hY9P2UIaW91RHuSYsN1aiOdocRc1OZx1ArNvlXqvabist
uPBfmwZld18iMfUpx3Mrc2k7Z8TIfcW3hdy59oQzMNw+x/nkX2jSZV8L5Bt07hldqz6QR7vD2bOx
x7+ayiXQUIO913sTjin+yIN8pNsidz1brNBuXfyVG49po5brDtOPT9OdKe+if2humNeR1fpDjGlo
7x7wmecb1Ystx4PvBq4k8/nNx9g1AfVDMI0r9tPhFjPFQTei+XiHrQKL1l8zPzyi9Ln1i1gsQqLc
+SHHIc5McDQZWY2QKTKM0h50jBmHnNiEtSg8wnYhyjmozAu/+s42mVK3u5K3kvB+gbRsdf0P/k2K
kKxNcGlMmvlu/W1A76wVcJI+hbqIvz/6E+XpuJ/4p+Ul3P9rxp+w6gFAQ4ae8kWG4mVWEkK0Wi4p
F/ZR2M8z9hTpB2rSzv/8TTdqnj+e+TuDTapyHQbyGXNf9mL9fRyKWb9Ot38P5MbXvS36lZiAMUfn
z/LiVkH22O6DaEKzncQiWLn2UiILKAqQApeqvI5zBXVnpPlbxhzbiKcMYt7xB65/GoD+znubI3pU
ubwvPPSy+FNpFW5v69rSKmXrM3Mwk7WOhMd3/s8EKBfjyUOXRCx58Wx3GYZRbmsxgOYnu3unx48d
epr1Cb3x0NVF4IFpnPsv1XT2UoPc/Gj6YvTKuIYFTSzA4huwWvUnr2OGFc8pvbnNKdhpDMi2pCK+
BX37X3g6hgR+tu+pxWYZOjDFlrGTH7MUtMQlnAq96EIQQYV1BoVdeEXkbNRuPytOQ+dLWwSpoLLx
fwtnpYnTx+LAosCEV5Z0xj9ByXywEPro8FGSe0QsRuD/mjejfeJ7cRE736VvoeRHPTK6vGfkbTTC
4oSS7fsbvvaVr9gAW0g2xajZp7XI9XUcesUgFaomHOoBuAUIuZuf+XqHINQMDakI+ra96ovKekpO
mOjH5M4qIRZZl1NAchEB+4JwgcfHEf76ymy0X7d4jA9Sf34o0gmsaGrNsMNnslSOv7oVCQ2s4Q3A
nI5iSLZgXwdCIrDz/gxFczbCVYdBr8wa4YlZOCL5Vz+12uuoSBaXYQOt125GTQjiUUVnO0BSrE88
PgI2/DClFr98oAx/lhm4tjkO3+YylqmWFYwK4aEb6POiVAFq0Fjar8T/9ZJYtBRDpfJ1UT3xXEBb
r/TwoVilmu4FiuX7/QwkL2sA7zKUPu0K5CITjymqLLdf/QH9ZAb3j7SeGZKouun+XNsXBbL5RgRi
eIOKRtBhHmzRwjbNuxNYH5XYy00EK86fN/A23M4p1VK7IOdxYIs+XqhPQmLgoU+aKAR4A28nvHyH
gL4G9iS0S1Syk4u4drjKgsxkdQCCy48TLlz1RGmBecSSmpZqpuPMdsDCTUt29J090uvPff0xRNjo
0kEJ7Dx2zmWXTeDo3uUSXtV3qDf/hC9LqTqEeoMWPIhxHfwOC0P5397FrxHTPq1t4IEDq+wfWl8z
xLpicvN3hZX4+04j/U+m0VKqIs4B2cl65g/W19D0gDsHQr2QtYwaD0Bnh13ozQtJaCfAlrVMouVy
9+HLVGKzeIMcClc6jHqDei+KNHRf/kUhTAhGdB223JmlHlD0Np2wvOarFjrdH3AAIbBzoWE4rQ43
3thon4FnE3WLUDtE0KEZBDr1BUSp0Hw7QULPkUS28aJfFQkYMKiOmqWn4fAJ4AnVTS7k/vyWJ+p0
5tkxk7e7SzsGxwzt2HB8smLnQjAWE3f/XUlCLcFNsADxRvmUB/p1+uQ86r7fVtVxCUy5ST6PKZB1
VjOe6+o2SB0ulAKHpcUZqjOYr+vPDD5AW8Yp6M3c+haQ8qAhpojJdNnQ88jFNm52N/06C0P7JXpT
G3vUfD+TlxQaXJu9U103NgdZtQD24cPiHQhjsVUx3yfltZlSBk+TlJlWtqxpVWBrIXhP8mBPXbR2
n5yuLX99QzKkAGifXa+yE/KlIfLkF0marjaFLQL2uzEg3K2IMmsNZSWV3NsuX/QfSVTrAdv7bcPM
xpz0QsoJ95TKVdsiwnSNJw5AxCclxluvP0HxfLwnDUWK7TIdC+NnD51H8UsEAj6fzxEPLr5eYjSk
xj6dwu1VaG40bzjLK05ni+nU29gOtE7Hx+xryGTROvXKrcGKB84CoPQ4tpotZSAWUHqlLTgTxTna
+LM5c7QN6Eaj4oILNs65EubkteWRWdNU83SjLDKVUd9vcIBqHOMul1mZSaNRmPn5QiT87cc49mHp
BFboJsXRUPCWYU8I4M9m4VJcmc8RQyaDaNoo7m/DSBEyclhOO+uhLHXJ/0RQiPp7Hhhy4EM+iZby
O6gHGNximHdYN94MC4eX3+TSe7b8kWLdWncJFx5Xc6n6w7SMPqMVhEHxNhfVvnXUvOfcHwqKE4lH
6DVqO1Aql0L4MtiJHyL1eNHPGc7/Yt3cVXBGfoxNLf9hV6l5NwfWsrvyWcjgSA0ZGvvGW9ehvzBN
WNygDAw6iHWIqspUr9TpcipFDg9JFgtF1aCmeVvx/0+ReayPDfqQuV3CXbwytQfTCXd0LMNkrUtZ
9c9NKRHsaD+2o90Yr6T/L2j+1BA+9+oS2A02cuIHiYB1Ywhgh65FYUlB5j8WFY8+Us8wK9jsWbCJ
i7vHp1CGZc4bDx1O4k0szw3/8S8OFN7WmT/OONgYhsYtdHSY/pqbiRICISMErO9/FZC+5m/wCt2G
1l3ti6V6UhFv2ieQCwJsbMuNRsho5OM5Aj1ytF6stsQup94LXfmgkoKjPe7IDQ05SRJRqeiImu2X
iUxpU3UDCN105Ge0EjfQCivX0rnnGp7jKcvLy2d8R4KwtOhLTNuCuBKyBD5yHlr5RI/UKT/fjg81
ZwmC5enFaWZRj4ncgGKvtliCDcu8VQFzFWlRi8a04KnwX8d8LLnuiudlx7JOsfNKZjtJBPEtCvmG
jjqQsN/D5qXONx6H9QLsXJZffSRe0HyiLPOrzLgF8vThVCgFtMI1/QxXWxMvZDBM7i+bMkCMs4on
y/ELbtP1oT++2fTmexZ+6V6iiKRT0urz5HrzFmjx4u1lsi7LUXjCv4b8+ncSj4Gei42jjd/4gvXC
ZWlaFLkH+YwoS9wPjd9qko87GiB6tMmL8yZ6KrFjSI6QnS7S1BTcugWti25gUqxlaz1YgdJB3t7a
CfznwhT1YKKf9KsrKYyYZdDb9muEjVdRbCD6uiYj9Cpql/E/AdMVzMAX0zHQcST5WOCihm7aK+XN
bmB30lj3Uw6Ki9SY8253iwwBV57MHmtP2WYGHoMv09V5+jQitng6ZNwvpa9yk6udt7zHCEnAq4Ni
gXBlxRHnkbkw8iVnJS3HUgWsrYwvAimCiXahPEGq0rr/5yosx3Xj24CH8YeJupP8FmUpXk9Y1V3u
ICxNu7AJ+y4BTpaSDrRdsA/JoF3Esq0IpYfDkgqchmXtvtEFMDio94d4ppGydeFS6fv1xgn7XB1b
rD2RirIi1E26TnMOe44/6CfICY0atJM+AOUp0lUPihsK4iMH9k1Kbv1HrnR/bAdxvHhNJ9ZBuOLc
GgoOncdfv9goz90G8bhV4vAh/nfTQJvgo1c9ONuPr+DbYC605Iy51hkt2k3JGFk+/n+RQTcw2JAw
iCxn1h24b9IbNTQmUVvVHPh+ol/NOTA8PNlRMOm/k50M2f7manupXsCEfUGo/eg9wxoPvoHjer4v
qpq2K9pW0DYdG1BE7BO/mTkpanhyx+fO4ZPT0r4qcq9tSBGPM0d2UJOfUSrYqD8kGqsn9UrhUv13
bPmIAF8CjQzDiTvlc7cjrzSmhoGholxxbpxOIzlirW6eUUjI56K15WV0JdBIeT/c2t5jkchEfXis
JDMqkteL5F+Qn8jj5e4aZtk6zSgF9diXxYiqaFP4gLZSr32kcKuCJv4RQ8sDkyq8OuhshEKAu69g
pIJVopLwAr8Vo1tHmxYEtWe2d5GT/hlV9RqlmlmSCj7hu9jYRoXo3lBcEOJSU0HBmh+e8aHOgYX+
3pLAtnkk5h7tFLYeM32mOz7EHZDU/JYJA64M4JvAxHoALXx4ESk4kqUWfv69V4w1finzBUIb4148
0KwAgbqPUUvO1J8W1YiIE2f+WpMTNfmypixzg/E7XOiWlt0+OMjlvvhjsqjl6YmEke2y8CdgUwzK
/f/E0bYBZgFzVsfU8u6aM4d7lSakJseuzqMzscL0W3Gfzh55PzFqv4K136hfvJLOI5Acebq0RmhI
7CE5euMkpSm8DnWO9bY53lea3+8BOuITT3fHYDDSp22KdDQOmTRwYyDUE47RqWoz+/uyvu6v1OWM
Uk4d5uavnCTz0Jzef31CG62mD+Lij+tVJ9pEPOLr74wWK6LE6FG0CRydpP1vsyxckFJYNdrq9cEl
X5NSiBO34jwbSDqfZ5h/QTgSmX6HQwF/zU1o5BZfgrvxLjeZkZSDQO1EkKUdktEUgK6paV0TwEJ8
2+lPGX6zoZJ1E4XgFnU9s8F6hq1GmATsA7nmCuFKOBLo7z/3D8NmxTSXRX20D95xxA0tOLiMUHI2
08YA5dc9djPHz/XrSLc0oJv0RGmd3QnL+fJW2Y5iJM1ywM694rfpEj09Xh3GDr1GQLZWaQK+5G11
olIHD3Lqtx8U61OFedC2/7QZxIAz8nDsfAnPUKWIfiRRbOh3eV3hHCagS8z8AALsprZibIS9dO3Q
lTq9mRTpei+4v3i27x8SNYRpA7iIw91z8n7VTNvTf1SwN0zHpquHmnGOpVX8ZkACAjigHK7kAmzw
jd55cYauNkGysAdwHZrbZCHoBMsa1nN8RPpnWrLFTNHp8VDWVF4+sVGQbZz6Vjm1mAPbx45rIFUi
LRO5CuYqtwpefyMknvxNd5d/TD5VrzlONKQjxN7R0biXzzGTDKcTOBicW6rz0lBLM4XATLDuFlfn
G29t7nNQ49+w9VlN7bQOUHsfMAia9A2BkkyPK1DZQPC5bbvpWUqbneSwJ/TI8/ThEMfU7y/kQWAc
k57z23Z9vR8LgHasrzzvWpYbhz3IUTcxA491O1lkg2VtQJCobs8CFnsBus2AcD+wJ26tRzZ5ueGy
yPRSZ0ue4EWhEPStmtpHVnJWGaqt6lbMGzqhH7GGI7AMXe26+JG1MPJk5BGeClgE1uc6+XTMaw7C
sWqPvSaZvo1hHDsrcTSspA9qLld1Gx1CVyOJX/oVkop1astWNZzHQjk/jlc0L/FuRoL3p7KLHPll
A0yMVlw6jq+U4UsXf2qM0zOoezhe3drWMQy4N7D4GXodIYc+6rHd7SoEQ0/ZdK+NvHZem+1HtfJD
yX79seqOP5+VeuvzJfTuS0CrSKznNs2FaIH0dYsauPNUVA0k5n+7h9JcFR33XXqZ595+YsBzQzIm
4LWwAKmMh+5JHE/2VtKVTvj7dBDnP51N3W144sUrBZeKQGmFyuyA3JzApUqEa/x37C3cXCsxZJRv
dr0iBIB69AfHm8aRLbCzVJ9ieKUYylmbRBLYO7uUfBbM8tw+i6X8ydWDnzSjbaD8OhuUHv3UExKT
1LxNmdXtriXIZ/ehezH6bHa85hKEO38i/8KIZ6STy8B5P7Y/oQR3C2vUxdJrdxRd6uZ5EsWAZy/M
wIqraHQ0UCKr0MG18MeFIuWA1+nr+0kMiu5gnhiYyqfYc0Ej4s6RGeu5YM4nYP07M8ZsaFR1WV38
m2ePRn/dlnpGTGpk/ptfHYC7YoeTt0G3P6CcDE2mAQQyYp3AG3MM+va/xt9rVFl2mfA+/26sLA1X
BuiG6leHoAlNZ7a/u+T4RnT0Z506GiH9vz0qKFULQIOnkVuVA+ZqrYUgZ9VydcZgscQ8yo39qRL3
Jv3wEdc/HM7GY3sk2hnQzwlmkHwXPHOSk2csU6JpYC3yJEwgMP3zGqElXNRFk8nIuh1tgS8l8ePm
NZszLLAWboCnc4JFy3If9C6PemMPKejD19zHupcQ/rI+qKMlaSCm92zlM/idcknKVQgDjqjNeXs9
2tLs6bM66+eTz9tjKWd33kneWzaXgyG387m6NYm9GtCqB33gHH0q0GaB55Pe5LqP9Ps5jeBpoN3x
/vfig5etDYvnvQcFTdk/DLyD3Ge6wt8w0tCOavkbmN+STeiwG2WxKL6EGZweA0jPjrY/xydLp1Rp
236t7BtUgkY8UxVrFJ1RoB+gEvTacoL0ToIuh+7Kb5ne8sx4xEzMpUN45dHXBb5goQYH606fKTvU
SxABjbK6KNut/sfP1/xAiw56ZKNIELrW4Un7CRw9HVQAxnMV/tP5ZCmUqrAyRo5uXke57t/kAXbU
vCJjbGsRLeXjl4lpbLIzcvNgNIhBJVJ0HWOXO3PWu28k8hFg2Sf9K6sIHdTUX0PfT90tM7x+27D9
quaiMR3zi0nIDP5DcWhZPNSndKELMDVP+XdNYS5PmEUNT7GVdd31R6s58C9cfzl5x9MKFkT3f7IP
9cdqWDLskSsab4X4klQSkRqhG0X+1P3DNtnBV1aFlOQziMVTFMcuBiamxA7Lj1ClFeta0J2f33Pz
eVX0tHSBB6hF9/xwQHQDbCylS/VkGURkY3n/PITIalv6CHgOJvEzt4BPTM/8akpXz4lBwWs9yr3z
cU2PvFfa5D+/bgDmZYmpSyC2YCOe7PFxzvdTpzFtQY/oMylOUpmQ9o4NBy1GsNUWcKiNPv9MbrKs
8pSu5JLJITLSELf8lCp1SPjcXFwI5Q3Dm4aKd6SLutj7DY/2w1LvVqqVlrvwHqf0ZKQDpOqkAQ5d
SJnEwV5RgaPeTfKAx+/beWa42aavyceffiG8oQrLP9la2OurR5rGWz7p11zLBlsa1QmKXcitP4Ik
m3/T2QkJaDhwHw2dlg1i0/SbjRbfItig6H2/skJyu74RVk/EqLYTVqSp8U9taWj1WQCp1me4U8Gn
1mDtpTvIKnVZztTAWH0YK/ecQhIfk1EinNVR6kNiPBzvFk4EYSEO6XNkrJn4BfMVCAXSWkubfdzc
UiIYj+SRwOMZvuBmmzuGd6VP1IV0Uw1fM1KSoSutluCiRVVMTwJ+bewKFfNwFmVMtUt3gSeWbIi7
d/40VHJgS4wycPx6B28gVU/FmbWMzwxKffVNxoHAEaNCQp8h985wIvwEKY6RzmojPLq4m1mrCwaj
p8Xh6Vc+QFS4ZJoALiGgEXh8cbjui7xMW6t8ABIzjcpwfp1JyvcVDESYfXdQv6HmEGlkR6fy7av6
ev/IQvc0D2XDMrlElwViKgFlXWUm44hh1eh10Slg/k9liHDQSvFvTnPd6hcA/ijVUENuXMhkGBXW
AQGw+IR9z5a5saH/ovIXg08H9HKcMWRa8XVtLs7KETarf/FxC0rzxUl3BHi4Fa+hsYYt0sbRZyc3
H5HGmCP/q+PhOBoGsxNlK/sJ8b2J9BpkCUeoe49tEWyOf8CwZsXKX/Svr1nw8mAuROmPZWV+8lNj
99RFOGqUxpLhTsnxj/RL31NLwUOlZIkjoSfT99OXqs921SpNz8Nkb1mZiSP7d1M7EKMMesF5kXWc
cGMeJosTRds9PcUPDLxufzkunh4SN6dXCJe7IM66Ez4g9rzfZx7tFrk/xKoTWH7qmvd5f9GZQyWd
ZjOvJ5l7P+DGjVsQ/Miq4RWFKlBCyYkFZQ7kdXCdX7TAz50071qSf0dC+Zmr77SrCWOBze5zeGDX
9RTOANwrMvTkCtKkpQ0v4CKxVh/cvybBrd+Ht2/BFd67lYDFUrNqjjXXJeh8guXgQuoY4/2T0d5y
VVE9KBA76xk5LpjuhgW239ukv3rSHKoliIASmX00RZvGgdO2dYA+W1A7PVyi/KUFFFyjucX1BiI+
lwpLXTEmp83BLGwhw7ESYWXIPoXeWDRKpJh1ztVz5g2GGl7xDH2GAEKPSSsIG5sGRwrwXBPp/ghj
JWBzkafJgtom5rL/n872wl5dy8PsZd80XrGAN7JYYYWfzzIKHxYfpeszeQ5vMMN60yug1rFf+h0l
eCC9v9hJLoWMnjG8HKNhivicvx9Vq+O+7W9EAYNAVqahRlw3XGwnk57m7elvkxJIJF9pCMav9rOL
IA7YvDrRERG4/5ahpjmYpeMGg38te8iKX9YuSAuzllFXwpcoVhBrLKP9XlKeHDqCcivtOEzIPZ/Q
BgCbYNzhYMssryKFGY4FX4O6Lf4BYnUUyPDy8z2uWNhQR54lYxiUedGDhrvESzSRfV/mzVwE+jIz
+l44jHxPhtKV5K8Id+XUgZxmAA1X4MZxEFYqDUIfNJZFwC1Q6wNJuNTDHFQDBzlegL3N7NvBDTgr
wVByKruljN21dl7phuPpPfqhylUyqH0VNR6j/B9QbqlTebMlXeVuDn9Ow5BPBdCk0BMwvrwJPbLN
9V4Xbe/VRXrdJ3syOPoO6BhSxMzEU6x1Q1xYrQ54UmewTLScHXcq3oEUaFCVJGq6AJGvGt/G6D/U
/6ZWnPVAUsA5MD9n2qJC2SessaysqA8jo3MtOqMywDiLjKR/+b2Bzt1SFw7hVpQDIiE9BpmESxMA
eCUxVf2L3sxfPD8OqM263vvHXxCm8ioCJpLLGdFx1qvlm9p2FMhGTMLQ07elp0JBthAT+6zY19rV
SpV+4nH7k4ewYYZP/qecX+qTI6HVy69s2yMW2/sy8WATH6efpxfedR6hqTfYxZjxkpdGBxAHknFz
OoVL2Q4Kbgd+qefzWTXGs/lZqsjhjw8oH277oTYuf3D/tg7d778VKc+QswBC8CMUCICuESBNK66/
5/BKkshkOTbWmvyEU9DWNXOA9fW6732l8dLLBnz0WNQfY/2JS1OBZGuEs2RelCqkXMd1E4Xvac9w
ITcxFUUcgiEJlYgICGdLZBuyk6VYA36NioerJGrMNnh00nnWMH5xTZq27kjjTIAX4SxKenMcWGal
W0CRyLsLpW0etPGA2tvtMDNOfWUBPPEimE1CX5Sw7pDDDBNTWFVvMorgqBbbXfO+/5cX5+XAppE+
irneMripCzl317QoO6SxrptszPus3I+0EBjunaXTvcMyRvVeQ726PbxHOjm4oUvJ968Unv2YDa55
RhYRP/NQY/+u1QDoeqK3dbONkSF+KXqtJtwzraq/4lmxRLX2ddVFkITBA/xt1VcxUyMTTQ9CNc90
G4eoHTq5JM3XqkHcI41UpCMJGEntGwC4HGmNFdhNHu7EXMbIeLEbHDcavqr5og6L4pQgqI4yAETu
mvSLrbSV4o7PMmvU/Oj/Le1LUfreJkUatbvuWAGipATiOht0FX5n4rtvgGLLcOxTsNdmbXSBKVoy
axKAA8/dImVqqd2I4acgG2dOiPbHwxVI0dX3lm4YflJPEY9qgi1fQbyLiqxnFrp0DFhJPkOIuuXd
fDUpWZCb9gYAFg+Jv5kPgUCFGVMCGSAjA1PFBjr7MqGyqMzSXwwNysnOV8YIRbZ39PZSziyytIC/
mTQl1fxOGkVK10YWYNK6Ryt5SFzhZ3MemszBB+U1+CGbCaU0ktRO96nIiDZcAm49Upk2RbIx23bD
Vfrp232X8+9TxjMztUFucCHpcTXgob+ErkH2yU86yNHXBDlIYsaQ4Tea6s5AHP4oklE01fxaglLC
dWH2ZBsbVgYVqYB12hLUiXsn5TjyTSmujJcR9S+7Fmqr7Y3Ebae841uhTGGDz0KGiU3hTLc3WiK9
2T1qbEkfLcq8hPFevD3b5m5qJAE7+5v+XtHrcfiPl5SuXLXv9RFyTOdu6T2rlEH8pcQLb7IcPU7x
VZZp22ZQWG5O2u7eaOuSfBEqMi/0PGA3M6oDrvdqo+TYd/qIlRiyc/IUy29tf/rrEzzRELgX+i7O
Z4SF97RjTfy7+Rnl1rV3s6dLc9gApOwK15nZWkjxg+9Z0r5LvLA8cwVnBMynntEBOc6OIFC21LWJ
a6St9006azFGVbZR33VZR1MtA5eBfsVswUOqJsyee/Y54ugpLd8aERGxcJMJbnWkRePzRMJeZwC0
MbQdxpBdtH79v7I/SUbuo6EeSmVnhtwGdBqBZH0jvxiTZXV6HJYIsoOITsp55UfdwveL+vp8cDJl
E3EKhZTMM0GaAzz+omjBYXHGEDm4pnk97lxlt2M469i2ZZOO7scB2oGHaaTLRNwyaSM5jA2KBwWJ
IGPmhJmAsCSjd+puesXOBNymkcwDvNV4kNzVM568EbOA9Q0nnuTY4jbirDI3yLBt0vzh7enzkCPO
7O/JSPRgfshTc9Y+UnWihmdz5XMKkPWsCTo7tjNBiBfUGOhDLNhCxX362FVqfsyK0evUsT4WVEKC
4fobi/XZj3GEZdpZgKRtL/iK+bD1Cqg4NKVVVaJ9yfRVBGGpOlwUqU64Nsyi5mgxN2q9EWZNOF/y
529xy1WmbBHFs5M76iryf4t7qwkrfYyW/JAWeN7Xwh3s6da1//Oh5tR5lTvWiH27bjt6aDN3JpmV
oCiN7VNY9EqyUx/JXJcXLwuDz5xNJaGdFfD450HDwFmtzr0IN3f0GIHlQ78e9FYp9ug7M9TPU5Fg
9b2G8y4FOg8ZkbfObHihqVx35+x9CsDRWIK0B2x8K5SmiuzfPHnI86YAySdeRmLo34DRvsWY2PFt
S4FmUQ1L2fOC+LXWUv99jQFGdGtCyADCR6N/Os6JPsZpcOfsblcVSJW9LnjZSZn5sbTAlpm9cbZI
iN0TUX6+88B574fKf+wIBRjL99XlsZaoxXjAVvwZvlVsntk8BC783Hi/D3/tiE1lfbzSdpZm6+4c
pwBNDIuMT/Fe8Vi9i9/9ogm/1psxsSJP4SoWxnD5r2UGXw1DM0FEuYQSM0Buv0hB/DCulhf7olKF
E/QAnLgwDa/sghUV0Ck6GhCpqTuH7hR/FKInFCuZObHV8f0evCgwMglaB/t6ZAaw22GZnS5pJMFd
Pf3FNBvES7XYkQNAS4PafTvnBXOoCUIobpw+smLO6LVOTcb8L8pQgY5Nzfd3ar0aMuxVAhU4Vbrr
YPlJFrj+Z5kfPUk2mgiYqVCYMivDStP/UYVxiGQaGICQT10WGTlxadWZsl3Uc8a3MByJ7RJfrDtc
M+eIOCAfcBtUp8EOUD+U4uoG6QrQ/iS3OVexm8PzOwTpVExoFcTdcaqv+n5U2K1jtehDmN/UUSKi
ox51VZGTC7E7zie2mH5cbNqWG8Fan1jULCMTnhHbEHJbKgeHzQL8RXU3VZ5s+gfX1C3sp2Hwq0Ah
hNPRVutJMCtGkGvJVPC1CaEVZInjn4JS298qOL3hhGTYtnLH7OBCHa4KxoyUzk0qGbkx0IthDnI1
uDTVE6aKE7IAmFk3UEhYnhgU8CQfQdu+YDAz5hsGX7qI2YgNxo0T7CrHg3JM4ootLd9c1/qr0tlm
ckzPMzE1Un3wVtEWVuQTMdLQfK014b/zB5sek0E/lNA3FntYbyl47CkV8vQy+X/UfaNRsZ9m42SX
hCIfUk2P/mZLhPo4rl1Np2V3/4ioSJHjo2N6rb63fgKJEYoVNqyHj8a2ntaeNgixM0ks6g4rZxKZ
D89ytXnBN8DnDkjnnhNR6Em595PoqjNWLG9rXX4Pe+gIUpFOCllOeX1CagO3QZz0aPBf1RMcTlq+
UoPZQ81vyrTL4+AsU/W9UPGnazbLT+nDuj1uL0B2aIvhCViaoWIWY3zTHWcyK/6k1/fZrCjP7WrM
S6j1wjsxUTf/siLjQYqghtoAKe4dgg31EtpqQG7d9AxV1n5Rs0eSXVCo1TprfkJTQRt0n+raJcvX
HCfp8AjbgJ4qpy0C53nA8dLEowmFfJPLcoDuvGJ1/a1uzXWtBNZscZd/AjpYW5XJJEHy65oBJ7LT
R34SnrqG7cgOHvblaCGUDEkG2mgB4LTMYuNtvs75M9UXK0gZMO3VenkUgWjl9OKKMJZiALiI2um7
pt6BkcjTxW8ZSEn+Lf5NjH8yXjH0vNbDjkpLvYSKk1oxKsMmQKMCGMMY2HR1Cj1vX1SLqVb9MOWc
EvahJ+mp97qDjc9iAuRgaHxcvvj4Tn7ApdDoTWgriI6aYpPBj89WrGEeBtIhXFhSujQ4NS3TIBSR
JJiZgat3ykgJxvtUhtZsRDYdA9weJERgwxeYLHaYD97FkNS0SJDIqHxNuqLearheTqyh+K2gPOMI
r0PDFvcxmLR09yLF7+wqH3QugF3vf/CNBkKY9OEVWRu3EqDMhnWZzhP+I+Wj6UGiZWoveQFgBMCO
pPWzS9RxDRDMh/c5KyQaJZ02X1Zlfzzb8UM/ax/rSIucdcwT7lYDPitHQJy40VMmWZOb86lZmpVQ
iEJWLLapwGkvD78YrvpOzwpV2EckeFyqytgQFJ7YmI6btG+tGbXJ/BphR0vEVDx4dwbzZqHqGPk8
kodMIKYlT86S5SXSKtjfSQl/QjvULVekx+E5ZMDbWmWENHBiu17MASNRArSrwGQwHGM4Fr5T5mD7
qERDsKz0u5WbHlFeLZJiSrjk+07Ml6DH4kzD+5QOkvffTEOluZ7Sc4EIDUm4zJEepOx1EK3SiDrk
t8cSAjq5q2YrrycKYuZx8Y2QPkt2uNjKBew9P2VQP63IC2ZylHcAGU5YyEp3ivCYBCC1CuTvt9LA
5RvQCA4W/lGpHGIu3Zm/ixoeVMGMIgQflCzOr+f12lJn9y1HLJuDl6Nws95lpm9ElYy7wouKAKcn
3cP5nFoZsPQXJdvDMbLNGbyHFZZt89/p0Pg50XukHR+V8qwEAoQFJSjSr8om3seGWRBYjyF24mH6
CgwqUTEiV4GWSIw6NrWvU3QLwbluigzfiuEOe9XegsCX9N2vIbelglKyR4HcBAvxep2liWPndgOg
HNBANVHL8XHbyk6xEW+Yx5yKF0U0XivqpsITJtj94deqHbV+vi/p5KlZHCFa4u9NX8s3xwI8hSX6
kK8HKahY5JMFsj0eDqOG5n+HetWoKZNZOdMAbMiSf5NjIz8Ne9xbaBvdhJgZVPBK0LfWucQBYFMn
towQySF2kMtiQKBHUcSr9AFM4F/WQ4Xh/Hj6GTol3pPYjrkzO3EEkGkYjI6WfxmDTr/EQ8yzORsZ
A+94K49oK9/GULwsf1ArOjN6lEUuCgiWMxJeoFMkqcWkP3BOAdx3cgQQBD4jTtrSZc2cRphHt2k3
t4rDkD9zR+Y8bUpLrQI8l/iEY0bVz/vUnTx9PTFMR3GGN6mZH/cO09P1HIv9SVbjDICjZUWacZwr
kp81Kkv0ioGMNT3G4E69XZVrJa+yOWtyEzSKMff1KhvKg8Ma6IGLuUgrp/nfvva43p8tlR2EZGlp
CQyRhdBpaKPL9uBKm0U4tD1EAnqiSbjeGQhDvSEFy6fEkyeAK0Ew6l799iT5ZsdApgi13BxzxWys
XZvg9r3q7S7z6JGr5qLOWEMWURCNQ30t6uwGFiGw+YpMCSqqftLwcPdiu9nzDXAKGrSIzrQN4iUj
2A2g4GbvGTh1VI2sOn3boVv9mSEe563v6NryssQZSv0sFna6JRjCZUZlxMU7QOCMRKqW2XuHOVHA
uZCCBJJVTWSrM6rHgdJDpQMzeUOueuitYfwamN0hkactgGZX3Tn41QeN/RoVPy3eUVWcCTxGqeY1
ol10YF3vu5YCEGWwszpuKd8f6oXMfBrFjbKhdShVTFIZyl1Dsq5OhkbWumvC35JcYkCC4fNW2XrX
bqOfxUbfBWEN29SierN/7YpDTgwQnAqesKM6P3GXdWmL+hYRm5MYwdvStvQmJ8IdR2v4VXiCAnz6
eSGoX7tdy/MiGLQ2Z5Agrl4dtwsb+TXLBoeOvASU76kc+lbRu+NWAoWqMNbw65lvO7OH+Vy5Zm5x
JsMNnK8kr+G0gNrbuGPJKKrJqhIKRQbGYCnknjG1h6Dw26bMbf0RReokwRDOXfuzePbPIs9Mhq3K
ybzEhsVbNKqQ/Xmx9qoTXBgQSl1ZLgN7NFJcECKyJNezhaGgWXr748q9XAgGigiUbetryP4nLYX7
8g8Olro9Ogzbh4kMSCxI0/4FwLBFY0Qq07bIKLayhTQytuA46bs7/QKn5vqHtCdEPYo9+WUN0qqT
1Zl0QaT8xXnGgCft2Z84GswYqSR6BdF8X2QGa+Iy6SEExY4IZu+ZpAMEtAuhlmZIGcqxdvJrWvR9
cc7RY0n8CsEeYzrj3htIc+mVQRBBETRwLD1WYfeOSjOory3mp4MC5LmwewUiSfocwma74eX01lsd
7BILOn222upEzNLdGJ34qgGnTGVv7iK3UY9I93FcWTGAfWaH2xictCCovOjdMxdQmKMxfAwBiZFU
pn4Gs4Ouky8C1ngS0PeJPC7gBs00fRS32FEc+A+pXW2hXtRik5PwFNeXdQTHXbkQODivDnBi1qRi
nzfKZIkoTVIRptHt2QmvS9pkOCJOFd+wYlFlnITzsF4jp58weZWvgytivsJFo53Zdt+oXCSk3jpo
4AxML/B7gcmmnsoulk5UKejYGk6UrdT2yWyhFf9D8azsDpWMan1mbe04ebXsGbBRZXJBw6Ji4y0a
AeqBfrpdjBSHW1v/oihq8Q4VEQQAK5IqVCjVwqdP7PJEv7fEetknoF/tuVdZGdf/XYTEPRRbgKt0
LlDXD8QuL5AnCUVIdVcuYT3WXWuoEHa9pl8QJbGrUpS0q+BIHB33aQ1FklN6I02mr1boT4cs4c61
fvcvLNSJyrkzeuDujCsTNrN3BnDzHMl7rsNurrL/O3wvnLUVJuFWdcpqF6sDUutx9GMTwlBnfxww
IwQydDXplYRr6OBJI4DaUB3s1fDSHkPdgwI4LtkK4877cmB1D9KUJaKmDtYIfO9EBA18CU95z1Il
MnqGKdHRxMv+QjSKiJx96n6rjO4CUEk/YTugFEkvSFkPLI1RJ/usOwwfX5Xra9GOQpeBRD7Z/LDJ
e8bInaDMONCpXh+cT3Kcuj3XiXRfqwe1v5h2/qFCi1shLqDgBnyDqkMb97NDMHHWWGoEyt9DtwFg
W5fDAApdFKiowZ238YXTZ6Kp6OIB8EMf7OlCwHe3565FyWK6w4wEL3yPaZS+oWZv/yM/a3QVH/Qj
INza0/V8i+hUGX2EMaiKMFcWQCzxlAkiZ4DH+3olfDCPYBbOTHVFN4UIY7Xh8yPgtsoYUzzj6UEH
iGTEv9s5/KmchTcYrRguYN7+ikHqRiaWx9OV+iFpFN/24nO1F7oVLFr2qnfQbHfgQfFKHdmY6HHK
pOFZ9/EUjPtKbRXCzaROlEF7BrhRxwrHqoumej1cgY824AYSF/ui64rfq7WPhE9iI0pVm4RXZaF2
pwz1nJwpgFZ9tOlG6pAP9ytm1o5Dw11Rce5jhRXnmpvMpsVarkIQGkHXpilcbJ4WP1HSp5iFWYQK
k0SwpxDX594Mj8N1M4XMYLAkqTw6ErrwPHkrbfbC4qJ0oknJxAGvayu+3BbUrnqr2WeCtgKF40KP
E+q3po7/fu96YBJ4AXmTrVMXrTv9bT5vnRMR6HWmWACzBjfXSnHwfmWKIpF4b9S0hZ8sybHmsljS
fnKpFhPYuAzbYHfc+sX94SxIto0ly4jKbpvpAHBQq2u3NahTZMXwD5aLauV90zrd5GAff2g0y8JW
V0lViXya+Ip+dUXRLX8FUEdPzTFxCyDrH0hT9BIwB6gzkKqQX+oITLqQJAGvjUb35WTOt3uKU5Rw
fPl/n0IUJPRcPVBEtxc+PvA+a3b7L4zfIez07whN2ukT52SZYAJyns+oioYQkFpdffTS2Hyg1dxw
tBrzSsJ+FH6NTFZOXU6QQ1grLybNGcNVwERqw6+vp+ELwDx+CW4Z/6TYCk95zMgSeZoLlIiYnOzM
Q3r++Pq51gYtVo2DB25Dsc+4F+5rzLjHCwWUk6mSMD1jP0yp9yYIjUN2DaeEtv72kh1q5Xlj6qWu
DM6CoJGES9j8k+br+pI1sktH8eFAPL2K6mXaJyNB5RFZB+PBgcnZSYoEH7akbmPSoHiTuDMoJQrP
aeB2gvZBvfN/XJgl61xIWcp0MIqcKPgVCNBBVFn42p8VMhUH5E6Rx07dfV786IMcBoc21NW3/uVj
EJGHz5JVnnthuC+oSNo1SPKhAVg+nNy5hebfgqlgFVADkP97DGF1/G5Ov8buTk9s9C9oHl0ISdCK
WPV2Io7nbbRbCbdUocBMzTGci09WTlwZeRsYBhLv+XdU+7NIAdSqprnV69EeZ+yJp3E7pvXydqyy
dx9uRk5NNkyiGUjRYI6GVrrDngBNq3L3ua8ElXU76Ux91fW2Qn7D1CgmfOIaYnfPtzPFIzniZWKl
gDEy3NBXsdKaOZot/dA8jJyMIcXJVS/XBvQVIz7eFm6B42nz210ew8ZjrkPI/zKlBd8WNsPrXOEX
2p+rU4rCWlrtL8OVKjlaiMgMs0zvsAGv0jNbMjo1ZAdHTN2y9lwY/h2yFoRiLJseKFsAnFl5JOho
TevWvIvl6kCKWNC79coruZXrVa/1yXxjkEmhXQoRXon2H7NIysEsY4CCGUKW0faPYrYqFnsbzuN2
4+1HCCQETjcEsja/tfOi/xXmVICkukysXspLz6u/25urhU2E4o99+97oqRwWil9y02AS0k7nF4Pu
9gWJHmicfEYrk52oreXJR+MRxsDaDZszrpj4cQGDK4xvbcEXrkYA5lndD+MXKjc75GLInKrz38i7
hGBowD8k+fcWtuYTnLQw9vDiNl09lXZ1hUzIw2MF16AzTw8towuzjb2L/mwH4yD7c960LZ5BbLqF
kIyNuLEY4oWevMOdxUkiZZ5DWXXypikdpI+rviRKWuOSJC9iWY7N0YBBhUUxmtBUDwiWwkGjeXSs
4t15Rr9/f7W6QWAuXjBDXlDOf9Rdd7lzkIQ7XR9VIwi8XRX3Fe5PN4/apMrl4n9Kc9UzuSizaak/
VT0WGHjscdGLgf6PBkpLLe9wMz/10rbdgR7/KRjxIUav7sEjXrqUEMrzAj0avHPX/w7O/nHlLPLe
vlJP8AICKeUz3J/dSENHMNv0uTDevXQgi4gKgtFOVVJ+yG2KVXwpfa4/0DwlfAbFYNRhhGRYLk1F
WAY91egJrfX0vOpnE+nRUJnNlOrmyAFJ9xU/SubimbfxA4tPbqXhWfIol7HWOC93xYfyL/FO2A4X
5copXV63ZjYIgpcGPrSJJrACIyG5C/HoUtDAggwfG19Fs3rpo4oB5Z5HhYwsCm/XgbwYrhKfve3A
utxgi3qtXpt8Kl4eg0vSA7MlFci2l97GGraji2Jbk8tm/mETtE463zfnSaPYdOoE9oI8RDk4YZut
zb2rz509QT3yKjzkXO6yZNZX77lgSslk7bepqlx6dFyBUrPYTMn7VIcZXt/7WFk7LoLuI1NJkJhR
gu1ySKWpt6xRH78dgsWptdOUT3iaFD5CN0HSUg7t8+J917w7WmQ6W/zjWNh88a/87RMkQ4QBsY2K
PRGfrfg/g5vnXQQ01yRtd0UecHUaWWAZz2BLFx0DMlO2ujyQN5Qoky6Fy/m/kS/j2IWFa0YVPI4q
sG5bMBuB4vKFSptoCba2oD54jz78cYil0wEpqc1bFtIS3FQRozWuM4f8lGE+mKwUO2fiuPOTDQRP
GIFG/jUei/UY7otNiXjQCMqlFLy1XHwUhmBku/K8ZjxPbI+ozeNvicCmHiMfGtecFgcMUz3ZsTj4
IXR60Kl8gR1ZgHeH92aNrAtKm5LOMZW9M56qAyn+tNh+UJA6SBw2nvVmv/aUiP7/7JVmZQFEIId3
QY1xMQ+vnsxOhtzKHWPE5fS+pTmrkLf69n0vWPtp5CX1iq8YAIyNSNJnzUjr6krIuvMR2Haz9Bji
T+cS0HKbj/u2OGD7GaCghsb7w/L3DwjkeJlzfV+GSRTwBjHHcX/GDkUtOu9fLbzu2zcl1mHkCqX/
qlIU1YUAuzEOqflSganU9qt1OU3KhAJZVs0aJd/mNqkDU7PN/oHfkQNmVrnwcZxxLd3jp+7oWUZ5
5IilTpvg0PC5AruifVKv4EyY2sw7ltTlZ6wPb/vzNHi2ph8QpZiHxvMdyjLl8lNv78PagKIVi6zr
2KVLF8iQRSkofgRMskIbcTj3Ao4OKOxS8Pr70M/9y/PnxBBR+ZvuI60lRbAs8mUcLaZvJC9P7xOx
bWiUeaKv6Pe5Ae2+6JrO6peqRdolIbndzwN3PvUU4WVpybDfXBw03YwDWOtev4Ymg5dce2xsKgGc
SpjAXE9qtWIo0vLOVsyuYll+IlBu9SoJVxWFmp/ZUaaB/1A6C8mAmNxU4TfoHX4p/5yHB/a7MzrP
BqJbz7oAyZu0FmEQUfe/KDN0P1bekSqN6gbS5q6rUb+lJ05AnySZSR5bBLMpgRtYVXXgSEBGx6Ig
5k6vP4oaYU+tYE0jL2F2517FPJ9TiFNk6xK6LjFoBwLO9WmKHNrsubuyUiqsIm5Ls1PAQhSe4dA2
Q0WgxAz8GiEYXfb6TqLQDSA/cJx6mb3DqzNdEsrBzaO8JN2wQwNidLIqHSLR7u3GUQNE9Tuenslx
RPNZ7dVsIo/JJ15d7Y8pG4tSDjCb/4otIz1briTdZjW3UcYaAiJGNMIM29GC6pqwIYAtMfozPyYG
Ks1jNK9tBErRiE5ahFCGObcboxmbQFXH2cPUKite7okUFvhJiXe8s/ek4D2SMUgY+x7D/5H4DMC9
hA2Q6DoS8/GxfC7+6hG49Cl7KpNIwwqyr9aV2I18qSpDSpIQV0wRRocW7STET5mzfVgjZ+rT+WLL
HWO6mDPVoYF3xtkszONylkz0g+4L0QrMCjxXeis9nhLXt0S28QCLohdq3VVBve2EjuY782QXbiq6
HS1W7MDVqNHgSm7tZaNyRhaTE6rg6AM2PUA4wQms8wMf5wSR77VTrATJQU/Inw8HkLRq253KK9Uy
+yxVd0uU9Cnfv9E4k6xAI+XHziS7iAE2Vp1Lbr5dU09EJ+t5RIIrCsLg3ioeBl9fJlaPPhwIIsz0
oSJVJmfqdxK0XkscrU+5SuLjUR+bpMjsPDOk5vKP7WoMmA/5N9tOxp8me7TUKBEt3K5NfBcYo4WJ
BHy+Tk7jPPYc000auoOn2NmqeSS1wlLUZSZZxT7gCO38Ixys7lTN4e3/LInIQJWyMiew04Jzb14r
vOJsPceYIWnurvc2D9kE1K5jv99SAIiiBvnCz+Somh3dA+8EGbmxmhwX5Pe7f+4UPDS3Kwvw5qN8
EroASW9EdJEKvTFZ/WO5nVAp6jsUvZzH9pawi6qrhw7Y5YlPRLVl9cQa0vc/pNIK+Gys51yptXRT
WmBNaKSM68XUyzXejGT8kQ/DTGe2hpuyan2i0O/wrXRzqi/v0el9AmC2REWrE1cmYbQlpgQfTz5c
b5dG9ZfY19NdTEcRlKqQ4vBMR+iwCxVNQcEarz1lorVJDaCcSbb1vXHy+CrbcRTjFbJb84FTsBsp
3Z6RHy6r4lAFM12l7/Yq9Tz5nIqzS7Okna8Wcg6uN3y7rQ/ZjJCEdGlKdzlE8e8CW3Vv0SY7MDP+
q8cYIY9jLBc/tydoMJklpQnUCWCS2kTV9bKESLrVfS1/Ti1x6T9Mmu9XzNWfGPzVsTGPlF/l2E/9
7FrCuplM2GsMudzwajFzvKdyo62axF0tumBJDCDTs+0vldkLC4jnNDhguuRdYxRSjBdUQ4iono9j
qr6qRcch4ILbeUHaFX0NjWb/+8EueS0kDZnnm3PFDlh1E7QrE3IAP48L+vdnFz8VKUiQYRLFw0rd
MtmOlvnPfP7birYMoU1oUTNIUnUI/z0MBrJi/s8Kq2dcm5IupHi0tuVDDDz5Rlay5TvqpWjXd/kp
1T6NfOhkMFXivhwxv2qpz6lLyYYg3vM8x2AjJNdhR/UqUo0pfVggYA6b3L2uhCAmmQj8Occu4UU0
zCAdOYIGtFkY3SEcPSjBRtQ8fZ8xcSP4zBc75XuEEd+uFxrsMEJHKneDgUpIcAw8Hwffb1SNOjLB
3mVepWiu5UVQVwZ304+XxdJdNnFzWWFmFSph6A+WTKOhdTpR7a37Y/EEvS+AaCx64JkwesY6/i4L
UKRi1ZCr0m6Mp0LvTh5G3scXOQRvsqpJLUwfUqu0ZjPJY6GtsiKcViVMbg/cvY/nppFqNitrlhat
AxLAmqSlyMNu68FXDErd17p8G8z2SG4xCf75soEYb8kMjTYZrQ9SMioK99dN9U+mEj3V/UvQ9kU/
RFu3S5rUFU3Qq6MgtptbEqB+uOnzkWBLL0g+G0aUQ0ZehymVUyzUHiTuXIH5nxEsxqdEbkeKp+Is
WehBvfLauW1QomdVIDSLglklDVbPaicYYZhIWD/PGGDFfUJW60BIjN5XeVbeh0Z4W5T/XCj6ATO6
J1NMYkZJyJCZnsB/+anS/pg1RGTbjrU7H6Irn8b0/OlYZLPp0q6XafkAQK42FvoHF0dkHr5k2L5U
aSIEqwlrY1Chmc7LOZXa0b+YtIZsgP4lNldnuqKNJuiYDHxENbiT+Xg/LyUNbGmabfe6d5Eqt5gJ
t1Nt2HzMW31oRTnMJsBGpPt9UWmeMpCJblQkq7eQBC5X95UPotRnjt0r4O4V3xRlirn4yYtxt/9e
vyaot8ZQDic90gEbIethWvr3r7ieeLU4/U61NVUn883/jWRUD90DhsLnntzKAtzAQqCwtRrLVKgO
t+EfsM+j+AjnIfEdX3TiNTqF6NYesh6aEFnrI1hFO0COZiTYvRaWB75dWFgXQYXBxnK6hfxUvwWZ
J8GGuJcxMHdz3yvC0nQs77odRTW57UtJGdt+qg8+uTELfjj7LwL6kaF8Ky/zWIHcQmHdpnPL3Xzw
tSaCZgDM76cKH0cyef/lxA7X0SVlUFvMDD7avOltdEMX9i3p5GXu9NS1pbFLvLJgsAk9xz+R92IT
p2UQBRVtmw/1G89V/elN2CP4TWsPBl10Iqo2xopNrlCWw4mZ6HFvW3M+pAHfA7/SW0YtNE8P6+wm
5v+di+kE5id9lm4tAmT2oGwTsyOwdTe4ez1RcVQ1ICf3o/dXA8Kpx3kONmG788Gws7uB5yZdIXD3
YnWduvCnYUHD9T5KbB44IoX99uYzCqyQ3a8TqaUP+lvhiFmuKxjX+pdgQVnlMXEZHVWzBUedkfsj
KjKGgzLJ9rLJVoPP0B1yf+/c7wrU1AJkKxCis3grtKwbVs18jyJXVtNEOncfT7+BXixetSFB/Bnf
E+JTCVpPisfThj5gMdVme7UexCmtwcZGGNGsK9ORDjZ9YWlamhZbGib/9f1wJ7CiRNpvvummrc4W
9G4VWG3SJBfTWq5jE/Jf+tQoKYV+XScg8MHlD7cHH+jx6zrSVxtRIBNmrXFTIpslpIw+TNAFlE4j
XCL0AJ5PLgAGmE0LmpMfx/bQq/xDEeRsbBzHl6rGGgc40oX9TWeP5MCaru3DjBYZ0Zjc/NNnA17i
o+xoVZot2p4wumsM8F0fHvNsRjH4cBqSn3lrAmjMfuyqlNfVT9v76G/1cs4VSM3UhoaCl/5usIGW
AFNG4i9j8Z5v6YSpoh0+GQCciZAN61UGAN3b0+eXxm0lN29lc0ifaQ9efkde1CY/VVPjw5FAHHrz
prHLRtJrCBwL52GJvHC4av2/Vctwzk66zWrkOBAFleVuf6u4kT1NU6E0Yso1BzSIW5PSMbjtJrxX
AsNXx4hdQqrEBTVlR2Pn3klInNr22OjrDjf0lAYGWeRUg23TsskacuVeUSWlXglB5UUJm3rFxYCc
0EqGz/lnyt1acNFRp+gMlElj5/aHeTZ4407JtslVhzvMMJERSJsWX4CILH7pOhwPg+taNgL6UTYE
arsFqAL7shmIWZZqDeVzrAxV5YwUnV2EtFdGTIpVr3RbNb8u/C5Y1gZca97QwHpZwgaaTnos4cOf
EWlJcyvtrJUNrPHFtjYJmwZZk39kMfi6RF6VYo3mmpURR3ywCgJta3y9GRUMpnmjm1OQ7C0SrrMI
wq1tR/bhXdaYct9nMVrCX9YkLmIH6e3GtxXLZeGETzGhL/tGybO6oB0qauXjxTW9rUiUdLOsGjam
d7vImIQZDtWJYQGSVKggFN3xPDUo5ZrW1eZoWTzEW8cA1OYj7rsKTjZd/iSdXDs1D2pugV9Tj609
1oOuKqJfw2rIjTxoW77MQ+/8IoFB/g3SZVT9XGZp2HyUpqa3OEaUfE8kdcp/HqvnmGrv5KXz/URe
q86zPVGGqyyibpdGBkpAW/cU0NFJI8S/7gsn0RfvvzQaC+FzTFnBKOeVtC+0qv/fT+2OMOGU1pQN
cCez4H1McSY+PZlupJHTiLQ1Bycljt/QC7q3RMG+EgTG7h9SMp4GP/m8FZCDJa4mhsPzwWPsc+Rt
OdnVRisX+CSKBSsokYAVbYK7PKD+L+iokO1iFNCpmhGfXf3VMOI3fqRlA+BHZd8blt9GriNqdf1C
aOCT8/PEMCZnw/zyIHrpEEvP/gxRp1DqRI2g75BWwXvOjB3qTMdYB3HAYTHjmJEwQ0R2yCt2AAA/
GPkjX5nYs72llKoiR7rrw2mABDjcT2w+QtYOwVg/5RE70K1PD60fj67HEcgsF/05yGacfJyfRC0O
qmVRu3mgyPuTGh2oWisD894N5HS758jlsGsolQ+okd4HNDzYBb09aGMRsOm4gbQRpAOjJVUeEVTF
q8SGOy2lq/x2UkHXKpams3HW0fD0Lska22KiAF9/UqQCi0qy7zj7je32vERHaWnRKbpqvCPzS/ya
lhXSMbjmGKdQHCyXsPABnWxCxvoSGJIEB9ToCUUjD8OtVgLgpe/nct6bZImgA7KXoLvLKpQSmjh3
pa0YjXRZI6ATjbNTuFNtbGPmOiIXTPn/nsdkqNkSAfptEaw2hkf0nsnPcMFyFrlJqUuVd7T6QI9a
9PJqw3xQEMhLWBEZewJb2vJNv1ThJY4nOf0m3w38MbK6I0w82oKQEqfoueX+3ObKGZSJ2tdxLfX/
mUeNq27kdWI47f7uyAGfhNTO/a/d6D5rNLnDgs5Yta2wMHlGzKoAXZbBK/nKZvTNRNXTvylX1w3W
x3xm1o3g7BAogzjttsxslYY8ZWyyJgYsaorAsBkYq+YPWI9yhy62RUfdLoEr1VUpW/hkuz83y2sW
CucVuWmzu/EucScrZzLEuqyZ8HrLBP6Kp+rnDPR1fPk15ZCqnZc5MCglROCl5FBtJYeKjmjxE3Bi
rLUunsdPGJSxI8SHqpvtgg34nqJZtRnc0J7m8VT9KSAXt1Yc/Ao6lh6T82dWYaYQz9qH/QjHFG+H
Bm9KOC6Oovu7qSP53kPa4x8LTPXGfODNX0jOyBzolGG709vaNedBaJg5SsCjflL0WH0WlbxpskKe
Cd9/6ELnsmlcB1zYg2i9LNK/l/Babfu7O/8MS0QswiH8hZXfcfsmSyMXMSYtvmLxlyjIeU965ZiM
Dd8HXjNjm5OwQTKEJBBbwkEUrEf0M9hZf6MalcMSuDQDRarVoGCDTfH5EkF+sPOQCkj+KIcvncbs
pJtyvNDcWamtcAq1f3Fyhx4SYqQ0+nMGs5bBriD4JFPoX4c8BV0sExDfLCVOt6AfaKKXmjb08LLj
e1cSTnIdAWxdhfYnCvver+7RcIO3uBRB+z2r5o8lCJ1GxqWw9myVmbFa+RSmZB1Wj2UKTP013KD/
0kZsfni3bIIW/3o1XCtjWNbXlO+OnLs90dNU/RqB8X3amKkxpskG6pkoLOjFrneO75cVNyfigPxc
odXo8TJ0em+RNsEJ5e4Y/TyjenX3fiML251OmrMFp+r/7SoH4DLDWltyKac/16hsrXDWkJFnLRYE
Es/VV9QVueMunzMgAZbhRGYNKb8MwHbzFZ0nmDeEZSFZUAql2QeTFhUBbUY2JyNzhS5CQReezWqn
nT75xxycm44u2gHxr2jQFlwcu6XP63NW4UDo8NXzPw4Pifs3CNP2bwWsUds41CbfCUCNqVkoTgNR
PTcgbblV2rgQOdT8U6/pHsw3fgJAwGD+O1wbfMtgpFEU0G1hlQsQTXb3cvgwAP87R+zHMpW9+Yaq
AyhdjltNZuNcDAHVXJAAHRETfe2hdr0sRIZ43zvipk2wAauo+5M9YHL5vAQIo5dJEqWB0hieUEp6
796b//u2P3CWqHNpxGhNNqRO3m2tkaX1OllhE1psDyRY+reAkxE52mUGojwc3efF0BZokpdheqrm
qA9HdT0gvg0j06ZvUlVo9T/HuRz6NQH4mSQloLvBNfgEBkfzGk0JVsZ7sjTQCqNN6/5QWeGudEIe
DQCzBRQa17Zzuu3vJMcMCLnfiX/QaPW814a4N3jX/O9TEB90CyQ5w1M2D54Yp8F7AS/YWRauzsEi
IOCTwJbIIuDuPeFQl0Pm8vNPLdyukb3hIMuOu1edGxaMyYFayzakItanQVm2WYly4FharT43Bd4k
tiK0BBcOGU60Uc9RXotCLKBJ6XmIRjzqJP2DaQFDN/nyleEwJKNuzQDTAJSRhAtWCJD/19Botj8R
Yv3I1lN21BW1lAu64rCyOEaLJ9zuHMwpX/dAPfrxmDrlN0sW1fhgr5rE3Gzj9qs0Z6t2IwDTLq0u
32QMzp3JamhHS+bFBZg3/3PZyXd53IBcGMFrP/JEmWSAS3n3EFsCcAg4o6pMAKs+iD/e+cgeOevq
VlrdOPmhtAJpxTPjVRKqqJuXloKCWLaNIQteslhwoVPcj+ZVha8a315gwI7fYF+87QShU9eFeruX
CWEYEKaGx5chYzlFSgDx6I0T08MaETGWgoZxmIJ0ZlP+TJcyR5Dk0BejkAfiGPuul1Isxf2SsVyl
8uasN85tkRq++QZmjVjCBXrNfvCaAqzRlafmNjYecXQejVTVR09Gj6YwbFIIFbxr7DDXFbO6Xhlx
ieT/U3zF/eM2bSCKZq1oVcHbuxX71JwwEwJvIBQzaD5adI6sNMw/wSPWZvW1yad5kew8WBzKuyUU
sZZGwVX/t/QylI3Jdi8TSUMS2T1Zii1tsVZbfBHhrcCtAv2EulXSZL1Lryy2pX7MD1RkcPyBt7HG
lzeY2CQl9KyTqvcAUqncIqL6CIb7lWSaF+Q451jy7IdCfseA1fq38yW8C8DK1ganflwwV5zxqv8P
7+CKjXHHVLjwjOyAw/hYM/IcPVOf+rDAFtZHkV9gruH80qhaKQGteVmLl1cGXndSABGPJ82Trqwj
gSoC6qhWIqo+3Ni4cJlMmNoqGRE49dm/JKUtmMrmMR4ZOMdD17/reZK3NTQ5CP9INF9PSH5ML9Uj
nLutu4AiJ0+b/zxgUoO6jNQwzXx3r3IfZlUw8WsCFqdx00dm3eii6fMU1Q+iAUGVCn2cFMImUzDe
ThJq+5gTxXEzAV3ZeZ4qqRImSKqi+xpE3gdYSKtbLJzTqBcVGeCBjqOp5EjIiQ4qic7h3CkUi17C
0kuquGkCY/dc8UIxGR2YADGX5pye16LlOxhewet6ndn5YkZDj/PJgN/2pVWvm9N3ZE5R+OSjDq6/
1xigUaa9miDag7geeZN8j6pBvIvijiZrOi++WPvhSmhZLdmrT0zClI8LaS/j4zawGqqsmhcktKCq
Q5BzBH5x/ZeA0+Y1XqdiSN/ygNe3dM/AdD6sheMm/zysv97v6rQ+gvoI1aD9AUaicp4+JaKHCUAI
J84kZiV1e+/AW/vHk4AnZinlqv+9kLRDPoAbdtVU6XND6twrsFZ90GlHS0CPp4t/R1fUhl0DEO6E
PPLkcgsCMhU1nfJR5gwudN030aPEWO8oALFB/oAB5ybvDtxLc+kp/oZ9UcRWsH4j/Vq4lQvYIEDr
Jr01/YteFRGv8XSaLB1+yvWTdfGZrFb6IPRMSytysBNZ4n7/4jqMhM9R0JRxVDAw3QWrhUFS3wsx
BS+jM5YLx2jVg8kdESOHHPPbw3t2v4iArnnThKPL7UWg876kG+nFHG1kQ2x3h+bPgcGyDV5tikqU
NcP9GpFMOK7pZkZ1QdIEPEv8Jfu0mwhqWMUBfWYwdRyib3aOnN4DGuPEOF2xyOYh8BmGe44Wovj1
VJkwjS/HeZMOQquv9cGEVmNPKVb7n6PZKgPS8Qd0oMfskDSjFZ1S47Q6nBPXxv3pa7gxzhSctzW7
LRdXsXR38avtOTA9l10BYXqGxG5M/SydSHJF52ZoMrGiEWjNeS2SJv3Xs5TSLE/q//sOIItOPxrQ
6XL7VilvHiQ40IZBDoRLTGnsJIzZ6uFNOQf18AnyubJfpmET+PkCe6rFWCFUuxZsrFDAX76HNkC1
I1EbxEjX0ivX6njMg8tswQ2bCjZJR5Rik6aAndSJPj+7FwxnD2fUWso19mMeMuxBp3kqVaCz1Sl9
wZSC6tzCS4GDvRLFtz8N6GQJlAyMdBowV9In/x4Q0Qt8XtRlTkztAISi3PG7GOCPsi2tG1mSj+i4
VlTCOR5XPFONQBHwVC3VjZBR1GM4xFBIuq0u4N6weDXl0A7GGzcyceMvDrCIn95uIo6p/DD4CYF3
J3RP6+Zz6+LWNQTF7wBDfPUUb9a9ZMr7Ipe2qGW7ynWN2MGvxwPatnumVUVuWI0XOrZUHAW20J1s
bZ77A4DOFewERRWkB17ooT3vGkUP8lkCN1kK09m4FpIjaH+7ygICtcpTnNuFdyudA73puvOjfEKZ
/mmuXahHaqdPGqfjplG4tIiQnrzMzdayiu25nbKf+ZV3wUI/cX5CvxiBz2WBkwn/saBfkqSr2BRh
cgur7XH/UCf8rP+upAb997P47gQhSvetPv4aOm2pKcnmIKntGwEj49pDJ+84PklBdGFdq4v5FhKj
l9Uk8HrFgCJaClMezBfWgXSQgS6MCb8mUE3bkIGJsIppC3lKG4MlWhDhtPDKIebVa4XoWPoF6cbz
6roGZKd6METaYy8vgzXi69/amtHBIsaR7KpJKLTU21oRFK9RjoB48ZAMZAutAzOf1U8gKYXmbJ1c
utayP0RZEYuKvIuExDircxJUhyGLLAxVp8uOhyHpkDGPW7xuiVZTlLj1BH4h7hJs9inoqed3lvj5
GS/Fub2pYj43FVqzU0wNdgGE6q4JvwCm52Fyyz3cP15M3sBPHRydNuXnQnnh334JF9CBydf2KNAD
WHdtjQXTuwK9EXy0RTNDS6IQw5xACQoeQfhQ1I+GfpTaK21OEqxWNUXMt/pG6m22N0SOU9omgWmN
FbPwU4uTbHoCYce9ianCWXc1MfBsXBEK1UMItFp6c4cAzdHpFj/CGM3LbK0SpjIsbPLLgaIMgY5M
0f1IGPGwuNIV4nkBwuaTJUaEhAGKynnEnQ8WVP38YL/AwBUIh5oR1kb4iAdJ43fLHSoUw3aMx88x
0P+yFvaXddhqEYxml65pRl6/4hiAcw7kWkHQ5QVdako3bQOulxvdACEU1c/6wOwiedWybjhMvYAH
lR126MiRBuRx4UyRlFNs8xZNxX4rZWrz/mU1nytrDbKuT7THT5ge3AeRDsluZGSR2cT5DF69Yisc
dMtr5hll/In7lhRFIK1es9e9KsR0cGlHcFjnBLD5nEC2LvXJlv9XkseSwfs8xBCiT2TmIQ185Tj8
e2Uvvy2cTu01TRcYxmbo0cHTrTVOTKc7yWpL8r2G9/N62mNFoMXE0JZUBwInghR3X9aE7wfkN0HW
xej32wDZncYsGqyCZwA3Zj5PeBiR4TUYpPt6AnI6/bGHGn+cj8LIetA+mK/4oNNKytVSvxFr/0+Z
/VZURxTEd6y9bJtC1JOAvgmqdZzuDXo2ZkbM1hSlJxqmvaQWNcTgkG1ynGzU4etgdjzDH64o/kwB
sJE2Jj4UgeXmzpobeCX0606AbJAsunIs+wOJkdu6pVr/17ic/7pVWLsImCyegISd6rEBGqX1/6Oh
fhMcau+e3c8qGFE6XSsm5Jh6yOFe346KeUD5HT0x1KDVInLJsbM4hVkmqw/UnKUHifa37UvcPtm4
rgE/Hb1OpM9d+2dJp8iF2zRLHmpucAPlJdKHfl4OLpN8LUmU7D45qk1R66r90u5GfbPuDnFyIK+W
DVxwC7TQrt4how7mfMAmfAq9SuBtXBgLk/XGUy+JydhkOS9jiAxjzP2MGSq7Hu6IbJzXBchoRR15
HuGeHWo4l0t0arnr3U3rzw5uTs6+AfG+gFbnoqVm9Dt9EVKj/yHpuG6VcpK/zMSopsQEweV3nTFN
sfr9R7CfGI4hOSOwLjnsm6HLcbA/+VOOnAzHAyomhYLSOL9A1aPnoH0LfyjNXd7bKqAH5erRspp2
QmfyOPD0w4Xzn470eCqOjYOztti189u4Rz1SUozLuWRCV8VIW+zss0wVXjq8Ok5LgzhnOtjT8vGn
/dSjWCQWRptkEg/cWtgHAABQWE/oEfFlcqxI3kALjuDVoy+t6RSup55eW3AyjRUhnIdEEr5dqPlv
aYv+SDfWwaQ+dduM0NtJxdH1P/50KP3e9jU1j0Ox+6GnDA55TsREY2XvFAsEzK9mU4PoQ0Ftwbs5
/rp5ONp62NddIisGxczGfuVjEdrkN3nFfpF3k07QDZAgegqkj19GZn7iS2WB2nu8SI+348v1BNkm
veP6oUSBq6lTawknSxRZgnr4GK1VIJY6z8l4MygaqKC/IB3obSqp9ogII60XTxuLK7ZNIZwkHrc0
Pas6So4pHeBvfmfgK0sWhe9meV0PmYJ1AYEv9R96CK1fKs+Zgoz9egsYUFXTcADLh2M4i15YbLGS
y4CZxdkN7slpvBXOUjYf22m4v4Lk4P2717JExnIHVorb2fzsxHHE2q6IYxuzPM/zCnJTxo+mtMTM
cgS0uL8jHzdmrk0RrSKaoBdtDPbrRD/8HfGQ12Lb/KINWwMu8c/IKBbV9DhJtMd583G+9r/DVbvO
UZCQhPK/YKC26pQn8rBoIPeZ4Asm6dt+uC5TCwfCVpOD6XJT9q34tF2Cq5RD4KY7TlR7nt/brUoN
VdPEZzvI9eDLAE1QjUhend6LV5UtJ/SWzNIUFzmNr8zM2RSuENWl+GfJbevCy3lRWsI4PSb9Pk4K
taO98f+Erz+nHoDoexiyT8GNhQBIX5SKelglNHybBap1JjomC3U+2Zml51I9Ju/kUzfCi2Eqkquv
vwW4zxsvJs8YVijfdVIsRj3xfupH+2yytPhvaGueZynJshkqyURTBsNTv620KH538Iomw/E9kbkK
Et4nyZXGSBRJ8wf3N/aIBJ69HuqgSQT3nzrnvkSwO6zRZDhfLMNnxbpz3BscbKxL7T4vJ5UjhlI6
iNT0bIuMK780w0CAMwUPT/1l1KPyJYODmeJDPig5LoJCPUUZ+wvSnVct7pqf66es0Oi63QpVfjLI
UARlodZ6yVToq758IhLF6kBkjoz/t5vfh75f5MzvrtMMoDQUodByCb8D5Y/ZvA8eRL+ISc6KK8fk
wM/QhMYxEFFMgwcT57YGg1ZFu++TPOKUqSTKHTFi6mBhyu8ASLK0UMnBQcl3F88OJVVT72v+e0r3
UTXqyxIb0uvTUHHHBa/CVhnwl6NnnacgigrlI+im3UwjRhG8Qad6BT2pjiLxUOFGVQh5zeh26NkN
9ykDEAcAapFUSoNHqg7iDvaVxW2DhBcAEqhwojFkWH1QetErkRSIDg+B1X80q9CZMWx+uPG8mr3i
wIvf1wWwyZZQiuSh/Z7mKjOINtd6El9C59rhz4pFAoe2Bq6tcYFXPiPLsan3nPAhXQGMazRx4Wjd
nOBYBw4q8jLOH/iUXTyrbCnFx4hXY9gJDu+ge3E96YqZtkcE1WeT6JPml6Q1sKhkG3COF7vRSK94
cJLroB4a382OEmyr5Kcg71VW+g2yNC1ArRandNGhCixHUyU1wKd6qciJ1hpUBCljCactm7Qvoqcz
zADQbZuAvfMDQwLpZAsfxuRuMoNkoza171Y649jreWzOBAphvF+AeZs/QVYGN3WvJcOji8YCAVI6
w+9bsHhoZ810q9Foy/8yezep347xxvGfBbj1ENSXIJ5Y9mq+D3n7C8XgqPmxOa2c78Qi3zgIe6CK
q0jAk54/RBCNGXrcA6mrR93j02jA9CIKgVPrpHmTNjerEL0srmr1oVhSkFaBeqGlk89f0IJ4qt8p
r28eHol6SkrDj6BopGzjjnWR/MXnDVUHlBZotg1SFr4dyV1gXjpshykzdlYfEcIt/c/ErhO0Motr
D4p1vkmxYbOIcghXTqbRNNNz6Ys4bAL8TVwXLWV5Y2vfUkCw1XbLeiQfcPTGydEZ3Ft3DzBn2IJq
85nKSf/ornKaAOLI3Hx8rXP9CeFYlucrmU2a9aBWXpv3NRkktIF1ONjJlNKUubTSwQ2n668mWy6n
ObXpAEdHO6Pkzj23lkLW2wMMaRdhYb3/RZTNzOhWaIAFgDNxlIa04QANLNpaOH+220b+RA5+5byh
HC9Lx6Wu8HJ69bI6GIonNxHIxo/WqHuncZa9kPdqP3bzaFT+aNndU3Rftw0zdJ1TMcefsju9LfLu
hWQcTVrgrTRBMIz28KzCvQPbIG3afuBCC0EJD9sPI5XaN1rHEHw9A5axupU0XSwJKRN2efihJbLd
lKCdjOSoTbf02qXsWYhv13NDDj7gFkEqcN0kIXlRteHOJbeae75XXjzRoZZVG6b/MnHNNj4IXcKk
kR1SsdleJWA8RD8Q/RbO7LCafC0RMg8WMkju3aHt2I4yTweQA9l+wAMHM5prEdgTB0ECLfhrK8Nq
mDtOKL2+223oO7bOXXInVclNVkahJEH/yYnPYGMqTzpZoWG54XowYLXdNvfQ2lx3OqQ7MtNWgV1R
RLtHCCZTe3fb0xwRE4j8dd91nOQstnJDhISMu6FKDBOW1UC7wrn5TY9CjAEvYoyd5e1yXeoSWSNx
n//SeHuQ2MfycGPFK+M9MB0FsEXArznQrkwP8nrA+37jIgF350XEIEv6OBErNwuG15Kp/nP4iETF
QawCXYSTj+xF7bG9A0OWsCdeFdDpQCxHgtE4rU/gf7/mhVilVI8sbBbBGuWoDBlAsMvzbQUyRv9Q
uxnu+lJja/I1IvWcGxOcuWldY7xRwd+3t6/+QYXlMYQN4LU9E2O9JFlikPr9GtnN+xMrF8LRIHCp
/HIfhkHJ/sz+zvC2HmIHTqyY6Yz3OtBssWI0afYsnTit9NGV2s5HjkIAuitAF1/2Sw1+Ic0RbN8w
l2qYWGfW6+K0PWbibbo5Ql6aQM7FswOIwmaSBy26G3UgwF5K0JedqoXXCDSGYmLhjDYyYlq8bGxW
4lDDjsEPILTVXYxf5Yu1uSwrhuVMdRhPZYuMW6QxIhrbWyUqhCOjrqc4DSwuUUETDWwOwo+WU43p
4lyYFMNfqmAM1NGX2/PFXluZvhkuRiHBBZ4KQvB/d2KcxnwWpeuJe7tR2q5GW1R5UPwxEAFxqJHd
tgi7KZgH5EtfYtOhWjE9b3Fbck7dIJRPlqSNI7WcVOBL0ApBtpPmPfKrX2AX2ITVThPu4X+V5WaO
S2LtwWDVmsZFLQT91GbNioUMARgEgI+tEsJ0NXdSU4vy3VFL2KtzSTFNqqyaVYpmqwpkiOver0Ky
u3dahb9Uy7v2Q8VYSS6eOJ5oeyWlqFjMIwkYftClmuuDr442NQxWR7Dy4HcSi0c2B+eNdkMoQQQD
NoA1zESD6vTl3XqdLlzAdH9itUTTV34yoqxyZI87u3vE4dJNbynooePMSPThPkyE8a/F9gu6rkNs
7e0ppX390KSfuLrXhy/Swvf0y3eaMHqDZpmr99YTXTdbsiWI8avfgud17/hABlM4JAw290Wn2Ah0
qhsFB+ioVCnMRHC5mmZAkrbk4oWj7y3YZkVHVao+KoUyblF84X+MzDm010KxedVeioUfu3VagJxu
vPHCJmSHFooFHLBB4EeHaTo7cH6WWqvd3bfzohTm11EasFPTy3b85YnNWjwCyKMkd+FdEekNq+Zf
/7RSBj7IqpatkioOhp2U4tXxlFiwanDdgazJw1SvvZN6INUn8ZTI7gn7h6S5et0PUiHCuymhyU3V
/WZEe6TXUTSGKCPmEz8tIOPdqzTqYhRnKxa3BTykd6MGr9+nXJlqnTdw5pAxr6tpTVFPcHtxHWrU
/deyj+SKN4BYn1p+AhteYHZbwyC3jItE49kM9cddxt89+YxirJzYcuRzdvX04YL45t8jVttpEluY
PQqAqG1Kl4yX3HH93THyP1hX4Lh45W4xbiWpYFMAKJoVQ2FbaUArzkbbbWjWg+UJLpSsuHdjdIby
KtLmbrGmpXTHVYUghPdk/a2OcC3OGqvndbgiVGVy+RvCS0KwCQVC8MiHg+exUW0u5xfUgGBhm0rI
O7tgFJWCIMuWySW1qoO54+Ik90rvn7zCl4zOomkTG+OonJxDGO0DwHSckMUiLcCTaVa+eeD9s94y
LJj94UK44zadxLeh3HfSPDloioZaeAM6jpD3r3TLSeE21fn5Y39xUaFb89C2EUXUPqZA83GnOKLF
tGDjc3jtLkckvYYw4a0ITL5Gxn0W1Ry5nOhhmRfsD2IeGLmFD735t4V0DdPlrB21FSac+G5OqAo0
FmMOINlbOzkLLkYCBT+UI6p6ycqpWzSK+nFwVg3ACbLmWwrwSldQghqjBzgWn1fOUeC5JpAGjO1k
LA3l9z0Iz4IFdCoEHVbPmE6RSyZCgrrICSgxt7d/aP/WRXv0UN0pF0lTU7d8QggQkh16vntMtGYq
y1eulFB562e6699vWAtyHqYm0DmDA3kY2hntHHizhq3wkZ6N3eokMPJgq9WF/h0RYvkglZmJa1Z/
YWGxp5tXX9TEYSiV3aogh7ttj4/WuMH0sOvE7Xf273liuzpmYt8pYaHPbpCKRv/r9NxM45/wvU7y
7iebCu0utLP2DwPr3zeMN9wVMHLZ+ZvgCr3sX20lo/imKGCBixPUOcXSLECIOJhF1psDswIbDJg5
aU+Cb6pOUbP/hRnzV7cEXP3PHy4GrOLmaSp8bwXxxc8H7/uYwh/t9r9onl8WGWhvlKuMhdGWm+73
Vvyv56s8aSkAg5hwdAzY3ETZLz+NyVieGmiUsbQjm3uHiFTcyLQ8vMGnqKIPQCibYzEfYpYNPu4+
305md379Q49u9kfElR5cKoRxr7DSuCbSAsAndI+PHuhAN9sAafzY8kXVEoo51CYLPI6k9p18jBXz
4oIxGN5MHyDjqw4UR21yz/+/Xu5AxPcokuwF1oGwVbWU4wKiq8658ar9bjCl2FKgNUWwXl0O9jiy
9q+w0VF0RanwTn+Gta92v7E/nbLWnMQxATyunTO1wAhDqhkR2QCr7Dnz/+3GvYmsRAEpSmieJ3vT
MU1qx2w7wo/HOwNk1Td3r8iaNt9rbEGSbFM6L5yBXFK8BEYRR8rXcpEfLe5wMjFoGQMgtvd23gTM
XI9DroJGTOvYTLDnYbjtDluAj2V1GjEWAJnqiQCOFDGhPWKBelouLqNVPQWerc93eil04/nAFK1z
QMR0CsXKCrzEXc7sMovx3Y/jgXD9zkZX8Z3uNUQWskqAHO/nPkaLUXDAyxXOd8c3IpCpzGEY8Hf1
R/kOgV8dwzoQiVaptRFpPGPuWer+gpwc1jgmuOi86yX8YyAnAFYG1v0GjZkOhu8CoOZIUIXH7bu2
y2pN5gPVZ+5DgQxESDweg1ogh1kgdqd5oy5xXSE1L016diXFy6lef/ojlbDrxhcdmnH+rlv9X12Q
4Aslo5NyvfC11ud8ba88Lbm9lGR4FuFZXQZeCNTjZF8i9U8yfHpOdNFbOc7uvB5ZCEsiuSKXT8yf
i7msyBcBCZNAf8uRYeifCMhzsNJ3skbVQqRxeY6xGSi/mIjGGPbV+lOnibgkMJAaMGrujTihwewV
E/CbilufvL0Gv0ok4pgk6WSVnaPgSzfR7gTcfDrjUJxM+xfISRaa1TE/DTLxkhEsuEQFnmWw/wVx
/v4PIz0TAEGUHxVTSdFpAuM1rbFQp71xrD5HodSoU1yv/ug2vyM6Kw8MUt5B6fAL6UFhAQw2yR7J
Y3d+/7UEXhgQN+EURad/+ztEZUs7JqCXVn5HXD/kDszA2KXMeK9tYNgr+A1/y8LsWP4i98/eNcQ+
28Aih4DpH6cBytaDF5nbNVGDPHuJpIrbYBu5lDBdGdQyA0K3ZgdArztJEhA+RNSAk3QTQ9gWE2Q/
bzwTruLaKxSHezEFw8MVo2YGFTgFgpx9EGpYEjuoqBK1FbgSpsmCjpxUlpWmbYkHrOSacxrlnK+9
O98wgw5jY0ccnxpc1vTbfyfmbQproEgs/9OPOQdTo41Zw0dyzii0wmggkSMzeuEyYgvZjhtoKQjz
TDFDFYDtHmOakTOChxRl5ZNzjcNVnjZrS9B7Qfr1bNVjtx19ZymXB4pD3cW3zTZMinlZZBXW9MUM
diS5mcwO/QSngXheumOHpL23trrUOABgsQcjixZYyZ8pBpYF+vU98aSbIZIpi8ifTMf7qO8zinrR
iZGVNck/4A3TyOu/R6vy6w2xsvGkVPILTDcx9B2HTF4dtnVwLda+hPrR1TrXH4uXYZMddllC81gw
fbIfZkQ+Xjar1KX9VXpMhUPJwYbin2efGjZS4t0RhgojnRzr6KmxX2cvSTJA8CSFsKAXjkJigGTS
y8YHyYXCrJuREULu67ScMkujLbZ0ko261EmfkizYnyx59O5ma+m5LD/4JuwiwLr0xmK8EQO11uie
2A24hKm0NtV4d2W0eU7X2qtLjqkK2W1VIYFHd/XTSl7W6QQHU923GDVYREmQIzhgRG/2ziHDIVqm
QuxsgvhEHbazP5MkP5CsIS0cV9GRdXxD/8xH5J+tZ3yHjhGBqQYVHjJVXfxwvHU9yZklpXYoHyGx
hegpScXVbqHv8l4QOUSrVDsqyBpRwQuYUv9lyTHSjrbxRdpoeW2Y32ckjncXRqGI6WdNBJrYpap8
T2F9w9dKteqz6WvHkWoQqGRNbocK8yq2RjhnkyoZL9lTZV+mB094zrtzMnaapozmJ7W+MVPtIV7U
dAmmraVEdJZdOhI5rSfv3tpgikrZaE4FSFyGrag2jDzrNM5sK9hIrqVV4xBFUVJN+qXDNMjGOiMk
gLDqA05c52szqmcK+QO8l7Tz4KNE/is3f/sC5ed25E05IdZ5SrtjlW4ZFy800w6szbJpVFcx3jWG
ISKZv0Cyn3gOxZs5oxKMrsCUxcv9T6Yo8G763rLjTYyAXkMJGGTijtEXf52OpIxpNMAzb1vxmoPQ
RqCuUeBs/SLqB3h5bqDVQM7U9+sK+ttWOl83IkGk8iKtkYZiUphdK/gSqi5YnifZk60wleVjXd9d
4DD0NZEzmvFEdl3yL79coLLhWV/k6Hbi4FPuvhc0JKuwHiOPob20q/TjbAOCirwcAUdWhz/vUGZD
IXDLzF0/ch+2YF8u3dW/Kb0E2DjqXV1v3xbbKD+L/AnTn/8iCes+JCLab/UyOqyQU4r+h3rzB//r
SqHhxVBWmk849VUE3+TJzCRNyqgGLofPFZsL8YuUC+sCR6NiyyrBFVr0/VOUlO7Zv4bMsQMJFnO7
ZJiyKmNdHZEX2rKWqUEF8YxVSnqkJdAPSYMjoS7peu+HwkCUYq8v7bD6tLPnwMzXg87yZ3bYqp/R
PFTt/WxrIp/y8sHoH54J1sIXvow2a/oulYAE2pyJ/Sjygx93UU+qkGfABXOvjovaSsLFgQrmrqk3
V13F7ByknxDE1c6r5c3ktWAWYfAgE52OS+rHlmKjs0VKFaXiZgcubWAusozBlViGEiL2o5VdWVtb
C86PP8iKzLt/zi47iisYkuElJ3mfhKAznrpVbrG5cG5OLIE4GXTeWeLSrFyvrTllGkxCRuC1QyXf
mOzDaWTDWJ2j42OsLzSHRfyP41qLChtg2BIfgB/tGKr95kY1Owmp+kbX+JDG1//JfV2HKT/wistp
jrz/nj7JK/JdOXLnOSLffN3Ek2ueKymxVqFK1iLjheOPMlpjf6m0cjV0VL+Fh3VvNjbQhwZt3Bi2
yrmAwndWHIcXIS9Km0bFHsgbZDqe9AVZpY6RHuUTEi6xhq/6Co7YXI3B00jCKYRvMZvv7jrJn2yi
1RmjLCcB5HeIGEjhvfpJC2+vd77TXmHUjjfbXopem0JEFFBicRONxXejGj1vB5oMANvBriuN8TmW
JvN+1WlEG7YSPMrQIP/En1Ro0d+y1VbQt7xoV7mlsCPgQDpAILdV960GDXlAqj2ihfEnpkCEWFED
393NwthygZiosLEWiUmntWyATaPcRPTyxxmNLLJ646xbAv77yrturaX4hpkMQaZBDS1w9ZSbUFN3
0gLOFjfE8hvizIZsGCGlvNuQw6GcjF0+xPeoyq9vhQdw1r1xBy8o2aN0r2fgVdrxUEiO4ZQOfZSc
uuk+IINnsUXbV3NNCvtrQkzpTBQp3NzRNh5JFVhMeGM/9fqZsl/XAMhsWU+aYkjRPU0SoJ3LmS3X
LG0ZOZtGHk2o4Cm6k0N04dFJaZu7ed4BSwwAxD6WERPgG1ZkM73KQXb+4iKTOHak6cleyrb/53Op
FKRzk1IEyuHQ0rpjVKzkUF8tgbDPrPj+l3pLtW5IEJdH1n9e2RXJXg9RR6Xtv7BDJsUlj35Xk3gy
Lgsk69ZQ56MuN/WnFvouW3jDddtVGfASCpMEXDHEzLTC4hUnPzUenqjr+M2LzbuBSRKnBRLSukac
IayKdZHGNaUAhIzC+D0/LwsAQroQBYPtP164wl8oiNrr5ev5iLrmTHo7b3BnRPGA5cbvxe/1OGkc
hDbJWow8856TdE6UP4EdSZzMnyx12E98ZcIrFfRkgddY0+gDTPjAuyCx34eOX8MQmxw3QIvTjpyO
VXfcCUAmAyQ8sLk+VeptXMp/i1J9hHzeN4zuglL1CUPpcixb3I5aH6oEp1ychFTHbpx0SgszPBob
UzPvgIpqZCwIl1chNHNFB0ufA8WD+pAPKaLHBnlporX/XgCf6k3iVEEOxZMnQC7rdHRrKj5VDLSI
qnEJ2wc30aZX2xHxN9NCN8wl4drVKiQtz/TX5xcvHRyLNqc2j1wbQbESwn8VdLKzbGVo6hw/cB84
PdsTl3FW9D3u1DWbiCB733FHrYRPUskCn1keBsgazSJvfHGD/Sle2XWeF6wla5oaa6LyPINwzZiT
2FwhYQlvHUItdH55+POjg375EONPcMhSHafdkQL7JbThMpzK7ILS5kVzQaYxvl00HSw4VA1Fkj6E
IJAQhSrzDJKldllLMZQuSXggfjU+m3MwOkNTIw136p9Mt2v/Ijan3oBSLAP/aBKdkLA6g+8278E5
4wRTBGpRmYzYtaOtmUo4UHx1rK4wXmAEf0GhF6NAbVnDeP4Z8mf55kZsanaPUSsn9a6O21T/YuLw
SXuc2Q3CylYaL0+bWUBS3TUfv/S9CVlknslQjnYq2vTsLdyPyXhFF+ZVMqGv1A8My2HmXx7RP9/f
Hd2vLwNAweUq1GnrN7cooQQgvpWksVI7FW1Zpc7CDoytQy7rHnuAFt9CZNUfdZ8G0ULFm+bjKaxP
Ev/+ppueH/rYltn/LVJd+k0W6FD6/UVQZzy8BW5ghIL1H4X1Om38yQszVWeymTLs4yaAaOFRpXja
wR4i5BQt6M7LA0pPDkGuWeyQ6c8KHEBgndoA9Ya6uCyOFK0DkBAtJp1AeCBHUfPq7RtrZFWfqnc1
rakWBDJrHMk1UikXvzH857cvCm9EzfmlPSR8VcgJDukrkhLe/H5BEI64eVEutk+HlNXb1FPnXfyp
JvRJUrNl1mWHXF4nWANm6FyvSIuhIAuHWPh8KBnSN7uRREMHVzAmibscnMEW5YEZF3x0ZMrTbz6D
Yx87aNZkynsZv+CPSmPQbAz/Rh1ewWeovzaqmZETITgZY6+VZrF+8mfd3UheC1cfitIQGtx7I9LE
RBkk8/8s4MdMgIWGLfP6GOcfz1dHuTo5zTU272bLQYk/EzTl8P7ivT8DQn3UjTouFYh9wRWrbI3S
IOpHwf/MYVAFSkW+Apzo2kd/WPpwBjdEkMJVs24ofKNtvxKX/s/xxHYmldy7Lah0saJ/uwEzOoXp
oEAZDlgWEWT1qVovbH780mpZULQbOpCLiIiB+a3C152QORIqyk0mHPjAv85Mp4eyoFKR894c3VAI
89Otdc4ixxS+VsUBfb9TMJRxIonEG4OooA0+J4SpyKqlG7et8UTHVWZTZFqDrl2/kJJRns8jGrwe
b3Tm8+hTs1eKEqdtmVIrB9HBbIqZUoH7LjOf9p2Yo/6/JGyv6nkMUeIa+iUL8BWPWjoUdPB8g4/g
u63s5jw0Cu02XnFn6w77uNgthYTU0phxpIB8dN4StpnNzVYJ7ZSNKoE+pkos1dVBiCnFxZ/YW4zW
xSZGumTp8/jW0Zf9zavL4ukZ+9LzIpPUfjiD6XVKyo/ItVS9U7yuXaQ1pJSa/XfA0o9Hu/Ab/Ogh
0oh6V3lyAcLHN3zGKYEub9ocA3ATP4wY+GBIxU2rtB4A08ymg6MNNK0QmFdZmLvMRNibmTmxmIvw
dVZ0w4QvpGIcnjS4IJndiFHfwH2lpPUWNN4vYBSg0ByLjhpLvIUw4bMynYuL9DLHxkSdRpaJFhfs
Ncoy2PT8jwsoggidwO5PmmPrQYyoYc09QZqvagoRaE2mCPylxCDjOUPVa0/3jiF/1i4dDQcL6zp0
wSa/xUWhG6WSTUp5CGVOyJrhH3C+NbX6+iXi6L2OCpKbY/UwAHTJro37REBIe5epMxsxNjCKzPB9
xyJGQHMlr7W3LinwC9mZHYWFgw9uk1sEvpr3a9YC3+s8ZT3g5m2kiMwfKFConQ0+ZD7VeNkqpBls
58YXO1Q5M8ESiVUT6N9wZXsACgwnMldfBkR0P0PdlwuGWAjlI2GFc48JEVy1NExgyUE0RpNTHU6r
yHTneZeqVVjtt5jl3SUFeR5ZzzNkRTG16OeuehlFA907riFeSuK0uFw6tB0klctG6NbZQozh+7K8
ZyG97B9j+bFcNrzHrc+YU1Vyu7xvEsiwQd0rkqtQ3JKc55Xz6LjEpX4PwGh6b8VzR+MimVuiaXRV
BBkSPlAUBkjHhXbs6vrvVD2u+7C4DKy28oF1SU9Xplkxe+k/fQTTXXyjBh8sPjHVLtC+2RDJDIXx
AsMJgHjStdJidsepruolKjGYkY+Vi65nalqG6snYIwvbufytybHNLSVmz7x8+mBtY3H75+wzTTfQ
Flw9XzeQUVOhQHf5XL8AMzeRTSr19F01FtiWk+H6SPkhF8gsYE3Kgq8m8WLKfutBC0REcNFUODMw
rr6S5SDLGe8z1ibCv2zoIvCZuP9d8pFZD+QQ2EW0fRSDRBox4zKAdg1x6lRAWYmcB+TfN77pvqvs
j9LZFCsju8JHPljOgSGAi1Pdi1rtko+wsInPnf7hy9PjZzOz19DloYNW9atmvHlUOmUX0FcRtaWp
UDPiMeIs9VfnufonfJQibdfsFr9MeBWIQeo9sFTvfrRcpuI9vrhyqg+wlbyC+MTLR8CP+T4EhETs
2phZ6wRR9FY+YeOIWPyl2A2jh2hdVvslbR0KvYtb7i2/cINStSi2Kr8qzwlT5lQoEh+3Bk8CGpFd
7r/jauhmsKi73J4La5eWzZbirfoumBpi2kWyjawJ/14+S104p3kxs7IrDwU9g5UVNQDTjUGo5u/D
8twOF0bZyZ7mE+jN7UGBofLe/5HKTQ6QgimlGHKhe0XIVIxl5SekZrJsefUs5d4bxU5Rktc2GsAE
XeiaUnUDviuVWsQjD6VS8Fa18d6/hINKOc+QQEtpcpu/IrJC9s6bjCdVN/KqbS6xX5SHC4ERTTdt
UlAd9ZcfOLXuPg0JW3KC1onSP2WEy2RSL5chwbHs9t9ceaV1f0vFIsOzulSW9KZiii02DAuSbTkx
XBeDh9GI9tjAk8fLl5Rf5mPljJHmm1hEOQtiynKHwhdI2lSVtNx0sTNaOYI+XItjYfScVDHZOVaq
v6O84QHX3VhW/8LqaMoj8NnDe+XPn+wy6DKbpqUuMZSuSm5zl984+4FQroijEGX4AODRAoop9Neb
uQfKoDfTsDhVKee131GJZMECro1IVl6/F+6JNM4G27MyrY0FRGdidjbSLDG/PasyWQgRJb6a8f8Z
d+TUA0iAnloF6QI3z5FOeKH+rOl19gk6pMawJrW1juRxMZjISxZvI6nvMRvK/bU6UxPhDEs5sYeQ
pmOHDmsJw5vPPw4kKBEYNA7E5UX0y15rRhqO9o5gxXtVAxzzvH/Fzx5pUmDdWmM5FcHSmsADi8V4
HRMhwZwbQcOlZaUrgfcTO352GLVD4LF4+YO1/LU3bPEnT+R1OZDZcAlo49yjRpcVHuzGii1/zsrj
zgZSske08u8QoQJcFXBngVLC48xzAMOEIsNiOOwUVBYDSxtZfkA/TTHLDAgbDnnP5vrJgM8gQcQi
0kdhOrcm0s5Tl1L9hgTk0oqZYSF+MDe+9himCanTAZUI7KbCM1WoXkd5qgQAak36fJa2KAXZIn9+
4BEqm6PhMOsIoch8i9sO6CO9s58D/LRots8RLpLEFYOrp+Dp5sGENw5Gz2BKhLbIUd6iKlRovA5a
6hlNxDEFwXypOqU/tjoK20VLLkOHV167L1iHq6nDiLdohmBxv243MNy9PNIev8GKXYCGFf59cB6D
N3JR63B9saZRH9n8CvSwzpf3AZmCGlD0Ah3uO2vNkCzGyrEO1fokPeWs7X+evEuiWqeCn8qCPRFS
nzwxnMSyzj4ZrkejvmucL9/cqsSmg8LEv2RMxjLnQV8IVqU0oVkGmQssGiH1xr5vgNrmYKLGMRFJ
Uev70GobAZkgo5GR2Ms4wIV7plBpMmy80I5HIN3zOs1NTrw+Hz6yOlZSWDwZn2co5+89uvlBZ1Si
av3kVthv3b+oEuuLGUgXTrH+ZWZlXxCou/QnBxVuMiZQ+ykkNtGOVNzhUnivJUUtPvyiBndoubNc
u/IYu27L+Bp7+JNL6ldnY+xIGe2/brz3iTfMrdaK1YgF1Rlh3Fp1jz3BiGK8VTkBuFth05mMh3EH
rx7SN/KCceBL5sDJyIcPCEbjcTQ8SfcaE6f8ApTKrqsmgXb5BCbab90R2Bz3YoubYwK2rIayU3em
jWxY8vJz2COB6K/yHQQCObww5xW/snyeEhvihe6x/sQojvD0zAaGEt1y28Hstnpg/3Vcw3LN4MF3
XW1ZQ6FCid3+5vYSDvhB1efI6CM9e2aXzV1Tn0C37L19Ksv5klAsrcKpwBOj/VaPxskHl8Ske4Jf
2L7X0fKqdRLtOzbuor+Pf1MUPAqXoL3pnHFm4kQpaBlsq8uC9wOXNDLGnk1PLhR4oyGuwLQxwwJP
HEydPbc7PzkU+lNRBWZzpU5QuXhJteVkiRn2tB4m3MaF6LQEEd9SlG+EeBKJypAJtwMPiPJM3Q9a
8jxXzObkRH5LE/uwL2HYk26LZwZLk3UmkAiDKyAMz/m7HN4pnprpCHPUHlKS+8tuBx3NY07twLhO
7WgJseDO64gJu7zpHPEQZ9F8Vgdb7Zzl9MmZK7T4CaODEkDjlCCk9MTP1foQPOWNYlqz+0Osf8Yj
tk4InHDvkUhSc+XIatWtGpddQeB8hYR2yV5+CTJFuIlx93aNFGIy7TjGJ8QexEJxzLbkmzUzUSgs
r7RcgQoI8Lm1nEbzDAZW4KSxqY2MqsSRzTuHKv1TxKfe0rUa+fD85VpYqu9qSCSL1NsKA4yh7+XH
fHBinHh5jbVcEKbdw78Jh7XW+mT9DwjBJNdS+GA+0i6/4tiJcSidPEgCX75epvwrXpvFag54HOb+
kcms763E5RGq2NurWZoeDr4xmuRDd521onIeRwFd0Qe/JWfhsvlMYG/9ki1DxEwf3tuNEu0ybDHw
cV2Ep0Kf/boBFtStod0wmWCz2k4LdAuV4PdS8WtD6rXaq0jWgR9ycJKLeu7dJh7fVxly3dyuH1C2
uSL3VpQa3wqunpZD2WVoq36rZb06K+l95h3BU0+hyqC/847SXdY/2v0OkdZMfMwMHObIqw8h2nCY
pDAr4+UloWDJe2qMgHxcIrXXbc6eozqgksa0KTNHIKrlotfPaP3xsUMYHdBRHW9tXfC+A+X2IJ6R
xEnFyRGidyUDibz/3g9qyqhJn5ygkRPr7cftlYJqy+kZ1BmbUUR2MH8TEG7UwpBuwfOgA3YMfLAd
bFI1+ImALSAzdesYl/dYOkzi3/kMH+sRVq6zcL9Oy8+4jlCU2YLRl+xWh6ki/OesCeKvzxvAr7Xy
3rKzk9wvoAOBnVKewykyZz1vqOG/FUpZjLD7cl388jimubHZs7qB0EDRjXg3bRK3NFmZxuJT5x3Q
fwn6rHKThyhsEMdvGMSp6L8+ePjm0+/N2nQx5hdLC6Yl2PclbqHGLnqWt1W1gsmntN/ktn+FWF/j
67VU7v2/D6TcqUFtmOhVYQW6cDYPZWgsoY5IBpj0X/kodFq6U9Ah7XPXryD26qWVc6TWzBlBtSe+
+ZNOWf99CVVtSEJBlVra2xiOGe5cBwUbZOi00Mz2+D7g8yYYMIchgFargHMB4bLImep2rAjvkffP
XcIIZAYTyarCB5hWH4SoTjef+sriDQlFJ5GfJTQq7tOX8xpUAr/HjH+w7toZxnt1HktKCvib2a9t
ficUQGIKQqgXTLK8tu3QAVvfJLSdl+bH5tOaUlvZbItTaTiSDb6BSUq1MIUKSAVKB/YXNl6b8DmE
PG8m69p1RHeEE02qzWOfmwBMg5SHXl8NgIDZ6YAlbFUalJeGuGfSGVjik9PwCymWzlLiCGuCeJIG
mWWVNHtYxJLFhN2exA6Da4AHt7EHz+PmJboOai/9OuUy+G8Axt+hX9uO6N/75KkheNQp0+unaWYV
pPnRDKthZyoAebBq/lacCfLwi51am03NMcrMekhHSD4R2UtgKiCOKfneYSmzRzxqDjcWuwoiOpFl
Gf5qD3P8dmddc40zt5Am2ulHJtl+qgxaMqGL5py4XlLsidn1tj3d/qLhno2gbes7ZdXSow20FH6O
VyQfYjW+3YnLhB+tys8sAHtg4Aw+EUDa2sTL+V2y93hMtYIYyjafm1tjNYSNk5IcdcpPhuNY0Q+K
ef7mYutUrRpAWnFlQi3TxgPVmxNFXAazGcPqGpEa+9iiFW8XihUkgPKYCBqYP9OdUemuWWGgvblI
L8QCetUvQhGgLtVoTOFEuj96wMiu3nOOkL+nyB2g7g8U4HG/dkFB64TQv3c2GXuMLxsPC5NdAjS6
P3wBRK3SBDzDzAadrp15jR1sjIKJJwIkVXG4v9HiDhlaXvJtZCrwJdYtx4ea548qIWws0FJE1vNO
tC5NdBTuYYEtSAEVOzFIySmaB1AMwuoB3k7FdgfRoO8LXI/dBHxnXJYpEsACkh/gKDsHQldgDe7o
HIfGWGT5esYjSArEGyOpF4jpWluDwK1DN5KMB9R0/Q5RzKYjjtEEzcwDST+fXaCeKazebW45BqU8
e/scnfsI6zQIG4LTHt7sY1xp5DgRqfSkhw3CoZ9vNnwbXGfP07CIV7aPhvxa7kn1iAUtIvEf7fER
lftMKxaKPqWMph44TOq9IFWI3tlPVEhi0HD9B1cZHzR7UQUZoFMBy/EJMNuuA07ybiEfeZKZfK7i
GJsyRf5CiGM1ACDW8c78+dZuzKpim/uod7ii8k9uDZi721f247obtnOmu8Wj8SxfCTndDB1l1YZc
AKJtMU6/16OgDdl938Bq6kd841G3/Ye3R0HgXWof20pfTNZyLJFUnfSHdo6YvRCg1mYqtwlBwGRs
yaz7DZmWR6P/KShQVBk/G6d/rtNNRuPsRXSEfudUARI4TXbI24L6GQg9XlRJSLiD9hVpxNO10Wsg
0za6fpr1/+qdHd3x6Gn9ZKdfrerIaOEBqO3zLKiYarB5rCMP+gWjxebOpf7wFV4zyjYGy1Xrdayh
bZbYkDBKsHofHWzfM1h83RvW5CKUNi3IxXTBJAD/4xmwknifTAscwiXBLrSML2U3EMf5biIz7ZGK
ecoJNia7IoJIvXNhX62TGThJIDwBZejjhOvA7QUx+IsekwgeuuWNyYtkef5jW71mN2vo7EKtRLcc
Uqybcjl/GQzkAqxaNk4i+kbwX8nD7281vnodk4Jts76+oyiG6XCRaGXpHO4NzP94YCWOvngErNTW
bv4HTQh/fWg7ohYZj2iw7gedbiFTJv1VIbq1PI10nWZob3RfhsbyIPLfLlv6Ua+dBV6yET2Ps7dp
QNpeBRcYb79+nAOO7I6Y6ft96KE6gmCbRU2D+Dw9JKxnb5+0CGRt0LqyuXafr9C/n2/1SMObxe9Z
SceegW8x2IbJceipS43YR4vDOGb0SKvSrTeubVFEZp88iPRHkIU/eAocvV8m3lB2NPxD9y0uuxuI
PoP/kMtky6GbCv9jZ8rfosAsXwwWdxok7diArR8uwiYW4aSpnS2g1akxaaYkKDtxNMiP718DIU9g
4R3TzpnqZAulNwDZWe8RohUc/c4Ojzcsc3UMmUe/EkbPgftWthz0s4l/Pp2Shlb8Ijr3kA5kNYV5
7FPaIFVjoafpbuU6GZDM8WME06aRSyV1p6bKcko4CtNASBANAzu3l4VV4fWLYafTarUCq0DLgVPZ
gAXkSW0IQXHCqTFJSrCBan3P1EpMBEOe07R1+GtMs18krpxTuvn3MoOJZol+zIPY/98yfIzb6lHC
BwY7NgyjmzMAPSABgb5xT47WmSPh2ucahbJKH5k4HGd73kTu1Piuupe8Y5qX8RTA2mhMIP1X4XOq
j17biPYnshGM8zkC/liJuqo/JgXqME0dEXH4x/bTFoRgkVlZQQf6AOs4nY84qeAqmZS673KFa6Ty
8A4ro5BXOIALEodYXS/fQauBib3PT/gqzWHFTFjwHb74NFBAf2LhANXrkbOvIbXbk7ZXmLOPWE4C
QsGU8c9tCSmBYKNbX6X80vyDviWGNyyRx4gMFp3IuAKHInTPg0c9ZDo827y/1TXj4D1Ql5HXJEg/
acS/DBaoWw/5V+cBuNQ39AfXBejxlBjnvobM3Yo6xGQVJCgg/msFGKcZwo3T5O0ptJHHm0Ik0SKo
zhA/Mh/9zL/ox6H3G+aSRWErOqI3nW+3rmJJtJcrDHeN6AceawZD6bXxh2hBaAoE8tzdJjTd0lVJ
3/7VDe/BVyETfD+c6bP58brvMR7YC8XrxgQJG/Rzoi5uCvD7Tkjg81uMpiza49M2kEkDr69l4sLY
hA/dsht36nj+kRaXL4/PZPbYXjtZVTRbKDLlpcQn+KMBkNxba6co6+ZWDfLvgTcj9Y0MM6kDuOs0
VdOXBIwHL3XipSpNm+jTl4gyq8Ye6XWt6fL/FUZfpNpyC9DojK8NIuzeZMKnEDWrr94z5cF458ER
Up8s8xdKofk4yFupiBUNXutAM+AiRNu3DXA56tkfDJHLGETVn5hUbWHhN1s9/e4lMfOWiUyKb2lV
QOAqpCJ331jAZkIMldWrSyhlkdeYAuZg+OA85w5KAeiqrSviMGEk+ZA6qsjfUnV3c7xvt6qR0TsB
o461JaImBw/LkJe6wt664kn8Vnm22CdHYcalz4rUxmJmaOKM/nAbaTt/mRQruinuQr/kxhggjnew
bSDA5LXUwhfIS4aB7a1KWjqkvzamusA4R0mabZurRjyLO50THFcb/iFvBXzuoBplZ/JqKAFiu4No
1k/62EyeY5Shq/JV2IO+4Czu8HAcL+nt2APyt3AqTpoeHtf+cwMtx8S3g5zX8YtabJCma2/xoF7a
mItdNBMuRd8GiQk4+GYB7OcPtv+Tkl0kVNC62ZbxI8Omg1cJrTO8eyjA7PqAPwQh+R+Z2PdLeIZ1
RM8Sve06yEDV3iuPwkY1ZZ5gMMRJ3lE+yVdPHdUrtFbAzqD5an5WEuc+E0Vb6RuZ2CtFK11pdRr3
bnLNwcpprgJnJZLHiyUD4xKEAs39ewndfG8T0DdSwP+qSSDtfZcbynNOiUpdyPjB05cmCSV/iY9H
t2ls10f++IpW1+2ljH/08yMGwkG7uppOzxu3m5jCa6uBu7tofAfcL2G1+LpPILUzhFRSgqmyOZ3s
9qajw3OpI0Kf7An7hdF2TDZpqEOMw4WtOLqWMj59rpvoV4sFR4fQSrG9J6ZfAta0R+6TZXzslZds
fZZa0goXLQoHHPAXQsZFV53nfphuL6oYQe1ffgjZLdVE6EjtNW0FZstaGyMdURTtzDE8UXpc6tSa
yC/3HCEcdC9IoCXFV7SQW68a22rJyLlYtJl6PjTLv65tpsJUgopJ7v6FD/5MFtzH5AlHKp8VJryA
wR30H3POgjL2ewdmn+Iosffj5RfI1Pbpo/EILXbNyfpO63MYoTYStLa/mbgNsFG3Oop15fQkaCEp
ugdxlT15VQN15OvxWFTReU6DdbMFkAJgl7d/jMyyXHIaRY5Trx6Ihd4cnlxp/m7VTUNXgrAXDpxx
rIUzbhSFod/mM4VuGPs8N2J7TMMa67ioyNsyu8/fhbNmLVmQwFlBqx5Y1X6DwkJcwf9kvVFCcdah
pR1QkUWWwB01oQ8EckchymqMH7deAl1upRXVMUc+gLRyFxj84ScmTriAyuhFnQWKZsLLMRNsp+RG
ZiAMT0kyRAWWFf325yeXWLs9Zn8POd591JuiANoUa+x8s4YaKL7HU8UCwR4vHuCIVepoEOszCy3a
YFBCbFFoRE//PF7p7vlIi+cjiDW/65pOtCOcFkoAJHBd2HzetkfvL/r1G6ZQm9uBTCL/EnbFB5XI
95VgCbpgL6H4d6K7HstVLHx+YjBK/xIpRFwIX8ykU4///53ntu0EzF7W3QMxfRbzEHCUMK7OwZ/j
0xh/NJlLC15SC/8O6HY/Oa02d/fyIhkK9Ao6JWjEnPdaPdnVfq9qAogcvdhZTQ0Ddag3QgT45Cst
2dIzgGO0PqQ3SX7LcrHWXycNPIQNV6VQbM1G54U3alI/BU2ltwqVylOZahDmzFngWGLEE4Eq0a6y
gvDCnH4Qg096ZppErvtQst4XAjWKREU6B7Zr2AUeznTN461JX6xDG6BuVC2/aXbss2fTZNu4Sb8J
BszO/S7/XmPTeUcWOqi9gMjABhg7iVAsdPGQV/F4nJdoAWug3L88yec3XjeWDtZYulAbyAp/aKBi
A0YiXw9oo8pB+9qnx0MmLEf5RdMuwijVjNzzPHzL91/Ay7ud3F/9ThFntv/bNQrQ6UNoLvOan9qB
/dE+KQrPqLTe03wiLy56fAfQ/Fa7HOowxqLTreYdxCO5PyZalhUrH0YPdCrbi8zP09NJG3h+w7+6
ntxf+ovjLMTbS0aVYbqkLkxbBGYz6ic9rUC01Hd1HHcTUw4wBrYlz1RCK9stUCXh/++Ee93YTBMG
1Woh0Lynsy3P3S/gqCxjOq2CbqxlxxwXWNhUBLfrdUoFNp1KKQs9h49HtREDk/+zTxNaUuHUH0I+
jCZFSbUyizvAirDMtZvFKcAo/XcckTF/ztHqdoxRzWi7TLEejWBpDnTh+v52be2lY/CllFNtpUdL
rqQuHEzTO8ptJxQR4g3D2f2v0+0/TuHNbkoR8t55on4d8Agb222yPRw6hAdOrA+g3cJm9hIyAKKq
fTkSJXEBRAz86G7bHAYlJVFIG7IzGUtvaNe0TQsZqTlCZ7KXX9QaWFxnquezetg0LAL+vP5Y1qb/
Q2dYl661JZuGtZrJCKHU6vEJah5RUeKZDrgBByHCKXJ28WiuDYKSRT4u7t8PYVnE13kO8Vb5r9Br
xVYuCefdjZTA0ZBVfCJFhVjSNkwB+KRStJ6PoqoFNgh2Q+zNQOMz1t3s298t2FMfgQI1fHozXlZt
i7EDlVimHL2PEfem2sYkhedLoGHGrm4BEMTC/izb7LYciSbO1QehFkTrMnNev3EGO36dEPzeg0tK
mPqvJ6jejhtt4h8upm/tzL6/aXl4QVm6amL0bHZR2vdQnsk0jnh3nZoJnUvo6iFFJI0+6wYHlVW5
f4hhQk/WwztNpzS9ck+7/fNrZDKQ84mkFb5NnurJLYJT+F6CfRSCk5MhrnPHhNSYslG+3AwPbCb/
v7r6T/m4zigdlFQXzuT/SfHgnfBlb/AzuGQdyX8MdKz3P0PZBgyzC8lBTOVzBHK/6qCpsax7zKDu
2k3+cgx+3suYk6yXgsq3IYMgMc87NK9NbAKyBWkTuSJJCiilkjBSRNIVTFueHEwKjDRzU5luMPUP
wsTmeryfNTT4bvN+OsBk69hPRSfw9VsxWX9dhMmYfIpW6qucBsuqyfMzcuPKfuM0Lf9O9ZLpjyzc
C9Qdtc4ULQ2HQS+w8EErUs5cevpayN9g8sqOir8EOVbfMD/RuQkA3Qt7X0p+Nk108HbggS+32CdR
XR4/YwvjGiZyrjuxojMN5hgXVU+1g7GOq4zSjYPMCg+sP2oI1A4eG3L8izRuqsekfMI15tSnEm/b
94YTYw4LW0dL/koIRNwM/uhuW2Ea8MvBpNV8hWTP6pDYveesjAaZfFTb2QXw0X7qsBFOBsvplV0r
x+A3/30DxLjMQX8LFYcMbhm1L9IWp8ZmD0WAgGv0SbkHvOBR1xMEImQljurK/GRb2RCzQZtEkpq9
k5wui18eAQ9NJe1ymSEuVq5FhR3eD+F6+2ToLs2XTUQzvNfcTA5/Bd5uRTu8ExuyVZcZe8c+/yXx
L0o7A3IgPFEVBQ7u0USrgwvLbkfxlVsRyCLqMwsuUbrefKxsRZtTSqVgAQ61qZ96o8OXcVGpdIln
rKmAJOLvZhRL6b1wFnj7HUWmRPQdN2M3d/hccowbtbwTmWcyrOCJrIAHaI8pHISypvAzZzFbjzP3
mguxf1XkyvbU7yGMdirEDs/eS8NVUfAGgl3VLg5Pm5Qzf6NVo2x7d4ngqCwCNjAEecGWp/yEgbUN
dSlwJRW8RLDWDHxVe6lhCxOOB/sHMol3YPAZwh9mXlKjIt4PNAMHACiKh3HnLFjGH6ka/DuIt7p9
dspp7cTZKzfusinn/m0m6yRYg7VveM4v9erj296kpdnNiMjGhISJV4NVkbga2zdT0LalOrJkW6wJ
HH+pmMcPY4cnYss6uNFea8W2rRPbmnn/RZvyZGjtR0RvhotJW+4AfKbYdrSMKZ+5QNt1UioI0wh9
eAaMgzHnpvGmvZwe+vN3xLRhjMatXe3zDMg6T7RNbcmeULVrVhvJhH1Ngynj9aU8FKVO6WRQIlMM
U0gamg4/HNon/cPkkIGiHRbK3YzImUk/W2E8r3rO/GKn2F6XqK8t0wgtvPbQokQcGM87yTg8OUen
9C2YO9wEoV52HwHsc/e3X0+XBroVYS8tJR93P5rB4Ny9mjF4HuFiLap+8rsuk0hPw44wI64Y5GaX
ZVFLxbXBQlKDMNHVKhzTdPQDoBTZiKVszcLfqvHjef0KDL/1D8M9IqfY4fMT9bEeXa/E70k4Hmbp
HiNHxDVntV215RIjTYLyu+4AipLji3KlCg0n+UES37xOsRdZbi9yvvi+KTTNtSWXhC5Jvzo889XE
CcC27peQ4DU8R3fnliCHkkRkMfh0yx2vlTzRQk4Dp0QSFGuxOAEG6fcjwioM8KWE+WyjPqIflV4g
Kc+CGGrkNBr1p3pgNGsfB6Ihegldqba4DSC4u0U+p/tYqadQ6iHISMWlWj1MAi1VfRM8/sdl2JSE
MGQCz3+ljYLNC5UEWbxUAUdPchYGNDFTVkao5i9pBYBFVqjJ9AKlV0dYaIP4xChLfBWIH44MOnZa
h2uKg3IUOrL7sUe8AaL0nLvmtNG0L1kvbdmWDwNLKBqe6quBAJ64YdYmagmUoCJVrNCkfDR6GOA4
8I1FV5fIOkXtG7MBbUK0ot+2Fxl6qjs4Pztgg6K8LbkrhqiiR4w3r6y7m07hzxqcau7EVQcBWA7y
/xTFGV6zpI+pjucqaCCGMsKHlnxW+T/h3+NECYpugGATdQbTL+meaRm77DvpdDt/ZIgCwqK/a2xf
vSkN9g0aT4RLt1sXcKeU2qSFNztwED+zVr+KfKiz7wt/ubvCM6zLYf26NeJzfo3uRgaLXZKMlK8F
pBQVkf/RykiZN6A6XpNyXX7WbQluja0o1S5XMUecZnDmlqVxZ5+6BOd6sl9x+lTgjAiHVgH7K3AS
T2DSiuX0JGK7PgcD2v2zw1CAci/TTBDPajQG/Z/dR64210m7t4rjcbTpfSLsZoOoxw8SK8NIkUsI
UNV85b7KL8KEUXxUlAZamRycEx+/OLSfYuNAfyCWylhso76wANaIstPQ3l+AAl9uF7RQRiK85O7A
uQc0O+FqsWYUA2UgjgAcGyTEIqbjRaRFMPIPwXWs855AI5bSgzmrjpNQAQ6sbzVoEhy+J9OtWblo
upguJBJkINpDxsmd0rONCOdL73u1Q/rQ/kG060+Lm8tuaEjdDX30qk/Ev+hSJCCY8FjrKhAAgnH4
ZhoD6WmXVG6cyh4y03qcBduA3FmrDX0S+TTTbGduQlt76sPVAi4A95+PCshSKC8U1+EKj29zaMXX
CMlynRGdlyhuIPPhjyp+4lJ+BkK5pIXPe8kZxDcTw8ogtH2FULKF36xXDapI+Ui7mKDFwz18hGQY
YD2xnKPbLzbbCe/yZj14KlMBg3wPjY5gg68fwEwdO4vyAUMy4hUTB6BGTvQgj3x7AHftLLt2vbyW
4KuLauUhVikZO1IzK6ZmUrQMLPfEuTMjiCgqGoD15vXgAdHWeIhbYZTYRGzjKW7xHAPQqPkm1toF
lqUJKnVMmfAzFhz335rFqKgsJ1KBpf+T/DGxZi4LwBBcTy8wY0Wc2t3lv0nPZwpR03wdZ6cZPWxl
kA/sg6UpeOYh0c7cSc7e5TWudmTBE2RdLbaL8CeKk6e4TqhXbW41WKITZTLIWHEswtkUaju78Vx5
gs/juGqgU/ujfWdySI3+iR9HEwf1vBblxZ9uqW1ObgEs1OojXZDeltFy/QYNsL1kNGDwPw27fj3S
LR4cbn9EKFiVM8h5JPvUb6fKDFhO5ZpZHzC/O80ZIsFQqrUzi5Wyb1cY8pr2T93Hq9W6+mCq3Imm
DJdQFsqXxhUBZyqY3KD/BAax6hMRWbIuH9slxPXV8SmSMOgBATpNMSUaUi6Y/u4ZlDVe801giQFD
bOFvA0EVOg+By/qe0aY1MRkTeoYmfr5B1JL61+xXMHqFSQ6q705MHoVo+ebpYmW33EzoCrMx8QGr
eAmsCYbh4gPwt1V7uHOaT8X/rh6Auike4cvBPo2fuPWqx+zgCcxBrPuGT2dAwSMQJkPNJKNplEU0
IDd5pEiZ0QlAX48cGhTj8c0m5Avktp33UeW4LMMgqi+HqpxyMWawOCLmI9g18Ev5IyBWBV/OGDv9
8OwNhwKWaZV2W7RNlTZyjELhhHnJMVqnVh9fKfCwX2y60svgphoukYaNxgQfzneYa2Od64Jkjhzg
I3Zssr2/n67RC1O8Isu0qqsyYYNqcnL6nFQ4bRPD67Ka03LVSBOBcnGInOgHDF0Fcxa8gRC29M+i
h711ZyNMZcl1aHhWANaMlHi/R68tNNf2zHChEcoI2l+y7vw9cYfnYTGMsXjQzVzGkA3wRF98OjbS
s30C8ys3/EnvziWST5GfqYgI6X1i+Ocm80UJHtHVlNjktVr6FA7IUJdVZP+v4bGWs6g/BEg1lTNs
hxMWGAQMO56KmT0qddWNO5kML8KP5ufj4HDssGJKGs3gg6M5+iZzKRYKw1MMgIdjUNAL7NTb64YO
fnn+znKwJQxUv7qlXiU+QdqMQtWen5dr5JmOAswgCtJ82bjtJEk9tQ8ykMXPcaxEC0HeD6LVah0w
VrWTL5lokJQ/NlwWjPYsNqAq9mIDHzXaKlp0jKKf+kRcx+kzhWYw8k1nL9MvqHAARYpVXSjbEaTP
X+3BoR9BlXQJGpAk/s7aTi3LwOAuQXrZYBwebp2IeYGOlyz2mgp1u59fJeQ/UCBBWg99ktrlSdRg
yo7HSjZmasB4L4E+oJsKudQN6o+TU97v7/niL8EAW2G5AjmJZq1gnkR5TKfknX5cUQ0v8iKUfmxq
AYAOoycbfWq66LU+nCx+DTFsV99/ZAq9kiIrMKx92U6xlQUkb6ynXPKLrrCPWty8DJ+qvyKVodoV
laolc3T9uo5EGeSowwBJHQjwTNAbP9hBkn9Wm6d9YeBOJj7t0cIjRCtbvgQt+DVm1N5qQ2XzIp+r
ykqjxWaGWjaXGLneb6rW1Gf0xKe9wqyRI4XhJeLgEYO7KpCjq+AiOEr7axHCy7sjJe47Gn9Hbw8Z
uPFq7uN70rDLiDJwo0/lC/LhLdfSBfJB4bFFkn7p/6bfH7/EbkcTfXZz4A7tL0DYZFyUwx8rwrju
DLVecET7WyMXRwvio1MApOLXgOJitiBT382YZk9iMHjx42Z2nAIJaXc1ICSXHXpUZfdNEOHxeRnv
eDuuaesO29+d5omta5Hhd6zd93hY1exfrYQm9EPmmYWzG5bDjigY1dcQHSyYIhTXQiwhBQQsVPTO
pyWis+W9tWxaNl2oE56KOh0ps0pmrQyaI+KF+2pRuwC090dF/zgpvPHCdqBEpA5vTHs8+0zf4bM7
rwoI8gA8D8tgQTlJ0TGFdBwVN4GmibrkCli/c/rEGjWdraw4u5EAKpYXL+KCyifPasz3zLZsArWx
9moYn7WCcnDIgz2OlFGXBJEo++2Me6UDorCy6B4UjWBBiZjQwZUENEA39Q7lnucsihRNJG0dQZGE
ejrAH9B43HHPQHVn13mqn0hp3sAUxUP/oazlXw2pog/FLCGEnlAvg+EfSkiC+uURb/w409AXmAvQ
xur8rc2qy2BSEEvjP/d2DP5HthfF05FIfaqQl+XBfrUWenpdHDukLOfwWxRAwaNsbroizMcWIH42
rntsIR5GoXx0o65jkJ5zsARJnb4cUZbk4pcDvPMIjA2aA+tHs4DkdWfa7/9M4kpY1sZ0/Nd7SwHL
0IiITMZ9lfU/5ulxrzjWeifq5Ap8gmxiLpOqirYUltDCjViMwAsvISDr38IOXmNH6Y9DNOuosAqu
rmgxWJr1uR5BK+qKVIvbjujNCjy/FQcwBmuRWBXGPrOyZYoBgNgRjZrtsK0H6WcMkj806XIyrhxE
HTwcxQz49FiWUqdbUmP8ycgQByb89up292t4TlWy9ZP1OuOnINrG0NRSsGab6Dpnc0Tma24Df7ba
LmqoYAo8M4YMLXOdrnMEseo7PWweWo/4BLQwtpmMGDDJeQQVM7GdcJcIkgzQAx4LzYg2W4Odr5Qt
QiTOM+UuT8hcg5GwjNMo/Z72RvzcJB7b5xvG4XD5FdUo4bwEu7IVkFts3y30abxZk47dD1kwlDrE
KhYv3WqpsOAXmofja0apkgufFpNWxg2dsL1CZbQLS68V2YDM3MNJaTuXGa/sfCsS36xoiSG1wXQN
uBxZm0je/3rxllMBGAQ/CP/RwgPAsjybVuJBUE9wu601ks7/8JOCoAU8VgQyYm1WD8Mrw6V/qzF2
X1gz6zKi/r7B3ZzeQvzGOVIIQiXxta5qPbwp9sZAs8xR+ZX4UZP/d8JYcwoToffod88Zncu3B4wF
79kJTqpJiU/qNzKxV+fiwLSbdqXk4Mabs9QvJMWR3ZzQBNyBXUy3RajIjB4FBWPtMqKvBIB0Gfdj
VYaW25wds0iBzFyrr4yM5L5dRZ9CGjnKDliwTus21rXYWQkLCLdwtK93W4Anot3w1PQNI11Tx7zp
L9lYBFeFYacRkAx61FjsulPgvW+/uqvFFhMrxUAj1ONjTalAQEJF49LHmdvUctTNStER0v10MWD5
TlWxlp7Pa67u+IWquwuA3pSVj4HONr/Wcc0B6zba9nzoQSUi9wEBhXqyiYXuvpiIxh8PXFDn/r2D
YiuhTelVjMP8dUWUHb4R1jdcTUyMGaXUxcZrGR6y+YYRGv6zQho8l3SE9ESBXxzsLldEiWUdQabk
lVHc3xhLIdGNqRnaDeo1kGN8oFczATPCHTzInfe/mJtGNgLoJI+oggXVbS6ca4u+TExmBfbUzDUr
s5pQQ4uW8/xX84pBTLTndnEc+fvHCh1czXxH1VN7hozmmxosYeLELZ8pEebekR3CLdvnpcube0yS
ojuJ82m0IGlZKyLDE96DTrhjn0k2aGEHuvsZy6W9Hz1IChSdz57Vn3GT7DTpBptgJux4sT0zLuP9
Lh6dzoHUFhiq6xRRYoVL9cp+ERqLAICNWzZFfPwcW0H/24dDeuH/mTuoaBe/+7Dv+LREoiakt28K
DXAM95rns2gBg395Ux3Awn4nfepPsCFKAXAsPRFkj5Z/4diGimhTcnJL+Zrxy/gfoX+0FLIB0i6E
x01W6rhAm3u6Q60DsJhvZ+qpr1ODEDLGaXRp1hx4L7LHZDCdRIiUCwzXtbG6vJyNXwchpyMATaYN
cdQgRrPOkYBwkHFiItpy+YVEjpcKSQF+WV36v7QBimpeHmNYPHzsJJubX69eMOurZlx12PR9pv5l
94eNqyP1yKkG5lJ0tV9F+nI40rlIjWh308TpzHc5enOcdVaD1daUJVF7MLHBIuXItTctUa3X8JqV
O5hPgs3Qxd5JjpOxj5yYoVqNXH+ox32RGC5vH4EY+WG2izolUGq0w89n4LhJ93UkIFzb8Y2cF2xU
Hu9mXZGbLarjDGbr0k5PmovCd+BePr4NvXNnRao6Ow+sWNepiT21MSOPmdPOQfukxhjssTcLeFL6
tq4Riekw8RAypjUeIHlp8sNC2SSqe6NSuGvJYSl1e2lSpVvQNO17/VnT3C6BWso0+vjf7w3d9OeS
/+gt7EhLjLj9XlrxCWS2M0MnaQh4cjtSj1+hRpvp6rigLKG60Ip1h5JOJbchV0SbVRYmKCnKSvOk
Gn1injAtT3qADc0lpYg/dlAeCz51QGgKZmrORATIvaIpwFLQwcoELZIoTw68ZQa4eldoroXyqgL8
/vf2Bv2olcHsQse9BNZQ+Ica+lwntCwHpzEuiFdlFADYViSxGR1AYzDS0nP8Soi2KJS6bqSVutf9
AjZPHu7nZxjsDUuPEcNZtZy4HSewGyIVfgmSwkuMkjjibQtDM7EB/8jxycXLeoH+SR7Jv/JdWuXZ
2CKZdtQx5wG8+kuyGiSDcmaIhxlO2CGSeuIaq3T81s9PAE4mrvacc5SJFnCZayiF5AFkRJuqKw6C
xJO+/EZUOmZdcqvM/Ifk9LOmfjI+3hNCIewZUBeI34pqzaKGh+2yXPfx/Itc6lyWGH6JVz2aWTD4
Z9UoYxwSXKv/4RPieR9KUJ7ljjb1M9M0Lh1EZzuzRb/ICTGADVyWq5zxhuSnKcRIGA7Z8Q935uRi
QNVCoBNw+Xo/NJaSVRPXbjYVIxgJcS0S003D0gdsBlQm+8Gg9pYP26n7MKd5+NKNpq53k1gL/iPu
O2dI/wWqL/g/JaMdytKo+fAA39rplLGkyKoP5Hkc+g99cwvaUeYK7iys+wQZeZlH8gJWwOw/KRDJ
6mME9tqezbS/U2KbyLL3l7ZnJMw3sF1VVS5CCndQmVEhBtl2mKJp+qIuwWP17JbLa4VfVFomiYKK
4V3a2d9kcYK1sxY2Yf8c0psRpuaw/H5twxwKnvWhTK8UITLlVCKI+2dA/U8ZcXd0U2WaiLhIGPi5
MTn5BHvszbY64ZAyQhBYhsh93po8HgiyEvplGtQPZRnqljJiVOyNk9TaK12bmK5/zT1Urg5dcRDK
JDzSRguavAxiPeX6Wf0qeeKYoZ++2kDzCrDS0l+T7fflMKFiPcH66BfyEK6ftEa4jqyEXXz7WPfd
udTQPBNPnE5M7cmI0Mt8pwDDkuhc5NuyhAPIC2tiX53VD98K+xE0aIJfLQyAB1NlAhRAjdnetco4
penfJhaJUUbga5TA+LTDgOThiFvC8OxMr09QkanDbIZyzLAG8ATqwELcBiT5yYXGAWE7Ts79bUP6
EWGzWdSpCBPXj4cDTllaGuJ73BXc73MxBoK5XIRCjxgKQYj4TpQwuyvAZzaSpcHpHd63WOK1Y7Fb
qlKie92nljZgEODuqe+WHhc8JBz9535THdxjnxkKzZBO8UCN8UM1qJ1SNYqgE4uKboo35UkTaEq5
bydalAkMSM6zrXOWoydw2VVjaM2BjcsDOUdH0CEBUNSk9KBa59Oiea3H8G46vaGBT6FfkoQX6jMN
TL0cXrXxaIoMQ0wfxlyGQtIcSA5PmkCLzoTHy19fMZPkm/yPxtwVPeHPsteIYN1IdCDVzf0vhECo
jPrk2kwXj5NgoWe9jPQ5eyY36nNg+af17W7GPHOL1C1HLo+OnSYJxbdN4P5wjnksDE0CmLsfKHg5
t4FS8GgvVl7JWMZuTOszOd+bZC9cm0K7wAJKAHTqx0q58OXYv/MB7OnGRPnLZcjDOYX4kaarQY6P
ZXMqc/ELaJQF4ZagV0RmLzVfSrsjZt8C6CtQYLetEMydlhD9ELSrE/6P4nGY6TrEhPI3nhnOlUqQ
iQRKgBMFFvk+AWHpRWe4KERoZqzBUMGaIj+lMTIHzDDgzUww5uTnMDGdXVGssVj/2DFuQRnc7luR
++W45VZX57cij/iHssVenBhEu0Gcz+5BHouxLHRy2kOQQaZxAm4u1o/EsMl6fu9lTK4QjUUJG2y7
a2AEa+EOG01FZQuskVcJhmP00Tb3gnvtWfJbb2gnnytKiNt8c1h5UXxElxw/UX8AfQkIkiLyFkCR
wGx6v5masuCEQr1ubWGPjgjQanHgVI25ihllE8naWl07eeba943NwE2M+m3JIFWA87eXkRLO2QBM
sQhlxDl1dLk9dLKxqd033C/J85QhjzaZIHE5ANZXHNb7wGxxc+4B4NWEZhCDVmt/jlv6kEK/qZOz
jhfrYLn5+NsyosbEwrErTf8GC46l7iGSEa/hVVX4DxHspmGzZhtdsQH91DToBrDSpg0IP5M4vFtb
pL4K8KOpY+2gic7HARD4s5q8H3dGFUmIpF7p2ZyuxiRDjN9NCJ5cBGorkbqg2u90dvOAbYf/LhPA
9Gw6c/CCu/46OcmCmxb6r6qpQuKcdl92xysAotM1BOt0Lhk9jZVAiNv+6tvCkBLLVpCsez7vF4xK
C5gGP/aObZq3jLP+bvAyKH6vGuFjrLc2m3gJfOXePclFkdB7GATMbQ1a2q1C/DeF48A0j88uph3+
cyxxOQMp/XzC65tO5wXrhkJAH0brOKu+Ke7CcOWn1WrskKZIqN2QyjRw1x/9Lq7cu8FZPBdR1CBM
ItJE0QDQrnji3f1lnGfJ5CQlA2c/pwBQoQlv8hTHcpWs+w0EYMGh0lelGIMRERhneyRLobOpgCS2
tlH0eD5uSOk+sc7Zm+ogICfK5sRxYDANGWur2cDnDo10Qac9wzD8J0CwvdYGaP7/dj1btkw3jBOv
J68+DqVDnjJ04ZwdXlJEZFzkhbVIk6CVtpWx7kzCZc/WDY7NvlSZJ2xTdQrB+L80A28QiX94Wxko
MLaXTwCKSGsiCvC8bnsoKVPydLlK3pzkizrvvlglN9qLM/xwIzdF4TXJ4G/2lQz44VfFxDv3/5Am
wr8QlJ2LFw3HcAWa5l/ymSGef6nZ7vc/wEPTOxJwFP3XgKXytZz/T4CUGjtoirxpeISWlnMIpmsW
aUsufJE+64l+TXcHalyQCLtJ6SKCzWTsSYBzOoT+gFoBXgdWgDHhmp9tDAeVfQ6dpFvHoHXCF4ML
oCQ74uA2NtOkez/cmH2lad5jEQ32fkj8jfvo15/NqWHOIFZSHstzNtmFLAADs+kiHTnLT5HueIct
zX4DB7ubvd34v4eE22XLfHTIgbX83+zTzVjbFTt4p0Q8ms2UgSh7BCgStPE2n5KUhFGjdwIFclyb
05Dv/mS77TUmad1syf8mTBaKeqsgPCz3cTzP0R0tNUIJ94jvSIR3pK79Bfayr/atCvGWn2EwHlsn
sbUN7m/omukSvnV/hx7Txda0UQPtaDtHwOr2Uwg0FvmjZUShwFmg97hUmHvIxOAOG7whD5vUkoGS
zg69cmPScJQufhyIu+bWuKwl0/9fxSdMO3lhsCUMXTTh+XvEM2s0z6i05gsBWs9mENWLtJEOi6Yp
r9mB0be8CVBHbHBk4ibJ1EL50uGKNjyNIRxik9XTVrRCE2fdwuoaEw3AXnQvTvy/Jq3mSimBjac9
Ow2mBf6u88W97QNtKDUILOfeN4JTe0n4tLS5gRLS7hAYI801kNCd/iLh4Ks4SHNUTzfAHL2HUxjH
D0IIgG/ja0vRvi3zZzXAsvRyxEF2sXEXyCHuleV48VGAH9H9X8g9sES1xRLcRuynjfjcmJGkgflY
KIMCPFXCcUV/hHouvzz5nkNIl6/hB5jQKl5PE5AV5jrVkA+vZkBN2DGviawYlfFTUs2eUQ4ZX7T/
nDBFn15N3HmAjIsH/+CE7w7srgb8fawy3oqAxW1Y39JNfJ8rKEdzbawmV/borB0mS4Y1z//xFkb7
O8nwCDVuRoKcY557XXqkbbQDi+bja8cuaU3xv3QFG0mAg30f1oGEwpp+Q273hBZF+cnR5b2s0Bqi
Y0UMsIQy+g06SkGUgHmkt8DMwA85pZ8+Tpj0JxOZ8z30OalnlGkSiTItNK8Z0BblrVJYH+kbTAG7
g+18cXIQ3Ip0G70N6fzuyERUlOtmvfj8gbJ+UhjGd91eQ/84toZGhY1+s0zoSzCpoOXuwVRtZmBQ
4tRWvDzTnfLuEeFhQQME6jTpMmnkD3JjFhMfFohgXEs1ptWNGnWCCxw4OVYH3zS6YjDm2zcVxGMo
qEaiBUPur1QMkkcKuZ3GE/PtdUCJP6tL5qZeQzHktSk5Y5ouSEdWjoJ2pwDpJgSW66gwUudnedT9
qLEbJkA57fiT+HWoFcxuiZibAgW/EBvcteRjYz/gUZTUPRknyXYgsfz4TPaw/wsCHs83ZlnS3acl
qZuk6mk38tESryjpRQU6gfwlYlz2jBe5ImYHZxbKveGabLjt48KH+FU3IGGe2CR9bWUl5qBnFd7/
idscTkxKh9pR5ld+/QaodwZUBqv80sF+Wp3Tmq9sW0jdToY8nqPWkodkV8Da+PLOvfVh3Rj5Kqf4
5QyAV45zJ5H8o2oT3jZRSA7ZK1jS0vr5BcISATU+XXjs4dJA5mgKiZTWlKT0MRj+DjM4JwDGbwK1
9cCwfv/nUSPmFDSXSBfs9ojlQXBJ8F6FVlJZgyW+obxTXi+mLfuUumLIpj39qJ85csvBmnTJBHfT
d0o1PjMZf+S9qzk2sS4n93YEdWi7C084xXpGOfqntkqz8b8MnyH0u1jd+wtdnanics4DE/n12mOI
+zK0GDzT6x2H0M9msBrMKEjotHDtbY/sRaN6YdXWC7lZNvxZYid/aQByLBNWhH926eMfcl5L2UDm
wmmf544CAPnLbLrOGpPp77A1KlRD+QzH9K3BC+CbHKKkOFkTBni/cGdflyZXxhy6/OUAcnQB1rMo
Pn4HXh1KJeVk5FPRbf/H/lNy8w56g1Y5UhBQ4OmVBwshc5aMtUq0vPETJB33ZA9rIw69qPerpXrI
yO8CRM1w7srBuax0WpOy8vTyf54SBVzk+EN5nPQCEH/S+8XJQZxCw4g/iDhnUQ2aoBVezdjC+faK
c4gzJHlpn+uC02W/b8RJR9Ky7WqkaWidmOMKOxwXQMQ+ylvaQqaWjQh4MS/C0X2flCk+rCpza04J
FoVWiVoNhkhzCK48zfBEL+4GBOqpsffEdOu84YjrcI8BRMtCMcwfUUViDYGsoWnGB/+vhMgJIXZu
CUKmJcljt/JDWcY+CxW8gLlKjS1uh/u+jGVjECsemQXWovGAfCjg0jHvK8S2JO6FIGEFClayg/O+
1pkn/0S+VCny03ClTsxoJusUg+YjCPyZVnmyOy8+eqi7H5RFLnCH8GjxznWMz+SqJxAZf2fiuLa8
4O3oUc4SynTP8ZtlgatosGvs8zLichHohc2fQvt0EP5SrL1FWvSm0EcgbVXK4kAncnD0YPlPJq/d
fQuskInX0k0fy3Ln/ggPA+SqG/tp2v/pttqj2A10iNNVBIsxPErCG5Rq+k59eCkRyW5fymzggBy/
IXUpPn0X+DgleABY2c5BZHCuKkZRk2Imki4oYnlIOWMBNgEyaOF5KpKCbLjwq9y/SGV0iYpgL8y9
wGWXCkTPWM2wY++lRTKJbv2pzDJTpeGXHbgqHlxQSyokM2Mnd9J2hcmZudiyR7wvraYGILTfvMky
OrQNDCbedgBGvAXPr5EDiFOYca6mpe3No1/hQ5Q71yRPp6OFVdr1aU3/8sn/bXWvy4S8oTXl/uya
gmyadI93VFlaFib4aJroLrh8ITAyqLViPasiZ/Bo/l59XLHluEJGK5E/mqG11OXyy67gPfUyof6O
AXPxyRxxJ+WK6FfPyzZ+J3wU6Jz8NBSuspQ3xMVa+hFJvK+CB5T/YyMHNy8z4dtSd3enEQtq33T0
SnzQiEJz6032CpZ/aR5tqiMrvhSuru9OqMSgumTVXiZpDBW/+xWUe9KzEJYJGCKGVCyGxOwm261A
kAXp+NRC/L/gVjCpTfOZGagoZr0ZH5qIMW4xOnymhWERW2gACzQZmLJtrDWHCZvVa1V8vIypaHdw
b4+PlsqJQW3OBYidJiP8mdRNMKUgazMY8Q7sPAurS+6AwrZDR/hM03qPpod+oiGLB2hSFe/t4Y5B
j54iLu9UR5ev2JUKapXczNVvV/3MAeQySzqYw0zsmo5cZI90gSrIGXroyrPervRmvB1LFJ08Pdwf
bzni6JJaCjBvTpc1sopI/qe6fSBzri+9i9sFGS11JvOsuA1zVv/zJLy7x4Ddl8jXkhKbCIh1H7LU
QVPL9nfCEJ+4UZlDe4DxunPN6g3PAKBwnPWvAUOqoPLAE4LIYQVGAh5lrBzP5Ukp33CLQB+l7w3p
2vgibNI24zkREWWp9v0u0pIZo0Z0pqhq7cF2KhgQ4QZXNBg6DMzAp2IwwK6p+m4DX+vc21zGyQWc
c5qiQJcnBN27kA1lqa8TKVZTcGcsuEPKKTfuQDnk3Xg8YjxFw2JHk1HqIdbf+guvivjXEsybJlcl
NPqzH+GXNiaMmaFsN3YJ9FGFjn2+vXDOAHAKl/9hgetMwYhCh29lAiq3Q/W5XZo1RGU1JBybeWVp
egMnwN9PM0G6IE3/q2iv9jzkuO0tRsgc372f/QVOThsubpuqK/x/MUxbLGGZSqY+JIFNIbx6L7to
y8euP8XIN/kGPg+cSzNst5gIwbtkRICAo5LNhPNrwXab0blmlJb0uDii2Gx8T9eUyjp4d8f7Us78
c4n9VwTcdOdAVb2pxCqFDXE+dzlauX+dBt1Ok1IZAHj+VQur9hXqJ2rb2F6yklMwqBPCHhWuFAbp
lq5/XXcdYfJzmToBEfodHZ4hJqz2Gli78kD63DwHcBaQCzgTbjxOT9YT3U+Hhrfvob3oz4pc9I8D
AtoDxfSiQbOZI2qmJJoRUvOm6169XvsqlqcnBGNyYkmtsAugFWZrmNCfaqi7xVUw1FhYxQXtSd6M
9xbiWOa/BQa/tNThOQDm5qcbn0ZFVG09tjs9Hg3T2x3HQgdagJksTMpEha76mzZT194xYx0uhDxK
fu4UaY/xvPsFfIVIcBaaHsV8vwH1Wujsoo8mZnA+nWUMV7uaLhfvofQmpENS07QGZv703uMwvCB7
AnFBFPM8xTz7Iuynv6VxN/6JgIGHSQypyERVfdEOCf6lsLF/c4cBcsEekM/Ddia8jITfod+sOUJk
hbHpmbGe6HHxZCzdWhysymByFAZo/aCRY7Em1Vef3ax2qUtOlVXhQ1lU4OkdvA+ckTrCuvg5l2x3
P2QWRt0BKD1+wGc3Lwyr6Jp+wkoZNHBoaynIToVsroQEZQzlwC6n03P1A0CQ5mmqZ55WDFzJWDYp
3JrVjS3p3/ZHUDo2dn6JIRySVTPVic6pXSd5or4x1altDS8k898gqPBijdLpOrfWtY6aajBt7IY1
EEQAnfLzUJlMwLEEBmept9T19/3Cborcle1HbIfQsB95UL6JRNEifYlvI6tv9w+5dnfan6BJcysP
yjftMYulBxJJsm0k59johP1OG3VbpFkL0rIelH9XxahesU3ejlq0SnjXfzgqLfZmTKS9WR5hnSi+
wJU/CBPqFCggzdmegU2aPdJ2Z2yDfAS5ZFXJEuoOwJTOm/BvbrYx4GmF62AKHWyLWjWYNwi3Chtw
opnpiYzqkapp6HDLHf9wgtYq+QgGuxJPVbeAt42AJr9KHLwOEoSNmrxpQm30kUSr3eNCYBejrJJT
BInYWIRtD1jXwb+3ghkpDBSR5/Uzgw7JsXdpVZCzS3sXV9Cd4k7wCeow26kCPplIzVy9+WAvo4Xi
56EIjimVPlhbmhNkYKN4Zu0wiuYX643jfKsJTDTCnXwpudgNdiIKn8yEiyvmgZksB01kT53OaQnx
3+ambW337qc9N7p4LRuAHmPtPu3sZfc57t1obo9Pq15+mumDl0scF8Nt2x2GDJspLZ2tOiZc5V0D
rOqrswafK0TofDC2drIlWjEJbqjPTktvlGDBu7t4uK5cvtmEajl7q38oco70cP3+hg2OtteiYCBr
yfD0Z/ErPyFqvOLkLDXnzX5JeCOGAS9DNIrcVT8v3ldZOz2pH43kmTPHhTtl/0VIWbGbjb8+xtiX
uopRsaJXaCj0tEnxW5ZahxAmVaj5YvWrPJd4f5kGGXA7FLpMUUus6wCUOcgOhBC39GPEiop3rWMa
CvJoFQJZiiGoSFaoPtMTJ1xQ8YSEYDTV1ugyUXEgQwhYXeD7xkHfsh5i7mBQ0NNsJJxYJ1DYsENv
GFjK09y6oue+GO024MeG9wmbn0meVYm1tQVF3h77aE13Pn6BBCaNrUIb+XUQKV14XPRYOy8DLztn
rzPd6ZgUIDsWrEMaVAC25QbSqSdL+NAshJVXQRMYRdX4yOuq8I9B3g/87rfiqT+Ff4m2EjAzoKtu
40L2rt0hTFUl9TOXvtnOFZWuB0SgfgIa8vrsswJ1Dc2KVG/dUC9ayiJ+63zMJ5E6lGmzm5pohHPH
t4dTKuK8A77c9KGF/MUWhuwR5ym7QJig3w3MxMpU93t3fVWMVyZFRD8swe4uVhPKeEJFCaaRlHN6
tUyFJE/7e5M9DiYf2zUGa6D/nFvMsSCB3q9hcVfRIbheZNZ0+cFyBOisYwHUmjuzKsuAq1unDdwe
gaTrrU0sVNiRMmkBrhn7OXvrl1hPipPruso/bTUgZ1n5KW63YdnAgTHS+CsbbDNu2ldvc2D61GUc
yPOlIelIv2jHtSGPqSkOfpBqtY2beuUmVQ9bK4HcYq7L000MODGS9Asc5Nktt8QbAFEgkzQG6Q+y
YDH1N2HKidDnzErJNgSCt9H9bGJulMG7jkMXUs4RIZMrRWOxvKC8sO5Q3Lm2dl5k5Bh8JgGSqOBX
0K3mCDSuE9On+Io+9uCRexDwW8/Vqk2wWqj3zxihNH55ai741UepwTTdBjf83pL+rf5PNbZtuie7
bHb9fAe/ldQGZ24GifZvgZslIdTQwv0ISyua1BS3S6bcJ46tzLWpJk17cK9ZUd1VLasf8RpWJsCJ
5hY02mpUsevZHCcS7X9iZMFftS7Jfngme4TUdVXlwF1gsjN/LhRgbsIMx76rvIy4tUW50TpvDWe2
NGgxoWwwnyldo3DvFNCiGkDV/STKn2h9qZVPjzz6rvjcNl5DwzZnTrk5vIutxzJPRQYTv9QYwXi+
2aACABXVFfdjMv/G1G3gmMUcTf3/TtYpFoWaVlwfvlWgykKM6bk2bS4Oqe97gpcDqLnRgjK35NJM
MWSBfB59UPxRgQna+SXcFLj4ntoDEucz1ein4rPa2e4gPD61S4EYvxhP65Q5QCKdIup0w5VTtzfK
3Nobq3YBiztGXL1iouN3QGieyK/eGNNtj1Fg4pQm85oDzRdFbJygd6Ze9jMozDQWjP+PQCeQPVB0
uFuUg7kpW3w40HhFWctdFkdDj05zU7XdN2W+YmuKVEoQT3MZ07FmoGQ4QIexvdvJTXlnzAbK91Pq
a9TvV9STEFjvk6pLXrsKWjmMk27ndc9gGNNlyui7ShOKgis1Rn2GEEsWJy/GR8wKIl/owfX8K5/Z
KRUQPvqSNLNSwxFSaReXURak1i0yun2/2eEkGWca4TwS6wRFN0XgYj8wmhkCMRDVtdxr/RYtouvU
Unxk/m8V+xj7Imr/HcAImilYL5POikhVPVw7dporqksy9zvwwxJbbqBMutVGQGvgWlrAzEv8G2Fb
jxKkIeWr/qW4apXQPYg9TlCoaE8E4GheYNbc2XaDGVG3xYV09t7xWh5Ak5v1UsAurb1FmTAkJ8XO
XVutk4mGNCuYn/cEO9Imb6FHmEFEsImgl9KXhOvQF9HtxqX1EBYhthlyHQFzou8ZG2RRXFGewRZO
0bJWepZH6wIV/WgRfLW4qTt8Lt8ZnvM14pS5on9W/u8WogQsy9d9vtDPCE1eHxkbIiT2w+3pq/P3
WbJB0wuS2yn5QN5kOGyqkfiwvOQNmDi+ORf4DDG1iKpA0kWTEIvZprvq0KKfwz+2CuHIttKUDvb2
GyeXDdKzkHaoqJdednVl2HdhKkJyy83n9VqrWz1GvY+ct97zIKDSF3oDTUa8h2m9XslmClbd5ttA
6GftCVsPgmv9AYPs3KoLJR0g2GJkVdez/hneoFeNf4p3YpEK2i2djutLdOyltns5i5aMjy2oHeC4
u86kSAOIaPBAN5Z0j44uLtZiSdQo/LNEgFQ+AYAsyfPxd5p59HxHqiTWEGEOKaUHVMJNGkdrhof9
h2rU9CVjCBYk/cR9OI1r38ksj+SJyIVaPezzzQJfjGGzaaYlbhEE/mQTxRSPLmK2QF0uBVBn0kLi
CopUBcWfAJ/0Qo+DpG+/8VHJtUu0JxTUH7NgvEMuenE5j7s1DQ+ZGfMvgbC3DtC7/je6EE5FR659
QELQtKKnreiiF8e4+1+p7cGYz3D69fOSDcyzG1vLlhkS037lS84P4fXR4eYBw9OTpKNW3OONgw/l
mhZ1SKFXF8/mRPVRyEemOw3bpgQ4qOwrTUWdsk6Bi4JBNdL/1cVsru2+IMElPwd9Dn8FGUQZp8dz
snKX4nTvHHX+Ag7Y+4gyqtz4KZqPRvDkK6rD5Pn2vnGGxSVGaLhYDKLHU2Oislq0BcJ/0C9h6b28
WLHWt8GJ/NfOmFq8i2AhoXBkMdQg3ul2X73UlHskYstnGaBKh/e46u0ncXKPLl9vFjYXg7ju3TTg
jqCrtHPAr36uOzAIBJhBtkZ+sD/FUk6Wxq9MPYTy63DbEdc6kVjBhZyusyL5FWLgT6DCizQCDFfz
lk3M4xuB4o91Q6BSvgvuGPBBF9m1dvwO2vNgBPdWHb78gLN6L3UAmQHvrC+bsf0m1bdeh7s4PICI
DGkeFMtjkgzYWN2rFPXG2MJVLffLN2TTr8DfJsOQF7b8NQxH4i2XdVlhY7jqwdF7PmpSYC2MKSie
lMP7kkE7n/En4iTw2UPnIVA8Ps2ZN2De0dZaNAwXFTPCWe8FMATcHqGt35lcTyHyjL6qrzopnsfW
VV+GqcA+AWeG71wSbt7L46Zg77wW1ODb7vzE/qFip13fqrw3W7fA2Oey+1j7AubTDUvb4MLn6vCi
Zp3dfXCm9WdrBy9VcTEOWsBHOOaVP1KhPC5uZ4dKYnB/Pfv5Kf40sGuA7KCEo5lHvjlWQakBGKGU
bm6+P99aT3u7VUVAqrz7SHpNGDvxGmfb1aInFoKDYRiZnjA7TEgJkXs+8+lmRmzU51mwK9SN+BJH
oE0vf0rxIv8So/3t6OFV/SUIXOfwGS6+CJRnvSuTVqakxRVDAlJa9Vdyqft7RD0ad1g7TKAZbtZZ
CuOkLJN/KjyhY42+GYDR5mPlNgCXiPO1HGJDTNckqMVlPf6P+uRfFabd+kJb3uCH/Hc2Y8T+n7CP
rmqjYD3a4v2dJeFlz/V7Cd0FnOY/GdeAMlv5CDO0A/yQVFVqbNRC4XcsU/CtpK8V53urrRpSkDNj
WTMuRPCxH6/xXYZUjmgWVfH8uVBvAF6uk70m95clYDzydg0aYJXzcuLh8SLa+kP7UjxG+clcVHhD
UMTmZ730YLp46qsaUVIN411qMcZKtFynDXSl7bf8M5JLH7fppSLtxPu7GI3WPBDnGLHLTOjyM+ur
aB0mAlGrLnIeMKaMXvmmFz06A+EeXsOiUpod28SG12rOOGDdPrkroA9Bv9Xlm78UD1YdiTRHcuo5
jl6gNx2EwG/fUCXS5nXmo6gksR09Tl/ftg86giBLk+Sg2W5Qt2aYp923JzhsHc7dK7JHOvNinO3X
Y1OCrndglrPIGUQsLqZmLpodZ6PGTx6UhZ76d+PSOMPaf3ghJoI4ax2CdVV2HNYqfsAFsw2l9Gz6
ckVfpHVXgFBDxa8NxjLPPdF48EG2A3VMTUZYALQZI5tpFvIlTfrHXfq2/kYNowd9qRcv3i+RwnuA
Ux7SPrkvUxKjB8Ud1AIidZNnJgl/DGc19lhjMGXgkSdzR9mhyrtd7adBz+yqKGqnpsAKxKcgp4wB
8W6sU0dgYt4oTTW19sGUXWNe8w9MTR3MDathpaY3U2AiQu14HweUM5sBBCCqw/r88oE6jTaOGAau
COATOb5jS1xNwR8jxaOb+YIxabEt/FuqPLmmjYwDNQZv6jfW1clmaapXlDmn/D49nvB0VrmfdthE
UpUM2kBEmMHYvA4BG+9m/6KKe6rDBBPBWLyZEtG93psAmZzvfLgxVBAdtl5D3sh9tZozA3A7DAcs
bbFcGAe37rBTU2ulQCf2AkM+bHdefKFMWvXlKcDuvA6qW24lrIn53lbVAT522P1itQeUmoGbqVd/
vtZKQkFp9be8xVSO+O6aKTqQh6zkkzZqzUM6y9W5tQwd+eiu+BW1GQt1SCPZeDfx3TiOuw1RICVy
+0Enj3t+xRkwFu6mosF8ZzeEKQSDwC8nDi5G7HmAfNfT0Zc5gnOlQTAJ156ti6sMQRIn4aTJYloD
F/w3yRkJvh3db3teZrCXMqQxWwWJnSe97yrFuHvF6wAGigbNhwiWpuNfeUn6itXZbOQn0RxbkIiK
cIJjPUQlCN2shXgUasxJ05A5XlXW/0kA4hzaX17PaCo0WIk7t1reCvXMlLOYTpzCjL7MPhtKHgyE
Q39LiL4Iy2vP3523IUdsm4k/0FKfFL3oVbkOVegp+xCUFPMXjSdvf49+i5cJIEZneiJW2DyIX6P0
QmCPdA+dtt9Ti8rbX4i87Z29HyMqYrQvM6KNrB3g0JNIeihOqpGp9FWkUsd2WzNU7hHcc48sxNXj
2zpeAGjEe4zyhkvIYTmlULNeN2XJIR2W0XIcfMpgi8lmLpA9v2QiZDQDBKoI09YrU2sPGfpqHSju
/il/XSOTiAj/kLXfAUrfyxWVN/gu1TSUldGEjLrXXuHTgFZt5x67Hx8SIlkWH1eE3bihmfrE97eB
+eQS74paeurOS64tjyH2NA4acEBT7O8Rj5XUXrDgNLClNNIyztfQq0W5sR+XzUmXK9D22scCCnz3
/HpAgjBkXUdApH6rJUZnYrTqxk/ThOHh8J5Fob/j9CJ4Qm7uETim+4wMsMm2yGjRU88EiYOMfyYM
dR4IFaECk4mDI2GXeOyxaRCW1+TX4vWSdfQHLn0Bj/kdP8zEcAa7PCwNgarXSkdwCnfzaCk83+r9
+E0vf7wfAp6nfZvhR6TzHeA5J0eRAIVkPqcM4TPtbIikrpNGPVm8J8Y4GOUzCikuVPO8i7xmY5Yc
5n2bzhkpIQ1vgC1NsDIdhfhLgu1FqrNwbOVAmJbmFUCStITN+qz5DyfH43n0b0pcrP50bSPUt91E
vhPW3VwCc3GrFd0kOF0iU/2vPnUCsYr+P0cPGbOKe1yFiNHs0RrKY7aKz0kWeZf9wFZ9L3CCEmIa
IEtgDL+NJh/lDHIWhrWSJaRe1Cgusti8Nkopt7HvMfWXisVkpxwbftgtgGfwdmRer0McEQa9qz7d
pJOtQcdCrErYuh0UuWLrmuNd+Tr4bfX7HkkXmVmNyXqjXrfdlSmb13nfl8R4XLzeCF/+4lwqorDw
5EX8Rw2dtGcLdh+0JtW8qSQUL+W8xc5iExUqjIKZVgJBust8A/iC1RcZiEBFRxqtkqiB5UcA6kYh
JY83wcV2a2hRMNG1MPM1CkqG591G4RrT2YV7L0Kk0nP+O+ePdgBpPT7VrEkKlqBvjX9c3dksoBxR
eBo5LaNiV59neOuF3yzKlV9nshFrhg21G8nbz1UXqS6/MdXaQtppf24vjICleuxgmdo7JUw1BGpf
DIWFUctZ2xmd1vPNMVNULjCzJFPXNn7riL6qS5RjRM4DXSi+ppRCXEuomgDdTpOqiwVEljWo/ENg
tExg4sb/VcVBXlMRGAYtUQItCCnrNioefiw5INjSRqtECxc5UD2x5cWrzPZIZi1ev33VWdSlU3ID
i0PxaVJ7dAhvTEchxJ+1mmFUAslpb1fJkNOE2FwFb8JMdoa2sJ9Z0Ti8cKieZlbIS2hBS0IQrzTL
WRUR53bx2WdSzQ3ZqzPnaSFUtNZZb3n5IW0eyy+eOUIltkZ1c6rK//xLkPlfPGo6L1LBsJyI/K1v
kBPiewytf6QH6WIIRFb+8nkoI8w3T7XSTQPlPnPmeXTfh+9kPj8nbg+3pUeVbrF0BO6nieBTdFZu
kTXAzRCs1k8gIIugRToClwGShXYMdIcVxuqLyV6rrVQaCyK70topjkOBtccmqbIcZbO0iQu4PfS0
W9Zt/LkfRoGYJY4QyHSxGJT9S0VXy8RQnHI+rzZjuZFsdyrt07s+kubH7J+6s7L3iKY3ykOw9pfl
w4oFwQqcXq0Eu+yyc7wl5BSasjNs80gSvRfbKGkv82KDh2BZF+gU7LBdJBRseEZp6mMyx0tsOz6m
ta1EFatDkTE2jqER6/50LO9i+6fbuUYUMm636AzXT6NZCBiKcicU8gxlx77bsAb+kWj1Xcm6yOrB
WSSKQyEbh8DUCpHCWKALSc0cXhgQiEyXz2reV+y9/I056qiastreJYBwZ/Mug9eb8+SyLG8tSYYX
UEE8+QvfWubs93PXVxdGbTRFIclFGWTzM0B0w8rYtBSVo8TE+K9v01wkk5zAjYUTC4XywZw/ge0u
OOD+zDvPsi0olgSif+Kd0ihyjtmkmJLMTvaRTLWave2Pyw5C93HNM4t11nzE0M1G56GcDwEd6lWK
yzqDk1vAzjCEZBAJ00esKq3bs7M/xMzTRtguIVyA98c4jBsGyTA83XJ0lWDT7/YPNTQk2W0D2jEV
dpMS5eXgshxo8EGS7sYO+Ayh/Ucet5a+mO3bLSCGOeYSMDztRKD82b8I6ls1LsZCO/ovQsIq3oD7
HN3nFScqqkYWf/5fShqVcbjUlp0hTn+H8S8XHhvHf5pCrE8CX4qyYP7hiDdYWeoataKAQ7M53ig+
syLUaMnwn7ZWEnH0EA1b/DpKkmZy779Hdhm+dOSFG467uxL6OilVRCT+COadCWB7PcJp3k9l7rAq
xOxgmHGV3I3KawvjCH+CBRtdrh4ZH/Vc2WUjbhVXSx7uTR5MptupjlW0T0J0NxPf41TmX+NpwCfO
XrGHgGslTeuS9oQW9k7wSSRZVX6DIBqckGzVxWAG8wIzBBluXBaqCxbdfvojgJlndy1j2Wp1zCh3
QpnidFfCLN+Ovsla3Tsq/1XBmI/XUKjXmVnvucgxXIrSOgGHjxAuarhMwaiU1W2exG5pZrwNKomY
w1U7/6plD7Xzm76OLJQ7+fy/gi6ZL/wU2mqD201yaNw1sR66X+IueMnYofEMGxH2p0kQ8AYK7dg9
OU11nX0JjTlDpG68gurZqAxFcU7iMafoeIglosxJeITnsa304cfU9fUbuNN4KPfiZVCI0FDh8keD
zaeK8HI4eiPOY6ywpuJMOkOw5JK+I/Krwpsottd+IGekRV0kHlysn5ZQeEj552+V9XGrFIBT1Qut
T4FQtBoZMCh1QtdkDCW+MIM9VXXbmPPsUlxlwhSh3g0Nmnu0okU+QvmDcDFM+xurk1wEWCNINQBI
D436siHfOnvt2xkUiR37zFrMADU6WQ2KTc5fvkRKdKjsWszCuPbLIoDF99McpYipYguzGZgbqyns
TwhXgS3nRJ8qDyNvD0C/0csMDWtVTEU/62j06fdAxGki3H35+y4VVA6PEIRPgmcDmqaqpAXdjULn
gpEDozCs+ttekWfPLuT3DnCa+bltFwq5xVKFKI+UudMTA+/TLkzIE4u8v6f1/DpCq4E3ldadunXl
j5roG4nMgg5H++9FasmiVpe+/hYo8KprKPt/rzDGCITQiKIU3WNBoexLUFSlbzVtLtDIjwWomHWm
uUAes/9CM8xptGWUUS+mEKD8G2dh1xyfQL/xGjuxGVwXVyz18+pFfCNZ2c9FBiO9oQP8Yre67yK9
27HiEiepKqR3P99plgmoulW70wRWzfvkIG63Z15Ydcq95x/T8unq8JWBnFhyXW3LF+aTAy9y5UGy
BgcZR5drXFhpuDh+GlV0ONEeJYDzlDH+/UUp6frjrWAWBWnHgLgMWXr9k3PnjY74MRnUvIOEjEIu
1/V82//6TeCXbimOCoZNtZUhn1iE8jZOOvBi/OtXrcNzFQYda9RkjqSMEuAvbggKgXhjp1iTKyys
zYtnQrFsYsL3aNrwdNYlHDqFx9btvjsARzuSmnMZ5ejaAPy/ih7M2PISprZrqPTAsEvNKWc0VXo8
PsWTNo2F0bJg+UVq67fUcc0pTtHhyZBQ/9XpncIzsbILg4wwtR2NPl/wnnYBSQXKg0VSBktnIjZM
dy21BZ3ndvSMsyOt5IsMLs7mhS+miTYb0aRhmLIO9mdHFZfG4/i3YvblENSf5lgVVNkjk5JlewCc
TBnPQdvZeRa3nTJWrwakx1QnEBod6wFCw3/4ZQdEqb/e6DWDvahXzkW8vVX+ks58cHiEQcZ8o4+6
QB3wpPOWat8UeRvUqvIAzub3U+MqrYHaD5Wm82Dw7NdCxlKnhvKPAy/6G137nOoibFHA51pm19uI
nxAMAKeKKtHn4RjvVaOzNgoslN/Gdjx0n3qe2r4gtkGjlPH/8EJwuX8HSh8epetddWQsQRNb0egK
7luHE16CZyK983cJdZSIGBbGGnU0VphyRhH5p3hkCN87abo0AIP7XqYQt3O3qnmOUqT03t4ICGdy
2na180zPcRoX1QlgM5ScRqLSV4MloDkUG6XYhKJtIaDNokktEnU60HsjGefW9jFhCx25DBj6wHJw
lYe4dJQzsub/tHa4SBFUGiHOVLaVV7U+iINGcDWJewEzCqTbl0fyliQNdm2mE3YknWHILYtzirg4
JPolD+ZX4ozoaXSdgpK97k4F1DHmgZwIDj3Fo+Sk5+e2gjMbnXPe6HjfEM8vS/dDvFsTU8Rpc1PU
GKoJCfX4A/cZV2GswBhT7FW7fj4RrIliw2QA6rMsSNDKeK/o4hqdHFlNUdrUblj48gJ2AqHT4olF
V53tLqplU8Y0Pr8I0loeMuOFRdvnN6dizAk4SrzECiMDrIjysHrXt2W9wVwMV+gY4xdM+bWE6YWQ
0MWwjhJKLR+2iAP7/FYYJein72vc3F+zZwsyc6d3jdlHC8qfBN9Ld64X0v1xDaRi0/11a3x9m5G0
MkHohkoQbvi2FCOyDaFPsGYmoGE/3872DB/mOSJMBc48Lv7Y1Mo7BWz3t/oYKVxeDMX9WQMxhBFQ
V2ExO5TYN4vSREvH0+QpIQsIaxqbD+E3HsxcNAxOY0X7rJQqt4LIyKDshSPnbZ9o8Cdez17hNoCm
+3X+bzDwFErpTzduvg8dv+oaqxU4J9QZDM/RERCT2Nig0FDpqOgqpHwq65kNR9T6Qmohb4Cv+Yi7
WvlauKPespGgB8fIQhv8PSIQJMpXD8a3G76zQn4QC6L7XPdGi8YzgPd7vOBEKmXiH0v/M8L+ajmD
tMvmyMRKrfRzRlbOEXRejG23hNzt0jtJZvjIATHltGWnKRHAiEnZ4D2zeKrTE/FPKW2tbk9/tgVy
gE95ML3WQFv2ifi05ZP5kat+Y467EzVeGLcKO5r5BfXOPdVGzUBbDAEDNeIEmR7u4VMiz+6Em+I/
+bZA4dlN5MIGEENBafYis+oOxLcdByW0YnYaBkq87SIUf6HFEhXvfffsueC+jlJIKI4ZV4fCgBi0
+6gHbkgPIBTX44mLnU7oSGQizpl4nZxSc+fOCRomoJd3JZCA/Q9sf3XwTjGPCDH2EKEwuEQ3apDW
3RezDtQMK+kncijg1BhIyoa3KXuf5jEbPFuewPtlZoj5Nmjj2jlBCcu+NzBkwWUq1/19rwgERgXo
77GHx5cam/p16ZxDwiUvCP+IK8HUDVcqIhIaGWlTHpxnjwGV4l0K9ho5kpLahEtojqfAxdkeN4JJ
IPRqq0idJHo5eKMsIB3ixFdu5M2iNtWcYMl9CRIto48Iarapz85k6SWyu/vUYGxLDdTsopT+E7WU
tvPX2/HMZ+WpFxVHIOmGAAj5gQ1UZBb4FGTLiO0CeXGBkIhCVo0OfNeHTjoLgYu+xtRdYLLlNQB4
lvVdPQAMzeCksBc0Emu1OSedgsqoVXGRNdv9ARxKWhAo+Qom7rVEgQhGfHjTq7MS/TWg4dJgYtsP
aJuGWqig3BZBDZMhhiC2jR6BJehXEb1sHivdKphCUaGvKw5oMM16y5TuqXJVnDGQYDPRUuObP8as
HsrjVFzYe4gkfSgqulgpqqqW1kt0xOP821NBN4af5qjYann48nNvMdcKJb4WkOYvQz41yW83DNVp
dbV3NX0yCPByhIy/lrTGg4dsmBfsS6SmQLbeRT2+oWysSqeOCGBC6riJgdYVLtjNymbAJ3i4864q
94FKvUL0hK8pVR6vkOQJIe7idJcaPRc17jcOenUj8DJPCVHNW3ZyW5T6JCfdmHdkAiOk6O3HhYWu
Th2mtFVmZ1bRx+dhrS4Q23qaVd4sh2HkqWD6jXyKo176pwOdsOyWYRzRL64XeBowmcsfTPhLssD4
4Cw54oxru8hVznwxlPAMap1l2slb6N3YUkOPjDPXI2uCTgOlVQm0W2xIWMoBgP6b7ZqhTPD1nr0u
sHJ1pgZVsKPSFb6EtIAE6/HK6T86sGVSFVkd+4r3h3uhfn6OuOjz1gzgTQMQi45+dxtqBXaYXHVK
pm+IriRQj44eUP/bXf0mWZJFIPzK5h/q7EX2CJQ2Tc/r2VxNwhN9kHfHGCE8wKfrbYxlaAU6H2eQ
jQidgCfBpIGJ3dhw6jfd7PphwlMMHEeW3cYWak8Zh4vfxO7ZD0BCmEsLEXW8ZiRk5V4GlEEEYQmh
Z/2JpRQalKC0Uqa7MPpxL6KBK5W4x2fn2CIay48crdXB4+WXcKC6J6f8HNSHgtd+8rjL9zN2r7eM
d7C+cEr93C3886JSGSbWA93A28G3Bl0BRUo5M0LSu5GvnVyy3lhL6T7upKDi4dx9z3g6dQFfP1gR
K/DrsNPatOvIA0r9j+HLd01MrSx11A2M/XKhdqqvdcv7orgtMNUaTNkxHKB5Z1yDTF7OP2BRdDZL
cwAw4lfNJbSAAzmQdCWPOZdzLP3OhsLzCvYJ3gRBFrWiqyeY48q7vVEueIFSYfVbsGbvtd3olNE8
EQpjV0BULt5yiozjLRUITNBMP2mk8+pTU3gR7TSwXUA1JmQfLbt1+PL+n43qXFyrmevjyio+dl5X
+G5fDt7sJmLLtZeCjgFPABsVtEdPs+CJOmfWwu49J6skUmyGCnAqxP3PWCOBfhwF8i0P09p0EYxn
mlQNwc+lUNhe5auvN7wEtLq/SydFNOzDgMXl86rPppQjCxCIsDm/MiBYNcqE2/PDsnTfE3lBDsqA
LEVY6Kcr/1Dxj576pgErdwC9y6st4Vw9DJaII4nZ/ZpxtO80MK/sHNIBRc4e/Albu/6f5um86x7K
0ESow8TcY6kXxMMR0usLZ9h8TBB0ffdNpcy1CkU89dLPD+WUScbjjE2C5817tBrzdxE2d1DzMKmq
t7wnYG33yS6Yo+eBTAUtXYAcGEHMRpBiZ+LUdbMJoxY2k65+STL2b4rL0XTpiZAMj6CD6BcBQmdk
WTWKYNu9eEE4HzNmVd1Is53Lhydu9HR0x/JCbyBq82WoGKQK95Iqakt/CmouJHQDKwyOVKa/YoHy
vL9ZClntdsTa/41dLuBNCAV8+i1U/Kj5COEu3kaj+fjM/OmUu7/ZfBImQGgCX+lqJoRnMY2TfWIu
FkXYenFkiJMfVU4QXv3RgUI3zM+l1HdxmfwZ3Cbfjpwa9cw4wDsjHK7XceK4sKrJjdVk42XODQTZ
B3dhMaVPpHHhDV8SBFSIGlcamBVfzFh+Rppjqolxodu4HJK9obUAePYRLgVGAqJn8kqtSJckxgIs
CV9AjHrWofpkl4ULQYKzof2aG/xlTGwjL4ek7ymoq1J/8jzxWyP6HHWZcxc0zC84TRNmvRXcg+in
qAvI8+WAXeEFR1FWnEnj8clr6mgypvXmrDIDAykTSjFwhfeFEACuaHqzX9uKeHVBPICJBlXx++6o
rr158QMrToPSV4juvewQKreRJovBbprogpamwBsV3QduOiJ7i+9S9sYT9syAYOdsSr0GnVPx8VMI
Fizl8kAJ7yu8hWYoLypBPchBY6FiYP707SPi0Vk/exuQWJCse0o/CFHfm5NLU+rHjnzvzMlz0wy7
Baz9+QcBBztwjS9dcVW7/gTr2GzHvV/voccsaLnkDRIpnwGywRHYMEBFXJFmQqv+wenLmGFGxaAw
ZSAFIMskOlPF3stKV5w0skGkMBCXwgBsWP1ixK9JiXsqzaJrzagxn+aqHoaUOV/dFBHLeI3Xo+vr
A9GUitvCXTaQPXq65b0b0Z5Y5eEV+4z+oXxAks3rni2Ts0Fzo8okuyV5FzHJEuSoXt5DFRh/oWsI
GMU1A0OYtfDSva574Ri0CfP91xkOPbWlKzJ0c2724OvUq6FO+YjyD4qK6IPwD8FGNw/xWhZpKmmL
Geg4rZ3GT8D5OorzagqYhxuHjrN/72njAGhmkXe9Jj+/X5jJxNvYuRvwqq9hEbIbQNIWizzAgBFx
SPBbHi8OBIEvBHB12dtMYH0yar2fugPl7nHc9Z+R02MryZ6EmGQJjLzEs1XIDJJCoRyoiXA2+Jv8
5wZYKPqa4dWXn9AeyXEnTertSjz2dPptl3lVBmuVvK4Sa6ILPLXBmtCjlO/tqbTxMKNbAYTL5TrJ
ksg5SuX0n/NusCbs8EAJCK8g/ZrOdD+cJGRh+U1ukJckmXIsyRyNbiLbUimhYCym/fWNSq55V/y2
k+TO8KjMJlKcBOhogOkS9URgahfh2p0Zg82Zpvt1SvLX3iU5JmZSHlMW5WTdKZVFAaKQPtmG02R/
94CUK6KZ5v4j4+4lxMUYIrpH7nEkPZBDJoFsz5Ya7PM6TdI/K0kl1SaD5RbNMYLnKlxudtc4Lz3U
ioVW7W1OcQ/I8mdoOZtpm+aVRrDVWxb10vP2Zm1a5YvtJFxaV3BuwIw3BwgX6ylMBMYUV6R5DDo2
MZbz6ppg2b/PceSyd7P7dMAT7B1aNhkw0q6310RE9jbJYpjCphXUe72VyibBQBwUy82G1baCK3xZ
efOkYGWkwEfVFxSuIzXAVD9nzRSJ7huGLBTXhLthnKHk3MwupPLvOtOJFL3wUEbqu3JIoFLVIM0N
7DfJZwlM6/lu435HBX7We4OHzTvU+zGZhu35VxRm//URKKFGmwaow3ImVXOS7XAEJ7mFPKOvxuAP
jfdgNq5aZ7vFAzpIWvypT71TORYXMvUKPK8whyM3Z5kzlgI5IXTcO5gRZe7nY9Qqrd1Aa/fokLYy
tDYS8aRFEMHcvBPw7ATBcEtWnVUTNhkNPQG/AmARFtWJujSrPsgPK4gILho4XahiFZgubB3QhHI9
7OPKZ7IZWqN4Q5L75zFB021l+pNl3JdeZ7pR2ddjJwN2CbmvSarO2MBddv+3lHYhVHlNJ35vhKem
AWRtqAG34yKXBJdJgfPUkAvdQc5hvM6ttFcqNCjggHSxRf2J74LV8BYgebT5IA4rngbpsO9Gy+lX
EwusWdlHkJErbxl2YXWQ/aWhzQfksL0Qgp2f76uxkD+BhS8SxlSaK15qZqvoKg0e3RSW4mMxTgTm
QGT1NhLdYksiYaaOO0Od1lDd/hD1Z+ALtbrpQVC9tGtmoEXsPK3A58+bVyqURBYP7muTYZVLUJii
t7/8OUNkVXpYK09lutDOg7UnNNfZTMXdulfwa1QFKUGr5jGFysl+E6IuhZk5oJ8yEiF5xWU6gDpA
hpY+LqwADTkjmUzxGn8cnd+ZcwGIjLWz2WrZh9qD9POw5g0TbtCV1aeIoNLUx/tZQSb68RyZYdsG
C7VWFjT+TLI4Cc5XDGJLEp2g3+Kbc/r++XENQyvX8nBdRZEThfgub2uZuIYE2Iq9QrrYu2OzXUAo
TPEBwQrrBx/ad9iL28VsmfWKQ07seEagJs34Pxjxlt7ojj6oeOoYHoMn6gWtigo/5LpdxjJkgZ1r
jgyeLeVSw5uDBJeArFdPC4kxaDbf8v6BANEHk2iUCKtiOfVmEo2fgs7+CF5BR1WxOkGA4FS/Kdz0
GT8y8p6RMFcPjzD/I//6H3J/LL1IkcCOwLgSk+qob4J4PZxMKUXWMMGPHcNFZvXjNIAoVlvdbOqk
sbf2t0XZx3n02Vn+LCMBe0exL0/tucTHxt3WkX+r3MHDDpzV1g7z6V3S+PzlwppfkNBytvcNji1B
YVZeZf4qObMuBpUUVXxrXR6K2y6+TtWGa+qxB+t0UXFOPao9GgMdC8oIRaDygLwcbawh/W6CVcRc
WsJauZW5FRcdARa4OFoDUR7kVVaGtOFMhtXbQqukt4g+hnDxtQwvvwSmNI74p33wSnqodxLud35E
jCBPX5TtON2SLywIw9iec2T6E1Q5wjZOafu+pVOS11mSoMZVYCJelp+WGvv5hNCH7U7PMELGSPlD
ZaKqOyb1SM73A434uO2GaIcRQfzfeHaG7p/UN1J9SzZD7KRYWt0SIrp5ykwmcLEic1xyxWbL/KfZ
sUdyGSA7JkSRrrh5rvMo7n1kxjGd8ngyjgiuQXo8ZSGJncDfe5xkchXGKmIQYOS0lRnWCeOwpWwJ
IHEmzalZfzxIwmDTWCP3Fovtu3kUrw02rn2tsHmfZm1WT4O6TDrbHT8DtadxtfkriDb0GSxLFcqo
kA2Q7KRJOeO9Ep3tiPmC/NelAzzGcJaX0ULaIf2WbZVut/u8umRxCkvBVL/RP3LRaFVcNcohdUiU
f46hQeJioOTwBfohThd8JqqNlpFY4EyJkpVt1El8A8ASB+BAaI3dIDi8iVqhjgSvbGiHayj6i7JU
Qd4a03hGo8Ru2SUcK5zSvXO0LUn9o3rE0kNt+CDhDlVK/6vl1qJPDgpLNYWo5Ik5q3kuLKA420Yh
7p5R30kx+YGc4teIIEAzaFo4w1v49Hl5RBRP4iKBtcMRC3DvMFFLgbty7z1eBS0jexS+QtDh6VCO
oAP1S6qm8iesOxKv+4/yzDzcIuKWKESeI1Ekj5JU/Zndqy6MGCrYA1Em0w2x/6UKhnPW3PLR8/+u
VhKRXAqpDFogHA3hmB0e8U47oMwzUONzRL/VgqA4pzNbylPSYuHV9fYEMacim0vzUOAE5IAYmM+u
ONgh6nDkWHieD5a6UMKMnvOmgLfZCWjLAfRakMM2H3uwivFgjbHWtAeN3NdsfB7P0COK3mxIHn8I
SqSMk9d6TphJQM63uSu5qnkzdhftyB3Er9hSltlNJXWHV150wwAC7BSzPX1Vpohzta8C0Lam9Ysy
GNDJpz9oE6/aupjM6W6/0/WM3wkt87Cc38Xnb2AVm1CD24Zp+s7CCqh2Auzxwc/qVL3gefciTpNn
23QuTWoCJ0r+3hNWtgaBaBF1q+bswPbNOt++kOJPZvdv/MQpGv8Oc0EDXV577XZiWJ6mQNjLlGu5
JvPrlXUbZSrjfXGrigsbCbkx5TWiRea0eHRv66UfEMZ8+N3Y51Yxp+YXoNadklm+1AoEgkric0bg
S7gDonkv6kiGHu8cULTPilMl9lNo67J80C3qOZpWXP0vKhpIktvmaCzkx01nsVpKuqbTiDRPGaGd
w0nMQ8U0W0Ainyi+K6SoYLCz0BX6nr47q9atZarPiBnmyWWp2N8Ptlz9jmsh1YEoJdpPZVNLPyRx
cfDukCE0Ec4m2gN8IDzJ6TyyPjRYXfBURlgk+2WYX+3CMbv0ajQ3h/Xi9AqGJg4dDUIvXFwQxXua
Ve97lNSbJ6OknNCpPD/oTsRUXkxiGahv3LMYN61SkylJckZhPkh7iarVz64FYGfDkAMaJ2yNDuV9
v3ferA2Vf4O5yJp7jOhAEhMbbqi0xuRStmkz91LJMYw9a8ySMGV7RUtpMtpJPS6FVBZGDmerjr63
RodGZIcEz7bQmxsHIid6GaPHohkJH4gCKhaVx/BnvaGGWKYAVLHT2NWXmP/uRhyp+khuGN0tbm7Q
+oiz8DBmugvDZTQois8lOAeiPqSSfdqsqFpfNzODnegjZj9+2k1uvj7UHam2OCWDZGz0srOVQrhp
d5+2Gyxz0afsj6N+0aXSik36d5lCNJ3HJlUhqWdLxPkd5v/kyy3xpoPyScSDCC3qUAlqbTXk97iC
f2lhXzjjYpp/NU/4eD+mJ+Khfbk0w7OgpY75WaWY0eGjVUaBwfIiPK8gAemof9U7IzZ56wDJkQhy
4kgyUQ6UbHK1SkWiFlYxf0uQ+3uB//gl4qVcQTW3tOFn4TeE2wAqXJ5QJdr4O40KRsSxVwna+S29
jXd7QTrbigtlu/YrRdxeOAPIHsqrs31UsxHtWvV0mu5jn+JqLMR9x/iV8afJA5jWGFZe62TQmjiB
UzVspixjbtu3pTTQdTz97xQEQWET5keI53X7VXQMAt2sYKyQohoFHVx5ixVaEwg0sZGN+gLq3EDQ
yzXqwCDvHNPVLB5cJdcL1oEnHkeQiLU6aaFQaAjuy+388iA0wMlOvoK/2Wx6ctDJmL0zGYB3vJPb
PcagoNVehKQbhObuBPTMFcmfTsPGXzovkvj259F1+6NtEVNjwtM09c9k3ElQhDLyXliTBgkMcfX/
b2C5RBbczQ801+49EMKL5E2V1XY1w8qCFNziPzw4b8ccFpMB3SH2wlcQbFbSTd2Ibztv+C+MY7o8
iiH51qXmon3k1Oto7gsaXZT/ui/w4RdRKK359Ar8A3OkiDrTNZ4R+hAbaDWGccDb7TNv/od/217N
kNKBkKrJi5G1l+N2IGyls20YP0wdb9nHHDSvH4Tz71euhU31dtF7beh8rXf7fAX4EouaFBVOrWdx
9WbkgbLTfT/DWWIswrvW4sOkJvVzqh5Ujkio/0w4AuruenLfIV/ngyOce+L7ONTNXBNNcvx503uN
k7qaWCkanDxkrj+/O6qGWD8eDSyHubW2Pz8RvaW4YMcuEEsk46w/pDK+1M6ZX56g5Xgu1t7a1tAI
5Y4qIBB00Rm+94SGHOKHr6Z67g1pOxgkIFpWzxchl3Iol/KyRCqPlNhYS8bHpbVVI7aqP6u8NSe/
6xS8hFfslPrffhQOl1wXxIzSjg7dUXTK5RITR4sleGNnX8jgARcBaIigcbPaT7/L03OF6KJ5+2yf
5ytgopcbFfPA8NZAoGNfqkxLtCfZl9Cwyk8fhuHmZdSvOWBhm0sz8ktQUSTtQ0Snb0fFUTUWmWeI
/0jkBA5Y47gmPm+7q2XzDTJFxZ9U4AhVgWH7zqOSt6omif0OIewQtMz7rEhDX+CJG8P2TEn4rm2b
u/8ZvL5ZTvyMUZlcFTdbzE22qMJacLEfrh3OOkpKYlqZBXX+QeFiveP59UdS8j8fdeiulCios09r
KaJ+P7pcLVZRD48QbfHlP4zrsLdNs74sJX9SQyn5XY6rInzX4yYAxROw0GPbPw4wJ6pNUTDtgKKa
DTefubV24ZoYan+7Ky/5H+8vf52Dgf68cq0heEzyRFM2dnUq3h1xBHhvFWEn+In+xqYhyxkYe09f
mVmXRqN1fda77U1PN7Fwx5azBbKaq1cNF582aLbCvM7IMrU6FqlrTlcSwnzwOc8X6ro37R9SEwq2
XaT+vU5PFPeAuUggt7D3eISl2uiAwwQzwB63JLdfWrfUzUscWkZ57IG/hqOhwIHUZCO3ljQOV6zU
krtzuyRpmsmsYabPLa50pSFOrWo3N8rBHOWLIsv+rYRIdvtBzSoKwAlupmgfLUf0jiJYclOHI5Kx
TDaMZCzWiOME8aBV5W2XzWBKwoC6G2W9DaZr49Tfe7LX71v2VCIv3VGo8j29bpsDwMG65A0ZJ34V
Nsdkip3gTnV1e4m7LJteT6pYN4oKFOF6bgCsw26V/wYGcI6Ul2diAkqpSTd/AojZZU1/DtZ2hBb6
ie7OV0Z6Gtlq6424ifyJuiFSQn0b0TFLb/rLbPEsOra92lVPPjT//OQuSPQkTmC77NUYR4Ae/cDB
4yaLzVJWKLApuOyFzuY8GZLnOim126hagy4hQLepe1Ovi5Z6w4OJLAP6vZicqrCFDw8u0wXCwP9z
rSkH49TZnA6x3rfCTcxnM3grHhV61nQ2i9Y3kKq3LVZExVZbb+hcEPiN5FHbVWmvtSQalmyLO3wN
4NeQIuGDWqtlFaCb1Ehd/gHkXEUlZmb22sEwQcg+TNfjXJvs6bpBuB+ouJEeM6jS1AHaJx0sakE5
kXUPVng0YmrWnFwnKwok7iAHOAPsU83nTIwSLy1zUHBrT6Lhsn/l1WclwX2LMbaSJK7hkp0eZiXd
HiLEskM4RtiCGvBNe/r6pxVDsRR8MZyW3uNJd3I6I7JRjrffCuS9uYRhZ4cq7vjVy1U2pRsIbaW9
q1NS/034biizXw0Rj36OcjqYWeZVcF562myTSVJ9+XmUoGGDMdsS9tICLGdbwMreAR+K4F3G/owz
XlMMlVs1f036uBvuva9/NEOYiD23OIXRegpw0jCgw4W7QOE/nLOQY9bPB5OT3UPas3J/ZjCco1tJ
suhyKWzx1G2zlJI+mMabkff+IS1N3bxQViyLOYQ8Bw4roSOCeA+XzCNDPVPkyvtHgbkmZZglJrw4
JVyHJB0QDuWNtHDYnA3W+2YjJXRH/7JGUbsEfHsUbi7MKbPWWY8km8ecNaxrXxy/LqkZe59u9w5n
E9n2WMI4AhKw8Ie7CZrYvsNdhsQxua8OzezGCH1ZkRvcIzEkGq3iTZ7Bxz8rcjfqT515hHqEstsD
kJT9YTIbf3shOtR166p6/0LravizU6Fui2blOMqY036yNSe3Pia0DQzSmhRkcRszZ5ATaDQRQv9b
nJ+ARoVLbKnI6ab1iTHKL8N2tk60ODPLyqUk8nBPHtMKyXYyJPUefaH9jnECDgocIx22XGP7tmF/
dDRHNl8ra4os01lOxpc7r4RDSqJRDvxGVKBpV8cBoBNmGmgEunmbetFJ7LsM6qWjKK4QzHRrnaSH
hbBEI0jmIVrOpkXO4dvgFG3y38HpsV8GZs5BoaLRl1//B1Nbn/HKKNAg/xhrFaqPwlZ/EbgcuAZ9
3De58gJ91n05Q0dzZIh//ByLYgn9yZAn8l6J7RGt2oMQw0VG5m47XHuAzv8iEg6hkETps2FLLlke
pIoRtNVTHTAO/s4GueQ9AI4ddX6oPuv7uZ4Tc3nkpQ/CuC1X+fbsJUObscwA16+4Rf9YJIfXa71y
emQKUhw9q2K20VatxGQfrBH+GbI0Me8A6Q+qMixq6Hv00muQ4wJtkF5snezLcqbh7GVQOvTKa2HG
x/Dgw34pfxAWKTpKLMcs/BzUfvNmfdtTWDDXE1ZXzSPPE9Ux0dupO22wqqH0V7r0trGrNFQrs+T8
DRDxvvt9F6SNJPN+Z4xYiORh53KLUCqK5ORtTfFQ6GaUb1ijwUy+GoazfXoDbSEX6cUDLC1L2I6c
ha0cQha7krukIvA3nlEKwEJhqhNx4zerk76jJOE/XeydPxqTwmLmDyJufcPTpWYU9190uKgay0od
lUmiqn1Fy8iOpxHG/EYDdtTv3PJfX2V8QN0louQSyudE2sbEJ1qEQypY9xQjVRfMUG+oaJLD9KV5
hkJR3KeYGVFsvax8aNTZmoSqNNixDYDI9ebHfKGU6DFgs4zcX+1Xh99SMoytVyeMH39vV1sTUD4i
5j7rd+sbDMdqigpsxAVBleEBaZeAgWGsuPr1db4DouPKXJjA7XGrC6B03EUHH3zeDP/0bPuDUtvv
gdQnpWG6hukj/ZFkv8VQxtAffbw0UZJatvEJuTkUuJaZGoCA0EJna+RP6Swtp/gSbecvbtXaReDE
1TmMV1NS3HINue/dbUYEUSxxU+bDPIZBx1snoOxtTuAIoafkbjzS7g/QUUN+pER/7l8Vv1t9GYcz
7N4MlJFMYsTQ9P9im/eApD5IpzITTrn8/6nBfA8vYTYQ6LFGzalJyweELHeYY8YyECQnGaueIpNK
RPDF7WG7VGYX8WMwPaE/gEzvEJ6hL2rnAe2W7W3bV8a8rZSxN1pcPGdiGYyZhSxR5oSni0+Zo/ZB
kOTv7Xgd8P9hcAfBY+XnJWMsHDD+2bW2r7rIaCwMNXP8S6rY5CZciWenlUNhqmDuL70XSD/P6oDx
m1wKdvFuhjSnwyH0SVyxDGALWPSgkhRCcsYyaTtkUxsf0sYwpoXoB6hJnmpwkfzDBjFeB3LaJcpt
4/X/uHakx4PJnYSX1yO2E1gu4fcqMvkyd21uO6loRO4rjLDgiJerLKQaHIm/wp8RC72bgjj2qfFV
Y18fJ2FbP5JHZAnC8UhKbPvFeTRnAMFpodwRZGovvoXEcP4k3afxdi6BrevDh/+xgsw/Oc9xp/54
pt/ZRWhzgaY2wi5RW3pGj2Ds8NZpsjXUy02YbaNS8Ax5cIqWtkudL1dGtz2vK9Vdb5unB2Vuw99f
fZYKhXlAO5aExHQxDbRyzku++Xc7Nf7hVxg/VV4zHNbljo08YfzD9pwKXeYePpzNDQRIB1KWsgQ2
mcCNj4o8a/p1OhMLx0qylErj9tGJjQHIq+BFyl3p0ib17fLF31aJzcUJbPWa9aGVCBi5nKGPqRjZ
FXM4/gdVPj3W/IpZU0gzsQeX8qSM/OFWvhMj1+rFKYPhnLUCUnIsgvN4py0MY6/cmKGWWCxbNYqC
6StBLnDF1WUunELIr6bQ1kJQyhfFxjjaXbESBmjcvsyLD7y+CoNVlvsV/uB4uzBYCL9Grtomx9PU
voag2y2Wo1pTlcFMtxdPwx16dTcsIY6rhBcmfLfMB3UwwPMF5CPQzAqrWkOGPxt+7k159s+70ace
ZqjaZ+K6DHj8pooG7Yv5QYH4zSBMuJ6m12ta/Zli5g/CEOzwQOLpS9k04Rp3o2+doaCKZtoCAfuy
hJXj4DBWNMztvmEgLoMWKoZf3buZqhPlTyaY2dVXF8OvKyknfKKACXc4CgYZ26xeypx1D9TQq7QC
UrnPyHPAwo3DwQXxmktbsZIGJhcupbIVDXvAhAfVP2zmQzUZ8IHW4ca38FAINT+i9ZH1tI1+CwLB
L01vYQXBjZST7XRR9n93/w71wwrphRsh3q69EfEXDwCHzvpTas3+qCzWx700cbdGP9Z6B5JhnZOO
piHWXzdHviRrMvqbEj22+5zdRc2LFwo/0XYNnpkHO/y/9vcJYRuN6lYoMywIfwxwVxB0NEwukGzs
DcoPVW+Nw5NFpW+2yppMznp0/iNF0KG3q/tAHTXriAeyJtLrxWL7p2+MmGJn7ps4DSA2sxMP5I+k
nM+zpdeKGIQ7Ygshu275cu01UOVc9vUQPQKCqgJ/fOFJD5vpfYRI5csdD5YDxGto3lo/vl/uqytj
ZKrYGZW9azuR0+nt58rYbBrr+8nd9F4OeSNeEOiKq36WGZ0XVq7O934I23lRnfjWrHPifmvysWI7
c95h9wvgWXJXMtmq/o5UXAbEOWOKZs5ovYG0cb4ybuSpx1vSjy7j7GaJatlI+JJl5+STbrKEqybW
Anh1kzYQAoQeml3DWipb5eeYmv6tSEyVkzi/3t6scREIuJnZqaOSW1z4VJmQMfQjbVrS5XKTgYU/
YpfLI9wAV7iG5MkiMzNQWdJZMK51p0eJD9kZB/A5yjQTELgTfY5opOgVPZ//TWBCyN8k/1Kv6HFN
IqR+/hA4x7J0mBbA6w2mLznzJSA+tfeilz3EPB8oZa31EAKTWgORi+rZ9iYIy9aomiziQb8nocCv
/sJqerYwdWl5rEzt3q1/Ii+RhOR+jOQpSGFJWC7exRRGkhO1WsLkCRdqkEGQSCq3z1b5NkLWPaXm
d8RIyQ6qDOeRqPxNlfDx5y1Sz8jHlS1QiQxX3TkzGJBQ4FCAVRR7dIlCT6wAG0haJd+CDnDBFPKE
l5TTY2p5zQXnjTVTkn/cw4ds66ZHi+rAnTQhflbxw89Os2IMSy/RxfPvnnjStkH061YMt1x/QgEb
ryKm4PKXKwNx8DnY0cr9OqEmUFpXoiqFB72P56TTacDrhwzGiAhaSRuqsETeFFgyWkLh5DsawAM/
HV+B4BTuXf/pmHC+AqxjSjYCGTFLbv/PJz6s1WARTGDt8yhJPA6Nn9y7OkqVEq8f/3nsyas0fYfl
40m/3J6kzddn9CoojwNvoWPh05FbtknXiGLDDTjak3hMPmpATZ9R9McdBEJlfe/2uaLdyqWKARDL
+T9v8bw7n6tTLAP7gGc8mE86zoG0PUY7OhdTgjHcoXOuXikMs3301VkJVDnebZimCROa3AjHOape
JUuCwvmJkXIhKob+xzsWK0Wo86dXAqCY0jFV4zhJ9f/2zZ7QxPHsQIoBGYoQ0solmaVI8vxueNIy
7ymWrGHi6oXgqmNOEWo6pyIEVEtmk3Z4mVjl27Ut1yUxj4yxvkYeKawcVpDzgp3wjmS52Bl/YvWx
f21RJDaqRAFiDRSs+9iw2KWDW9CedRgOz1yoPHD+uf9WelCQP7TRgkl8tOHbxD4rxG4xcw4T3NFi
CWIgOtAX8nj8DXeHz3BMziECegeb3rxFI7N/AkQiSc4sWRN3f2p7tNv/PBTmMhzh3k3bp5dUDN7r
bLtfEpgv2yWgVbWuP7wHnCHSLpl49ulH6kc9iA14pPgJH3F9ZST7TDCbE7Np08eOu8vzBqh7/yOV
Wcw/Vn81N/AlBUEj3VCICJBS+GwEIqlrvHsAn5dOH+iY9tU+HlOW9lVl6GPxMltA6zy6pgjawPlS
VVoYig1pT122Zg23uB2PrBcKXDcJLvc1QNh8VA9hkLsnDx5//4JzC3RFBllvUFoyv8aEbJE+ufGB
eg8WutVX+fJkPRCyqtBPm9CCHVorQMArFDw0Ry/7iEWI0s70yuNZFNO77vAHKhEYQABNznl0s3Wy
A3DfVZf7Am0C2QlhKufgY7FTMBb2pn0/F9/lnggcarFhe2z6U3ft2k7ODSqseYx/eCfiCEYP1CEO
E7TS9fwFjC0XnPVgnX3QafT6E3kXuOy3drudGzuFk8OB1T5f7gWs4ZLdCydG2x+Ac/DbFtvPxBa4
qMPz1CBHZpTTb0n2KFLh7+JefUQWAIxZQHWoI4yKLIHJVLztprnOQ3khJYoS6YvOzDl7QeDHVTTg
FhKp6OfLj/It0WgVDEfQfxXBaE48PwEsmpQiae+ihnUCAGVnMd3YsjGxNVc4iFuXEg5O0P+DnwbH
PnMQDDvmHYJTTmUxffZTcsQ8SOyrATi2KfqNnKhHAF8VmDWYo3AZ+gPRx1QK6Aw1Sdjtlrdg0XNm
xIY1/3v3uTAypPk+FvKLZyGh7r+nO3ZgYxIxMTk6Ser3+J6+7K3HYlWnK19FNaWDIHtEeGWzExgr
ngwyJG5CgzzUsGp4Xa0tVW0Nj3NOOim4peTM6E3IdLYOTv/Pg47BezFM++zhJR1yklBwt25iLd9H
/qsN4uURcmjACmCuJOj0OJQ8YGKdNeGTRgPyZr/0T0fVdlSQ7XYa051WfU5qhDylWh31JI2zq9hX
PyVKS6DsuD3rgVEx5aZEw5JNyw0Hxsit8AogVQGUcG6z5AjEhz076XiqasZvp5HACl41rJWL00ny
5445d6ojIK/bydOfF+73CfkDVda61qCeY2/5JslAb25R3ktrJ6Rvm/wgLHKP+r9n5+h4O4lWG1J0
dMgeFtHLEVcbL/XSXw/nrQLvyZrAAZ6Z5POEMSxpvUntbrNfhqEu+Bvd6xcEqCIdgGk6Wz+4oGYP
S/CnkLYqmV/Me1csX+7yu75EeQ/XObYHjKDZ67rHITYby0VDZBdH5t/M2tkCGymZXUuj5b/YudOO
c4fbCMK7uN6zbWRSi4LeM8I9mAC4k6gjgKqiaxf5+QVAqX4ULsa/iNgu3ucW9dPpXHZ2tYr2s0Ig
FoAQ5txi03qKu0lJvzUiKr4T0lpgAC62GHaPpelfgdO0RNDDzkm1Jf/LkSJnSfI1JFLl60XNJscb
xK9X+XKT0UsSn+X6w8/V05cOo/lGkdVr2j916N2JpFkr7r4hByVv9H44LnfADK6k97mkM3Sf1k4v
bdm3u3dA7M9f7cB0mRw+tkkFgUo1ka8X2R+HtlaicV9YhJS7M8EkMEhFIUsHDfvIDbkRQECSXk9R
5p1hw1MuOl10TolcRnzrOdkVQ8oQRGxqfO7iF9T5Y0HQVO762CIhkPhJj4U0lTofmIOY5jSvFgAl
xtICYtlIJf0HDrlErRzrEdSJ9TpV+wE1qVLcZgVSRkgVRX1nWEZufOzGIn9tXAiLzB44UAM2HoKJ
Pmnkh6o9UIydT+QbuGYlaVrH9P7rpUBuGGdqilP8A5XM9dJh1/xGZOD9tLCMZFbLIAG6mqbTbrd5
No0CaCbeYtytSyP5fejg4aFsuO2sUICrYYbMi3yro9GRAcYjHhhOP4vPxqK3FmVdB0vgsyn3L8GY
L8deOiYTWl8Gx5uN9PqngXA/FizkqvowIAdxyYfFptTYOEc+ItYZoAlTqx4twDqX18Ou59ty/B+c
JLk/iSNR855J3fTyulhvjXLNd0gmTf1xsJFO6qF3TKdzBOQ3wKz8SonJowOH4Cnwaugvba5Sy+Mi
yqOFZGPR7aVixcd+MKvUwxwInaMWvd5s60P9nOVXRFOl4QkiLu+Ttiv9WVbsMGZlzg9yADDMXg6V
9nd9zcATe3VBLg/2v3kmpb/8Y/RqZhsL4PwbwVdUnBH41zzgoUBr6ZTNTarEN5S8AYTc1wPUSlH+
oij9HhQA1pCUT34p9U+7kbNvJhtifTC3+KRp+ZMnKYaC5kKjW4UwpTFiYW0u2Hgnm3tm4ntfURz2
TaH8wv3PlTyIYAjSg+JUkxifRfOzpjXbTCryJqWMDZeT8V3H7U+ERu4z3ed3UIcexM7RSgKFw8VD
kPLFV9qXafkjQubWGCjdODTc9DbbI3GxaG/TP0VSQ6elKjLrpHjnu9KmQ55+Ez1u7zlUUBGJj/Se
ywe/qiYzVhtUCOMLCh6kr+9DINt1j24v277lQkOEAZQfnUV6TECvAO1GfOmAXUBdfLiZDGVScbFZ
Hy3eiQkfPGkeSjrz+QLrv9Ltc1m8Ly8IN5qRBRRFgPhb+Gfrq3T6CPyQarLO64bEQpxbhAq4O4TJ
a23+xuWrGiE6fnfM4gowx2bIKsgRWn3fX3nCihAGufQPG0jTava43y1KVSnQqWM8tlOu3m70pJZY
nmePLmx7SEGthg0/Wrh6AuAjw575uXNfqaHTZSy1KlCI7fHNl9ACz4TaAWVC8WBxWWO/mRijxRip
/T26QrsqgvlWVNhP+qD7oBBZ2D7B9x4lvhxxVL+onLZCCpt/TrcqSc58ijDKBuA++P24n6DAtGtg
ck8xqYNY6rvcfxe+uG/lgr77MUTohrI3bzsGqeV3mhygeXAXMoHVd/o7J4uBsbMpnS1xF3c44vnL
zdVTj41XqOAfeJuBNsngnehB7mKAoXXVrSt7trjiPEUlnpG2hJnNbcvMeIT3dTJKe1i9ipItFAfL
YaukT74fAmZY8ZIlVnyjQKBUlgiorO7ZibEr6ourbVmfY9YHUlxDzAeNrQt8xNmZD8LKkcp+Ropz
tlFzRyilwTWOkw1OxU2tK6N6rF8GWCIPs/BhFBuj53tyQWh7oSh5+NKS2Nr6ioW38rQ1WTFjZE8i
iYiI5au6k5BJv3Z1KW1Oh8oI0mY51B4FBZAg2tRMy4XDm62+a9hlQyr9s+nNHloOrRMJX3cLd+Xp
rH5WAHa0mcKuJOhsG9Qaw0GVWB4+uMuPq2av5xuwP2CcpA2xhymvEVYNWNLtA6WvBg2m0yqTztdP
Gwbu82/u6XwhsyIwW6fujROtNtkEkGKwmD3aoQHU4id6SlJT0+S3LS1F/xuom0EEOtL6wL+geArG
Jc1ntBxBNF2jdyrrnPd9s2rl0hdijcIJKmdRQfQwRmO14mv7dWFJkMJK3CBkLSI+Z19Aw2DGjPyv
HCmIlNUirM8lz7Yt7f9CgcpzZLVKW4z6vUnU971tKynNaQgr8rUoHyQVGYC3n58xvIRpGXPDaOBh
6G3A7VULRpsFpp4MRkc6sOwePQQp6yim6WWBXRHAsonynCgaKZwWm3VZ+kRfhj2gNirkdWK+fb7J
6MycMAczKYxfdnuMuP3ISPIaI9VV/fK+O2AQeyeHLdeW8yvnn1njOCLV9p+j/yA52PaLA5n44DNw
uDMlH2GzWeEWLekPzzFknUkk9XVMku5K50OMrWfbHf3RVdS1j5JGtM1OzlKAnUuIJHh+98FQtMVB
MDtJWI0vOy5OyCsKNiY4aPy34pK4lDs+gwgw0XfpYbDPXH10YYlmwW4icWVmh49r/saPSmf4XuUz
UW1TP1zHqvk0x27t4nm33OW62L2GguFKXUl6w20RigZL3Mbw6ngnIP9B993BRVAM6Ozlz/2p00i9
EhW4jK8MB2KAPOIK/jIKAZ1ak6FFOSOLJGn6tZeVHDCx6o5Kt/7YBN5RzTAA6Lq9EkGkttRFZTwn
rgMHjFSKA8S3LTNREAqmMAF8YNn5zun1domfnWMfcoD1PMdJV/0IBzG55xw8mFCKMCAVHJ8Zk6Js
ZdB9YH2FZrckHm/Zt3YuW/Rollbv8Ht4cQv3I/fnMPn2VcDZOf+UiaazXUFsWXhnoZq7bNLSMEbi
We/Z967GuleMNPVvEIDYvuFTQ9XbpMRvUs/O9AQXf9OZfSqgjmTjIUtT87ouUPjzvNsqJYS61MQB
LEElJ1b4AE4kNCet7UwDIbywEP0QAUPLoWG65Hti7OeFbgg0DOog6PtncfKUVUwG4a1AyCcS4vk4
D4BHx8Bn3mPSiePJF/HnO7NBQv2PpjqZ91wVjQJcMohMhzDXLReA6AI44p8ygxY1bFNPWUWUyfpR
LMlZIIRAXge0VXJ/NQSSrkSPC33pLBuvu5AWM398YdtBtHMPfBp6beAs9ee8HVT6boRq6hLnFhtj
xmKtSSgcoKqTeQq6s4P3lsQc3zCRyH4+bCBHP70SkvyRN1zKDOHAfLbMCCF3qXklRAoJqs9+z7rH
6MorfuZCpDJ2mNFTcYp9ZrogavaGMxupZ4/6GNnJcTzRAkpwegWC45RxhydVBO6c83yN4Tu7aRZS
i9Vp30sRsGoFqZirBYc1brFrakvm69LatdTc6LiyVcXjEkiRUO1ay4Z1s/Z6d/O+IOe+uw5pZBRX
KMB8evU1+QQJyuKw5skbK6dhevbpdIIWUD6rbhM5E0UBJ9jSP0A5K5rANAwsjjp2yv6KCn7gX5Eq
cpBZnuEXA9+Ksav747bWvFrfg3VyvuyhLmuNuVfBehknFUD7Om1vpp0oxnMbSC+PH3IIj1Waw/mu
n5Pwvw7BSYA9R6HbBCCXEAl+dJXTPl2kCZlZywrkZKI+miNQnjtLjQgW5i9WPptFDMYsSEXJDrN0
F8sYSLtJj53uAC8AzUsq3Yx1g5THnSje7eO/b4qzJv6+Oa0TRSrpdGSddLnkf7Gi6D6wl5p9DRiy
jgdp63O9NXt0fxdv+0zpmlIU/Y4RTOQ2xYwrApblviLlDBiRciGvXyMmA75h1TI/X4kS/2IOUBFo
1G+6gSMxrlsTGWvR3pzL45zWT3Ed2xijSvmQDJ2dF8P/nVxfymd6rLw9phMOrNGKf8CRGgUd310Z
Nc8eRZXDGxsR4/siWDDwsvgfegk8sdQWKFXczIJcM8nrVxB5JDaLvHx0AzZJSejBiqmhLjZe0MIr
4qH2JBQfTrfxtg87hI1XILubL6hSBbgOGeFVisEobtokU7yspYNo1ZsL/Q6dH2aKdKfyNtrmJbsw
LsIyngFE/2pqIAIzaF71oCBGka4TvpY7yCReyX64c32vOUQlkf+x3m2M31BUzhGwInXD5kMMpC7W
1XfYI+OA2oOX7lGF+M6za2bz6gMLxIZ0E2DluiqWQlcJPQHxzcHFNVl2utyQnfzEfliIAk8ifOIi
B/xlM01CVnUfe33QtkAF5SSwnLcgi9USCCc8peHDKsMUlYy9tfZGFkCQexUTw2p5qBNDJQyYmj7F
0+EAElh6KERzVMr5UFGwb/ULTRJilDT14gyONDCfwI/WqccEyBT87o91wcy/MA1JcLG2xITPKCcv
gogTmotnGIhkmMmiGU+tIrMidj/amBYv8e9fXpr++T1JFJyb6BbWVqsZBDJMwjrhVHrSNrO9X2cp
hXMxOkiuElQLavxNKT5k5DvBq6kEvEtukNegdqbQ5mMH+aAxNkVXHbMmrm8J/UEh7yWr7BzC7SQv
T6RXS28mxpxwruQ6Lk6Jmr9pZ6NQ8ZK54Z9XFFjcNfE8w0mWrr2BqjePvxK1Hb5AKFr8LzqZy0s1
Oaj/zrargkwq/kEuoKLXymZn/nrTT8I2Z4epZeWe5YWLwXFjuHgvjvgDYzDNHmPAWwED1JmNxjo5
7R4H9s7PDtQXH6T9s/xVD6G1Kc4ZmLX7seqRf9tyF0gY4qu9P2noTYdaHzH6dcm5hJF2kfGH9Fj9
AdHBHwH6XXZwcndC+5503iMD0cUaiVzx1Hj39Icbiv6E50W3//cHVwELgOvtxlp7AO2NSjL2JR3W
FNo/XIbQGFYNIEhtJAbGykv5Lk5TkSuo4ZBArP20xIpEiMaQVvchiQ8y3/mpFTdOogDZDgkjA/uL
9CA+FI0xj5fL5l5VQCJoDgBx/q4hZBqvSoKh/wXymUG9n3VpqzNbO3qJMzCdnhcLGwS1Nvh/PNbR
ucQp7cTWJrFHgobL890m5DrJgcdT90U+6cXyWRMMIOfBbRosgFQXEL787vv6teYjjcZHnfpMocCq
UBpUhwV0GLHjMODrQMcN2O+Y78qncofQsJHCfnwgVAM7PMRzVyufaMr6wlLCBZZobY50PtyO/Pca
mX7etFeHFRyB8u4pO2/P7s+1mGydc/R0VRnBl7hK6+WiZPdObZyjYfqLQWHGd43tK72v94nmqKwO
q+vTMOwlXhdZWa/qrhnS/VHNHgSWGpB226659fPDBKv+GBQ6VZ50GH03C3+ITJlx+9HHPCRJYPyM
gYMkWyNYlOy/jXrObQxcRUh/TSJqVzK0h4vhYdmA57RLRKprmrWHixfIy4HxXhvDiy3xE7as48+R
J9greQArBS7JFS5WJTOemDVwDBPcCAxgXQA+MNSlr/SkSKl2Vji2A7I678sS5G/42VdcoRhETV+M
2qKOVy2z/50H1LdZZ8lLUlVPPp5muEgmyI+yICRKjlkfgi5PLmDRVTSyOC/7c6mHWJvgFIw3YvjA
/TQqCKYK46u21yf2866Cp9hpE/nQnVNQkiu4WOIaznrjSY3hpG9MOHvqcVs9pE56WhjLGTC2gtyo
rJU9+C1i0EVS/J91Yb8Qgd2Us3qmGdnENBx86j3dacMAA/K5ywWseoyscVirnNWs/ONVRdhBr68p
9Y+7xhsV0CgMjbO5seiBCISJ3+0jixYmPUY4v8bH/zVS2J40HDTZSvDosg1hNBJJIHok5pVeRbTc
SOA3UJvU2IQcPNqHqgh2zWMB4rANX7EAkhvoDLCFdP7+QrcAxI1MeSayxWkZRZtD3hmit+BUGUMj
ka8WmzORtAkbT75f6KzM+ij+/l1C2UC7GyymF7PUlJaJJXEJyYnO/BfhFzWAEGDr0jVCtJ5WGZLL
i6ldQOQmDc5wjBQar7mSJBqu4+P37eJtjXPmT96ix29b5mPnq39grS38Iul0mihETiWmcIm28xEt
AjiVL9fHikFWQgrNcBnWBU9veHrz8jxzJRodmGQzH0rvQGKoBOx4bFhK+nPmI2JOFkx5dXtGrlsc
/L+8SvkN67Hd4yVGWVdXTg6URnnR+Of/oGwV8ZPYgmDnIe6c6IdqzmK9dkpoPur45+Gmo6f6ECnn
v/JfA/Z1hMVIHm5RMbShbFN0r1ozAdJ3kEUebQiDcflSzzQSsfJTBYu/WCZJSMwKX/6n5k8QVzRj
MLZzH6IiVfo3PPgBLAMLL2XKxz3v1IPNEqoAkAd7XXUTqC/xGjylZ38dKbnL5J4leym7O9omSl5z
MAxFyxAmxRk1POksq7Xfa3jTcfPoARHLJ1v9MngBMTTivvdPliQgdNvyRoO4uep9FRf0wDHrXLDT
Z2RRad35DYDOmFOtdOdBOMvb0WOEXLlBPpIz5pI95RIc0xZ/gsgX2r/IiZx9FCHgDVWhXqYGjxqk
aiEhufXcHc5PiwMbIjcN6qa5Hvbkdi3azFAIGkrNp2mcRcJpNcAAa0Y0pFE8Q5hsB43id2vtCt7c
RF8ktuqY08UjOMYMNmy2f+xvApr+pVzfvs+t4MOi/UcmxFVu4a4OJEqJ/JUp7GW+vbRZTnmeeFqQ
Ow6SyjFDptd5q/SynTVG1mJpYldcwHXMyJVVnAB6+Yx4BYeGdKGhuWQefqePQhqYs48MnHja/I3l
faIKhJ52GU+hsPt1MNcF9gBcWdG3i447Nfeb83ovWhsNvO2XgR/YQmmqM2EmBE0BSowQq52yY/wR
0eNDthHeEpGlWkO70w8cblvMEQo+lZEF5N6bjFM3ACmf2uT4vMrBD6Dx8j6i1cU4m4IwTvv4QF/i
UDn+Ka2VrYCgXPsRs1RPM6ZNFmPoTKcUl1stwzFcBEr3tfrhtOXTEHznbacII6222n2yD3Bup263
TozO6RYKHhZ+NWDdC0rXDIfdygxEik9pFVQHBs/DBpKCrJlfat0Vb2l+2exdKJAMD5Db7XKEnTTT
1OTN7Vzp/F4n99rG5bu3wEw/LaW+e7EIUg8NmUDcOyYZLGe7Jy6zTa4RF7xF8yrClWCvHpELYDOB
hX13lMruewLOZUecfXtHiVBdRhSq2BtGUb9mNvJ+q3t3+0Kq7z6BPIxNzt7SWXsCzBGvP3XFScSq
nvk6AXl8AkP4KsNV/Q9T/9bcjDSaG3GWs5UqZVdJ1+dbFQss4dakjhTWPOrFGP1Eagjq8t3TC/FV
gYwcpCHjod69vM/UpR5kSgHR3VEtZePyZdK71pOI9jlgJcTiL3A3nSKFR5mXhX8lc1LwRgf9NT8k
D1PeW8FZRlS4yzbpuRJRpC2tZ1UDRI7G/YKqVt/O6o1WJoV0bAkOxsCv6JXOsJJSZWRM5UjMK3Ga
oIdFmq16yIvbRaZV/UtSjisA3K86VlFVtn9t88zytmQwP98P8dr+EjzT16uUCc8yJ3dTYsG7bSmw
0/bD8HaPp0BJo7RF8k7t6mlixnXoqTad/U7CTDRLwlZXc153ZihAmO/U3sL1ekQHrhe2idgkikf5
VuOxWl4YvikjI2H+VrjEVfa4dX59USfY0EWQqbKct7Og0i02QOAmMK8ouXr44kUA8tvyR1b1Ze6k
G5+E8lnJ0LPl3xDT0Tyc8rTG4NrbxEyymqWeQjKGtCUHhDHYfiMyoQDPr5hM/xyrzoxiKxDbJCfX
qh5ceQKTVpT7UDyD0Ok1veJxUe58+Jp4Nw8YntuxF8+OwLeR8qOgoX9X86RJQQsYX0Qt13lXv6DF
sIISDubtQmAzdE1Fz1aadq+7zQmcrs6ZbnBYDo6okzejJ+rf6uyH7GM/9h42HLImbfnaGC89VsGE
sdZhsXlH67+b3rTRBzPF7e/yty9ZOFvFZDaMbNDEkLCLBskrNIQ86oMNBCVN7+H79jiIbil+/H+9
MWwkbrjimFei2efv8r3+30buZLsrX9jLMcJRaMpo3aTQVG1nFO2ojZevY1S47ORpxXLV5snYmN4o
7FEOwhv2ujFZLA3KWXCkQuiNhKUhEs6Z/UOuhPEC8XkJ31vmskWNlGmr8XXfiU20rGV+CK0C5PO/
6jJj1qh0h0g2Uy4oCL4wBS5Q8NbaIRcGFUcTQSO286ea8SDqrsjnfHkk78ZIkMvP0WNwS/ih/TWa
8tQT/VavDk3GRB99EMR+4l1UoADvLGEjoVnrNLtunzYSApwPUnMQSGgTdlYntDhZt692QpIyjhG6
LBkuGYeU46YjSJS1SsRS1UXihIA3S+NoS48psonBGFXRjpVG39+HI2+FiP0fwwFsWJK6l0m0ATwF
7bCo78qXUHraYF/Muy4TLxxdR1igbc3rwhJ+JEnT87ht908JZ7CwG5rWxL1VYcLThA5L95XjzVUI
28Hdg6MbHCox7QRjcZJsUkEePaiMqXWPXnTUmib+g5ozhesAMKgP9G9SR/j6oZpJBkykW3m/W2uv
XI+y158x05HSwrfxDWOgVn5hNd1i1+foDuYa6bRkcpVutSeBpPzL1BLFgLdc0wvwcaBBBgQ47TSZ
mIyVNCbCOMM0O7S6j7eHqTbtZ1rB6xCPMdacrawZ+Xbib0l6P3dq5bG1CDrD3g88oBJlnQtUTjPT
NqlYwmFELzVwqzmbw593Pswsp22B+fOsORetRNP9CU626SBt5BF0BgPIXGoXBe3Lh7mHf7CCoawA
YcDRc7hhVJVe+PTHjSRw5EdMItgPVtq8KkGZTDm/yTlFxsYgWx307lEnfTez7ERzmJ+Wv2bIBK2F
XhII1i4sOcf17JMHJDPJ3R1EKV3j6NR8DQJbUyQWYJtkWiQtQFN8dvg+K4zs/Q1O0VaxlNjJl9+Z
DuML2knCtAnIukcehYNCpciUS+QZAiOG5S8SK20e6oTP8lgg/8ODCwkYEEt95X0rY21/LW2oDG/1
NGmneOLkGPOnP5c+IwEtvYH+FIBSNW7KwD7OOqWubKNMv9l+oqMvL8za9Dd96ZN9vUOgKHQ0qV0M
rGdPVdGXOHfk69IAjp9J9mLrc+Q3nwYJ62byqRp49Ee0twMEWIzD1cPl4484u8peaCulIrxPyztl
P5P08HWCSLLom7Ji1abCXjeirnI57AbQqcAX9zXgyurVCuo3EmkxTITt+ucoYYkhHT0jEKW9/Y5X
hbY7kgzdVvDFikeApni4dRQs69GtStesmrJY7baLoXElKj7l1tA0PfcILGsbNCL/ZfDRUMot2g2S
LzbQ71nehTpl9WNvtIam99LmsydTIMiAQqJyc4jHmn+HgBE2vnKGKHC+Pgc72HhkEOnSydKkAqEq
UTr/HnPn6hE/bQrR9yHF/IKNlK05dolH5hUXKBz8q4txPVHT7t7tdZSTBvZC9v07ACGzDyP3IMco
ZpCxEQD6LmWLQx/WyDuWitmPkgHZfdofmVEXJF+ciKlMRqaemrt98gAoVhmgQCHIzXr/L60o1/CQ
9bd0v14bRAkayyLzHG/sdBeXR+YZIU92OT9WMvs0yLH7NNoEXk6jXSAiK68UvQjC0QNC4oElSoe3
t1LMVOm3kPpYhSdSGYD3mN14Ay16qA2jPbnFj1LHhKwUXxKRGNySNKj7+QkKflOJM4KTvzbiNxiR
v4FISRYT23LMyfR9C0I7ZSyDRH2EUGXbtKw4I2OL4IJsih0oeYoBT8XsXOS55AfFfXjf5/iKpsx+
+krQr5oB5uF+VP0awGZgwhwQkqRxmZDWw2YzpPG6V7/XlQlYqja3d3CWjvAA6UgfEV6fX4eM0n9X
F/PqBTIeCa64TdBthYe+z+/MQogJJR8TP7nb1Vs9WzRfOEECCgxDNqWvwfsct3UCWh12ePeU9Gib
2oiBvOocYaJ++62vSLwFxoO+WCIIj+cYtK+k5e3J9NOQrkjAUyM8SGcmBMFB8easGg2ttQjJQwda
qdyxd864gcpvQTGBTbEH21INrkgPfkqTDLym7fZYyhcfcpfbg/ZG0nQbs0sc6I/Omh1k8XoANghA
zJYiKofhfJUdgBLU18vEd9gOdVGheFCz47H1UdE3t7bVN2moH3ZpzI15Gu4jgXg2kTCUwJa8It5z
3oYnhnEBK02W+did/fjb4Fd4N3IGAdG/gG2o98JuqMgMUM9yTDGlnj2qPdfToGpc0zMRzjKwCD+F
eu1tnu729i68vW2nqvdpQqdzAv9L22DhUVZEHRdscaHuaCX50KEfQ+2IWAXlxczf4010c2/7Ww6e
9dBQGHBXGOgOyC7TXr5oMzh9n+IVkxNfl4m6VYxpApoMf4jV5Gtv8I2fYxsJV8vQwqZKoKC4Cgng
UWUNRYEKho9K7w+bj1ZRR7jzFJwtFZm7bWk237AJDD4g/WiMN0dHOuDnQns1W/Xxyusw8xfRVG+u
CHILpeHKftIGLWhoeoe8QfxERLoEybAQZhLnPKGoMrdN+uyfRI6jrp6GpioBLrkPdKzOduH/7dnT
iCiajCMXsQRutlLwpbPLiFTm+ETGv0FNWazgvY6QmH1HJWArR+uFwsZVqIN8o6uu+i4FJb/2IrCR
ms8GfU8SF+59F3WEmX5aFdULfmczy2fHuJva+Ncynwg38wbPrtVUxm79y3MIjMGz97JalPmyvwgk
4T2EeFgklndGsQNjTVO+IkWlk+Jj5GiqMsA0DGoZkZ8L+89CCtnR/9DswlT+mWLNSP4dUcZM2nF/
83cMtHCDv540vt92lJgEWslGq5bOSAew7pCk0Wi4kTT+N14aaSWalt0XHsBi/azS0zI79UdxyhAZ
lsvQs/TUMsllAu1FtsgYwzfTIWef9FsC/I9FUdURSsOVdmT8xC4VlMGpCmz3EO2CTEu9jbj23TYt
kvU12Kzr3HGQUiRPgs2qh1a2C1AsM5Hkt01PNycM+WKv+iFSAh4luRxzJ0tx5r4fuAHX2+IAb0Il
ClbdvOkynLuW8PjV4+CxLrWEKaHealAR7OUqF57RzMEFV62Rerrq3ttSK58UY+KCOL+6oLuy8Ov8
4eABRm6rDB5jdMkSjuDF/q4cMTrkc1XO5C2vswWAUeYvJ709WUrFmpxFB0kOG/PGqgrNGtIpifN3
CApY02CGmat8gImC+j3oyAZ++OrzviInQ93KM0KoowDmHkFDvfNnMqjpA0ebBslJytPBjQP0a4fO
ZpTocS2010o3uvjd0VDPWP1gz6qR/0+w1TlKKZjdpgGVJx7U91cywavIY0CZLVW1E80mtVs/nq6n
KdnADK92Ove3bBPknd0/zReJVsarU+5pDI7GvrTrfUObgKnGBdWTJKKH1Ji0+Rlyj+nXR3ThO2X/
Z+CcZqEotjfrm4R9+JcG0+HuaxXCYoccDBlZPLe5IBY0Ut2ePQT+W6XXaK6msN6lzsVCg5ANyJlW
LL+TcNvrv+kXEjtTLbBNnbo6HFys1w4W2d2qjz2nIzoIi9e7bIJ09GwPaxLmjsa5Vv1mHmHQLR+E
BjuSClJs2vn6KWiUVfBZjPH19wLwTA0aWbGnqU3eiCmFmW1TSO47CqsSnA7cawAxWVqTdATD0Kgg
FOis0mcGBCJZnYI6wieNWX120RFfyw3gss7LD+PRV2Nige/TXZ/phRUv8dW19jnY31/EFQdil5v5
rJoMHufUrZMOaCpIrmc/mh7R8a7ilurces1xbqKOFeFS7cMzVVWiubWLIYD5JFaSBSARvGXp9WdD
OP8Px/02s2mt+8nPSWcw/YHrTvODOl4K9O0j+O5Zi1Gd93Wr3isTC/XMEoIdxxPXbBqcKuTdDbhk
Xqk/USPfjfGR9O0nwLc2ickxI1SQFAOO2Zc8GGdXTgzrtrV6qWkeGSLiAofTJ9DhhVV1Ffjwu7SS
uYtCgwOeUocNh2C+kapJfcbpNjm18kGVN0aZFlkCSGh+L8VaPz2VSQIH5cdp2bWLZBWG4y3N7ulV
02Qvx8TvcaY6L7Utsuy5EgBwc0j57dn/S1a2zd3Uu4g3MSkWUOY22k1kg9kL2Slcvr2VCzWruHrG
nu2GbvaS5Qt+TBsIZQTHjkHgQ8fHmo/ygOCV1PEM/TnN28AOB3V1SR+fHM/8JpMfoK8joqYOEskm
E6DWpmQn2DQ7SZWK9mSXT8LQqDJATdxZTMipxqpIrhAVO0AYNgFeRcB6TPll2bQz7UR0WpLKNDBT
XJil59Uvdd8Sd8PndvUSu7v53UHC1/XjMRLgaDDP/Ubv7kAPs3T4FdyxmdvrotXBk1rxNmcogA7p
CvlJIXufxgea1Is+bNQre3luKd+0hP8eykMwjDJKrundKOsIBAYt0mdXWp1zo+5geOE2/dDFBq17
6Xdmmh+/KzYqz8gOuUZRjF85Wq4pzvvSDOHbopMRikSL8PxqMCUSuAi0xxUQf9c3LB4mq03X3+oC
Ajrjv36ng4l1qRIoiVOrT1kxyLLRIIyF6KOm54aGspcEs16liRkDzXQ+dLaSm6JlMFdCRM3oKyXC
9JFEyXUH6FgXoUgpRAmNwnsSq87rC3oobIINMiGy0fhuiJKYEZJYHSg9zr4YLyueQxFtIyjhQz5B
ZQHF3KWB2qAr/omDN7IRzq5dOmCixrB3xb6R4OGli1NsCYqKnGScpBshRw9bGoZU7sgppWa6Sf/p
PUQkRBxGke0MubaEMLam5nGvKqPvIoa1FCs5I+vDeQrpSVOmcczMHELp7GdpGpZNnlShRP6xgHtp
vmWysGeSZJFTI8Ktx+1Qpo8NS7B5nU3UaUTOnNA+lR5NkJc40le71pRkgopT+WfK+AcYgmIVu9QO
yMpDojSGXBqzvBA0NGm9ANosU99JQEpIq8Xc7tK0Gx9ZdJxorA057TvqJiZGEA1LRRTJD6GwxhT6
3/N7KbKIEg7idHxp1QvC7zBXbG4XTJOcAgxUvnWxZSII6WxxCmqCYHj/6dXvfE2J/fzxAKP+4+k2
dRNrZh4QIgU2XsdIo1o9hTH6BKTUxJbUKpHgSZfieKOojTbj6MjVj0rl29TdAPAHCLK3EUIrJAoX
d2q+APeOuBI+kdzd1tJG+hwD4n9/ZGdJ8TaGpMCIU7CMIEznbvlL+6VL6prZmrZgvqFrAK7JUlKG
eSLlvc2xccbfuMw1qUBkjA3lov3b+RtKGBrmYYcW4+QloJhaTovqdsFpSjI6M3Po5i7iqgt7A+v6
Otivc88pyHPgZ1eRMghLEzIjnbcWjzjvwCW8wl/zNX6zb/A2cKFHX2JhHjGnQaZi3yf2jg9fD52y
xXhfro2oiOIJM+yn3iRHcXdYOTn35HI9fYNH4QFiCU1O6VzgMN1ts/SQstPjTs8Yqnvhc+LgewoT
4zEX6addKKquF70JgldjTweCSUhZHlitxGCRUFmgLi4AvZsjC/Y3/sCYHnP0t+eC6W1py0AAZI9U
bTuqZBguHdVdWykK02gWpw6R3ooNh1Z4JOt6vr8VrHxWMMN0gE7+lRPfVIOTWFLBy1VeAOOs24PN
UTymkUr07l5XwGRbfRNDmmcyFHWZt/7RyWf6GgWM18SY0sdLe7YgExhn2qzwGTmlq5+8p9l/VfAy
VTf+KdLj9V5clYnuuS6LzoOj373bPCPQs2o+cPwLdDVaG1d6k11HWb3443LtzswG71ue9gIFc0Zo
j6EQSI9KKX+ubn34dTX9hhEsvuRe5qGuzH4EFSV1777tlci3jmc/UePa9VApMHyefNKWw4j4z/2a
FUNYp6H8fc1WaTbuFGFMV9gJBLEmSvDS/R9z0Pm0qddSFS/wOig/iCsf1I0bdljPk4WY8bH6kK2R
zNeI8oCniHIK+zzhWLXoTRiTnciPb2+E+NYz359K5GQh4SBWgbmMNj09H/IM2yl7MKA4Q9wDzIYm
aAqw+haYuMmvqozsZYIHpMOvAmdu0iAELMUjUcnNnl330FlCnaDjg7EymHMLABDvF4bHWW1Kk2Uy
gngTu9bNBNQLYJDzZ2ug3W5AMIPl/saqBryoTmIrgdcsdxbLCaBM6RdAaek5Qley64ClPAxqNSzV
gE1kFPT5sP9DuM9/OqbO2QP8NME7jeL630DcWCRtRWqFtu4lLns++14I6fdGkPpZR5k3c/kXMMlN
/01GVX7LI6BP//GaBgzVpMV50sqNuOlRBpdRl7evNJAwAntkYV0kpDk8t6JU3PH/MqFL1/E1puvB
UwB81qPLCEjZm4yitOMyVPFy1+6l6OsqT1m2oVvKwbdnHEvFG3RSAlVmtTLr5AY56lqeqolNIRzA
GAds6oR2oMKgUyxwynEGOfbwQf4TTl4VEPqoB9m8zDUkUPa96EaNsBPtUagBNLPcCNAFjTlNaMkY
oRwvr+ckvJXgWOfKoG9GNtza3hTzzb9PQ+mRAa5PxRcNR5ONzgYd0/MBjJXx7LWLS4WviLrdCJv7
SMMfiJ7+NDNttCn0+awytOV3dNboS2WU/u/8RvLTbn8S6nibwDq29MIcjDiQP8PGBQyNySJ9y82O
jaHR//WBoU485bPzNhOOa2gHAU4wuWTPh/MtxSEhyfC1asSBUb3JktnBN2adtb0mLGcszola2TgR
sOPj9UBdOvChyg/vH0I7Wk8qyG9UrrQSMs+r8276Ubi+YSnNs1M1b1/uKYUa79IiJFyiZWxgVzLt
xsxWqVAP99l4IjrkxpB14HynKws2zwRrfp/1Jvnc2Ko7I+/ZM5XIouVVCc6DKm4POX6ysPbJe4NT
96idmk4RuhsDRYfTUcYwR8jswLY15qRODHzmU85N5swRMlN0Qlln8TQWCNrgOZHZjQLGQivaRroL
6g5iGRohCPIP2ItL12BvTPZLRaJeUQ/0qBEhgvXTNqUUpFIQW3cTesWEJCJBmI46seI6oROjn8EZ
MNJPpPeJHTFeuROxpNh0XWHDGBbVafgYQWEUSScp12rLey/3tQsN2Cf8VTOtTOFOTaxXuXf6HVbK
5PZWOf1PiNtkLVu6YL3k35rDEn5NNTqqi0WxnhzlpqFs1lVFOAXvGYaYU+DQIfdeDSqKNbsY4nWZ
U1yK+/uitU/agi1HCKcBFozFNkfB+FYlUBwSOtlB/CdaPtfQ1GgTfNjG3z3BxDYOMtVIjGesiN7t
RyPbLXG0kd462aKOogURHlU4yCHJx4HXYPwQH7uxKeRh8pxPhXZ/jGluLl+jpDiC6amSGZ4OXn2k
4u2xdC539Bo5T0gOflw9bYw8/rkichD65TSdE1lf5eqF+GzXqyIQKcEO9XGW4Ld1Hr1lTiHHgFpi
BINWOVf+rjlmB+wUIGFxEgjC9L09IdWaZHx+OUN5MlXlno9dJ89+uJo0jt1xIoNYBWfVOCJ1/Ros
t+fVitLbaed+V60J9iiDqKceGTjN/KzAXYnDqJN8T1HjbvZweHTWjYhFtvsf1lKsJ+lDGkpy9HdR
bv9DV04/x6qMA71QXJaKHwyj7yWYX9yT8xNDSGRJ7ShD0cqhYSinFOBWfA2PEucRa0YH08YxnCR2
cNq1idlyUShgOYMK4AnJDVdCp1thZdqu9aNvFGQ1iP8aQoyWZwL3AHqQOQ/KaBVmsG2Y+fYbYKU0
tTiCFQUUZ1Ardwelf6HPB2G65nOkmZmp5fd5ewTzETCzhP4snJDEL/P3NYM2II2M/DU6ngQBJYIt
5M891DS80m4CQDjYq+bd3QFYGGrpFkzuXUdtmfww0kvYJrr8hZX2+i9pSf2qTXO07k6QhUGr9ofi
zeFOsJJs+LaVApaaBujbKQ8WqpePh+CzfDT7lEq5E7Kw8ueDbQxHIf0eZtRbY6r+DAFFBDWdb3tB
czlz/S5t29ZlfGgj3ETXOP/AgjQG0OiAnQTG6G4Ez/HBJr+hyiwSMI6SU1GmmcGCa/Idv8pPgxRw
klx7voXiQF73Z4ZZXTmSQCGh9MTxl6XBt5y3UuhrUfuBSISw23tzVtHmS8LX5/whskhfpiUKs+yY
T2DQSNqMy2HohSYnhjWcTWHiPja8+pwJ+xdNSql6MlGXGXF30W3GTUoE5YBQTG1Wfy0bkKNNQIiS
xWobG1DqOU3hlN6aJgN81eTeQiXt0nlF4SJSnOOa0XpUOrdA9YdEwJPYXPRICa0NyGp4dT8yVHT4
xcFBnrTD72CRAO1jC924YeJByG5PEasCPkvLmgER21gJqFdqL33PRCGd6qP8Mh5TrQWuHyyaeX1B
Zq5FOJiK8768FYqRhTCbcFdzqdvg2rZmSoiOoMbq8i63B20u2kddES0mPoNFUfpPZuxkCIrel+ev
LDR4EicCRLNVwbq76/xZbo8PjJPP4qco1sQ0AxZGTBvaAEdtyGLXVCJBEeHiNNrLnUJvqTlZpZk0
1H/iqvj3VctdRHiH3lH1xD2r+DSgPjthMR9olcOeQDbMQksGw6VvvtoICXS1Ujraet54YoOYQEAe
rje/+WripR7nI6u9zQJtIEnO2gayp9xPHJ09IF23EMI6vONY2/u/kxD/jkAWzgXqBeKEV4LAfYe1
0MaB5AmeZezUMLcgpXaR7BRcPTI/x39vxkS7d9ArVRAt5gRaO4mhDGIvr6T9v4QgEmThq2BM3kzb
S24XXLHWRTrSELIbrlDHBZWeKBqf6UVfKNie/TgsKVMhCOFMHuwgyDKUZ5wUw9MmSeK+5C5fYA39
VADDbIgKeEc+/Phm9jlTyKRfXuuFOSiUJIHlj4feKNCwZpqyf9pX2lRPCs7Vew2RMV03xhtv+llg
VJDGcaw7WRSyqEQI+b6S8nJiOBYBKxo7WLbkc/ltrvqjz+e8pEwNP39zohpZuFEj8+UwiNgrT6hx
S4FT3XYTeIWkAPxS3PVrKiqb002ErkliHtBsp1D9zVnl1GI+rywvJR5oVNW9S0oyrLe1KR6AdddG
gMWT28Dzzap1FaSEz8sUsz0iEdsuKWvNYGkq1Bmf+hntreuGfZP4OaNlMCKBt67Swi5+nFyXPhuY
sAogjBqUY127FkzVpv5OnFKTczbCDLzTV3TDh9xBbD9C/zb1rAdr9lScUR466OrtF06PCsnAg0ld
6UNLgjWxOPuI/ZFUMNobRPkfuIwGAalueQ07WsGw8/oognVbxCtLl4Wqz5QbXjSt+AKcrI6F8K+Y
H5qiQWcRYsp50mt1oU0lyaGrKq7au0BxJvH9w8+JRA2EWu8o/v10TDJvuf2NgGzWtnTfI0B//XNd
BypWbUr7lUjS2o3qgLTgLnAWyRRnC4mbjrdCX/wEH1KPS6ldUhqpuZ4nbPATkdlu22Vzc+97Hul5
COUoUvmzxScq+yR4U0qALSkKdvWeKyz/71zofOybfnVBAcC9orQWh+ZTZxWRuFNAuxFQNS2tuFaJ
QIJ+6BUlSz0AtLLnC5hNdqNqUNQXXX4baA/y92OTpUdVpOtxWqMzY2FTgmVYfG18ZbhpNre0AgO2
nMDsR2yVtz0/7PwuGx4aYpVE/Jkmp4GjAru+8dARIxyXYP2THdFxrhdvjHIYib6DaD83C5+V5J05
6Dvxu3sU2n6M8Mm9ciNhBlZuwdfM117WTfOhrqTKFOz/3LRVKvFy7zpGvfkjsyPIhSz8V3UBKfF5
gxJKR8l2PEUkCbdX96BwdJWS9rI4HsA7LqpACOXkD4W7B7mrUpgBbMWjLgd1iLoTOXVJebriR2uG
+I0tgDUX2adCIriIGwyX+uC7b1reQdoXLhmqh6DQXqeM7noudcLXAXAX2ymLqkZ4FP2bxibTBXcF
oW8Savo68iMTTPP8ZkS89GQFXJc0xJNn1wvyPt7GXPCmj92qrmEI3a/w+IGyTfgHukiJ+lZhyWBV
grT/aSmFB5iodgExia+IhcGbzKJ6bBP+7NWd/gpZrRFhvDDb2DEyklm15mwaygE1Wgpn+q2tG2un
ZfgISQXm8zKuBZaLk2YuJSGS9vcqCBJLNhVTruC9r2GJ5fAAcJKVOAJELmcgVnXzT6zibHvLocD4
hy8LWcXZs6ZZmUoFA3wlv51DhUyllzwpPiPK+4+3FevqF2U0/13fv4sR5FCgenHffz4bnNghl15r
uEHmGy8aTLHZ/xV8Rsa9ByMQADHrgWGJn6iCJbRfSL1RwJsG3Dp2dvgD09ufOLsCpW+s2PmMYQvk
zfdbSCObJ15WZF5YlqJ78fbVQZrc9kGmB+XCYQqhXvDWIZFBy34MQueGkrnPo/Ut5DwmXIEPB1je
Qh1e9//Wk2MMAgEiaHeK5jClbUYBfcc8Sm8sxkguUxltJmMkJahHVOBz2j/DWux7pSgf4BqNW9MN
OhwOcDKoZeaNmYqmWSaL5MVnNwQddpaRJo8YK6bQ3ieaj4ez7r8xlnb7The9NqSHCBvMmyeSw248
u9XEgNBQm6ymMW9CJgWku5NTsxJOALDmZ3qljKlAZrvifStsp49QJkna7z64LlrvGyu7uMq9KRfB
MGoJijU1ZgPixfQdvtSJTksGqUKZa7cBn9wjA8qRBP+bdgXteW7NvYj7kFWtdgfOaf5cU2T8Vb5z
lG3YNfSYMFRU5PLo9aEZz4LtjzsppeicB3tS7RBQafK7r6c4Q3p2WSSds1ajhBqTOswinMjr3ScU
d6rdy+6c/CF9anBtjF/ZkQN3CFFTR/84b9LX5mtXA+rOYoNnYr9NPULpWiXdKWBxlrx4Qrjuhn8d
KdzOEScjSD/C5RQcg5a1CuWgf2Df0QePBnB3dHp8dMsPrIFvGMjSZac+RDI4KS1Nq1dn83Zke1aS
525CVHcldJ2otVM6aNRMyvbCL+dOu9tV2DITXw5i9z8+atG1QCM68tZM+4Ebe5JTibVLOqWJuDSc
wV5QPeO2rm3nqTJjRuaHYuNAeqV6isuaxPkjv9me9oPU87Ft1tVAH63Fdzj36Gh41KD+gEb+JL68
VytUvY5v/oF/w5QP1JJhE1NAr2HY22wiWUH1EI8wjo1Y/xE3uaGz1FY81Jc8bNYs3TjE3BET3f/e
VuATszqglH6vn3muf7NJAPA45nQSCOfpVohdLk8pLQ63TuoYR2iO8YwJowI18Z5TA9nWp5KISKss
/0dkiMJmjmlLyX6CY5i4Rl7oXvJwV04Lw0FwDGwxdISaNMVbn92jsmd8L+vJJc3JfM6DU799rOzU
LKgOtbpoIFec2Xv3JvVmNtR1XQoZ1JwoiYWA2uYe4Mlb/fU3fVo5Zyl9DJdRXJfMXfy8Jo6FLks5
HLwuJbuk+LKxnfAcHHJmf5sSMXBTVEk+52WRrMzdRtYSffjqpBNu84ROCRHRoFG0yBdOU/fDtqLN
bFqeBhF7bUBJ9RXjoL2w0DD4c64SfQVLuYwe2QXmUVvCmjBcPc0fK2vFITMwt8HxeRp2rQS8eUy6
B/1E9wGm0kp0uRkfiP75DYX6jGmx4uLROhwKQYYVb5JyKtPPj0cinR+ww3yqL4O80vwZO3kBvlZR
TFJlX2pg03o77pRjLlpCNPF2R11FDuDVm2sPz6o9Z/nZXjOMzFG2cdDeUzGLqIF1YKh/iEWWFlJF
Smn6IXeMoV55YTLiZvZ43Ak1vRRyNfBLIDBp4LeeX9D+XIT2c3AfsgM6lunRYGCKzc7mwErRX+P1
3+DQAevGdmjN/734bDMLdM8vXu2re1BEqMqZvfnN44ytzJBzYikQwnmCqmGijPDeZemSI7bFIEJG
1RoNtbVR3DzsXqVekupvHqAgKo1MdDTqHF1VLPw8ivA7Ma901S5nbrQGJ/Kh/1YPoo8koSw8dJs6
dwBEtmJWCp7FQ/dvZaJgP4teL4sVT9pYRDF6viLXa6a7mthcpbyFBaHdrkZ3OHssSZy8LTdE6dHa
1R1nEDctSCcwXUuZBmP3clQ42c7AUiGJYnaL88EXFcH/4lTjpbXZwDIrcRIv7sfVIZhaXZzzOIy0
02p0yN0UfDAU/Et5Kd8pLyrPvzQyBzrxD3uh+SImzONNGYbbb09ptkx+RBwNWkcykwwaLFPzHTGc
QddFeQuXKvbxNoU89vYfbATjEsyZ+ILn8dEhRVGvboyf5KId5ZiTj69LlaH0gyeQKo/oBZkzAE6z
vMoLvep9RMmAXVjP19sWQp0g8VdVQ0Noeuu41oVuDD+bMwBtSwYTnRSfWA7Facc0xBFHKyiH+pWn
6aNrJ8pMa5HobW2VVs+ecscFk1cnHBHHaIli04emUTbkRHBStZhO89o2T9ZCByyzXaHXgasKie6j
Vm+Nd2Nd+dvbXSaf9ITq4m44COmy86ImodUpepRqaajCI36VQwaMlCUQRLTfAqPQFd5EL6TK5VGH
hCVWiRzrlAoQAiimuBJic/aYa3a/8ZdKP/tLgaFyTNZ3O2uKNE53tXLkclHCUwcY24TvKz8juxVc
AiL7VVuQbWIWVuVD0u8VZpK0m/+9YxYYDqJM1eHTWKlG/OfmpZA7b9JTvVv0TdXw9fbxsFIRS1f1
8Ac0wq9byR/a3l/K2oQ+sEFBfD2trkNGb4oejJiRvZrIUreAFnqYlPNMdXC4xeinaXSRxVbmOv9T
CtdyCpDm/SXt2/vu0MTxTOiNxyvy1n1dKRpDjM/n3Cj+rCXpwCV6wuXhmyurWrtf8XjVfxn8eZq+
Gc1rMktZBTAp2PMfSTxQ2kypfugfzolyOm7TEEV6P5DlOWBgNOg5hurzTqy3/8erltzyM4/Prgfk
eim38R8oz1jX+V1FgTOIvQiYjTd00ih1WVdNv7CwPR/PG0zbx1+z1FknIlzthjMBOpW/0Zpkx/dI
2kzpQDVaVkQ8nm/J0HGDfEEz2Hl6b2zkGQu2XWw7HpvpZH2tbpku09/it9N6yvbgUyQxsARqtwAP
NMfw4KgyIQiV+VCg8s6Paof04AHZHFYeJmBAsofD6JBmLBsOAWd9nBaUpQO0IK5ujnmPkOM72lA9
dhDMR+V1HGmW8flPi3ZMxzBs+caoZlrPM9ai+Jf3Go9Q83G9AuV2648Ppcj6VHbmj3z7OKxSbSgQ
NJcudlV07hLea+N//Httfd5QYLH4cc3aZM16qvG4Altk3UqIBU3Dj++kf8QWz8PhBW8tlEn0HsB8
RSwoL3kUlFFmYHZZ+0ZtCjpZxM0/O/ZEO7VBw5bOeQotwVh+6LCEnrDzmqT7TipMdSMEkBvswU34
CjzGZR6cK8rdZpBartZ0PJAB/jOCY2fnMn5S2DGugHmRYk4Bt10xWfbM1GdGSUg4RkXYXERaMFpk
dxWZ2c50Aa8wgqAa9cO8bArQKPqh4+9qEhCLUwdS1Acxyn4qX9IKLd3L7NM/GWIXuaN6CDqsreZa
rZsB/0j4s6jB/HaxdhXu0hJIAtLVBNFiBihHb7o2SWg+dvlZyYJAUpV2xR50YHGsVELPBGhYF8Dh
D5IZztqptw6WAVh2maGbriHj8ajiI6Ih4txdAx501t1e+nGVYslPBC328BMdXCWswUbKCn0PnmZk
maPnHhHpo9kkNyxSE1wVoXo2ch94N6dIMa37PA4GbJ8gLK10QweWtQchxDt3qOmKJriycVbZoRdF
2yquusr/7P9KFRudQR3vhMf8U+YrJrKSewEQSVgz0YeJWSf4SwNtv4+XZoO+9MRIfxanafxpAYaO
i754FUVRnULy4z3MdLy+XYgyF9QAtuXxRPa1IVEBsBIlktWVzt6/cycTcolW9GYGM1zHG/tqb+kl
+00lStloFaq6EbBKrRDVKsNsLyVxpM8uaDiGlNLPW0wEWbDG83vFKs1ZsiFWGqhS3uO5A1SQHGHm
WWDB2OcmFs99tk/umm9bYgg3y5ICyFwdNGNPqpaVVBgmEKczRAKJ8wPILhlDU7hETMZ/fj8EnJjc
AXVk4lu3WxNwe+nF59LxNgiL6yLwtsChikSfw7JaEZtKpfzy7X3MTXdUYeZJztxmcGxjN29WQZ3e
yCoMP7uBl09tNYK/im3J+cUzDVNQhhFdJnK4G7e6aKC6voHrXfX2ARqSRCBiTc6NuyYU09ShG4id
3B3FpIO2z/wf9pQgbkke53zz0L2IWnU5332bEE3KmLyZR+fK3JZVJ/yjo8UYX06WSiEGLOZJl5as
9bT79NzYoMRBpbO2cXc5555hmpqrptdGFxmRxCDIBOksXpmLwxE1K1WMmdyVHvPE0CdLB70JaR6S
j0UBmxQKcBInyjS6HZSAwQfStfPNIGpYoWPaY77C1JplN/Z5/R5ImFTt38sesHixDwhSkKqZw608
sufeh8cINZ5zw4YnnU4cNqPbOC+MoWITkaZvz4xPZ9CGYnxOIR6sRToA5cTh4+nIlWgKjNyA7nV/
zYj9v3LBh77LKNmcyQEHLsP1z/xTMVNGdZanyecrQ+JvgDm3gM5kSu9qXGy+CxKMMx+bVmfxCNBV
ffYgENgdaA5tzSNIuTx8zI+x1p0uMhnVrsNGvgeDaJYm5GSIq1cKK2z7C6/ve5HhigpUCRJMwEvN
v5oXKXLMs7+qbooW4U2DEtNzk0nMDG6+jm150DohvBqL4ordJTPHB8UvHB9IspD3TtS76IRsxmVx
QcOfDOJb6MvZPF4jR3ANfOhJTGdrG7GB5PdzOK33PtU4hhgA97/hHIfvheXWom/L1p2YvYzNr/9B
6JqTXiCkJrC1aq65k6R+7oxHDyoVFuZLnu8Scgifk395ATpYqg4L8afKzQhR26MQYX4WjSsLM/NV
uLWvSe+tipGOXPsKwCOql/IaXUaWnJtliuTcpnALuXg8Q60rHGVhUraP330zbWJBnzDIcn+xpQ9a
QowNSfg+SSFY29FAd6ytg4+Zxs3CyVBeH9K3C1mWClEMmuJLRuISo9eg+/A8EtB4B3ygSg9bW2Nq
13RbNA30HjWPgCpLbcEM5yZYslTa0NLd9JPTqWW2Ycv8GR0sRgxvkTFZ8NjjS1uaq0DTpHvIFRZh
i/tGPSL262VsBOHWOInokwgx4EWOo4LeiMe8xjuOJDb7rn7p3AzEEDct2q92gd1zsANEzjiZtJ+I
FzQICgflclZdlWGMMFikftZY6BOwmva9VTBsomxTyBV2IYK3WiSq0um8Oj2Xcyuw6YlO2G3GhS6x
2STUXR1z83RuzdxEUuehjj0PZoFKRdWLUymymoBElwOMQLjoICown2a6+2FNVEwnSbAiWEcatCXA
ZM/HLxRvMlDtZXlMKaYhF8j3D7MBp+WxlnPoHsqcNONhr8UMUzJPmu3RVd+o1Ln+Ez3Xw9rHdfGs
Uh4StgC9rxgBIHfFG8jjteJSdpojp0MlCNZqGn4PMkM/tRumcnaMHnO83CucGa419ojcbX6suDLa
6TQ18k3uA1vouzkDQkcg5EGcFWud2OftY6KCOeC+XMrUXfjP6hUMV53CUYYSgmNS5qhlrouACsb5
hZQcD6P65QNIWELtjHkZUnovCrdCP9EBiYbQY4OIK16+uhI09WvkiXYeOfiyvQaLa38iFEGLlbyM
X4g12080ioWlpjgfPcrB0k5HhPv4y57lMMHzXJl2jhsVkn/ReS0FlQueqGWMgqTdVirVHboKnsnM
435VRQ47kUB3htw+LbJF3r2IjXB30dA+qM9ztdfvX8ZRWrQu4Lrr8quz9nX5jCEp3n2roqw2zeAM
OVyEA1Ma629Wx+XBtIqk/4CdFiW6yCEHGQa/B6MnVapEEvNQ7od2p61ZJw/Xb202fDgSyh1T2lNV
dMsv79qcFD0vBU4qsCugBCJBZpvLF7AfIyEqoFqT0c7vbPdtJwJMJrie/jRtXRNgUyBL2X2xKimt
AkWRAp64AFs+vIdiXYgo2oQXLVx35TQv9vgFeJTUcau6qvSMMkjYlWIi0TnAblDGjxWebHS9awLL
7USt+tdsjDYGAoONR32LhIJlhlA5yKU2FZYDhVfpXZZkU37L95sy7cdMIBNMtP+t5w+zdxWWM/pw
4fZ2BgOJQYQvOu9QbiuKa4yLTJXUt7FBNPoSMz7k2owNaodBfmAjxunpS3PbmBPTgP20rvRyeQQm
SHeUzYJu1E+S+kGkYX1/Z9BMzj/rqNWxOUH073U7v8IP57CyhPsHdd2Hggj6A7HxPmBZmNAQ7dUg
LpHPnRjrp/7cYe60KR9AnrdGiJ8Fh7ZPev53IKsnNQtJvrQEi1gs2qh9ngTaKBv/ms/NNTxO5hn1
LroR/+3GVsb25bDeWnvSxLMkyDGMhbiiSmaf/zdkXw47x9bVtgBGzkWMQ+NPqKE7UTuUFsDMMzW5
wbZGoUX10I0H7HHVVuIkx5dc1m0toCVpcSL6DLtykUH5LUD8PC50oe+Y1Og6CYN8ig8ILDV2u+AW
CmRO8cMYQcG5Y+9r61djt3yW1WVvSPAwW34Cr7I0N1OOYUus7wVz0Kc4V2YxgXPlVSbShkeHJ3TG
Uw9ryaTzq8G0N7qT+HRqAHtD7THJQQtxa1SYhmg5ngASaPxzfGVKhGRBAFK8lE0972yswLiWmBPk
qiVP697XUV1X1l9NQukWmSq/MmRknByICOjp+E6TknpXc9Z6d4O+IRJwcDqBpykfKlRiSEQ0Y6vv
4AxfeJA/xtKO4CXfpFtz4dKJlBJ8CTIO5LVq672VjSrxFd2S8uq7Ni503nJhufigW2haZ5uQequ/
6vwNTAnMWIa4pBMdr8jISyF7YgPQDGQr3p7ef0myadYOYgvqHV2jPs4kY+ALM9p1iix39l5ZS+O5
6IziiP6mkE0tf+/MUYDRGsMlmf67S7guLQp84293myJSN4zQL7nwzZ2havCNq651MMHb/q3laDFh
fHf24QLVtUgA12sHTisrNaXVQrM8XNUT7WhFbyNT951pTMD2zu83lJtGTqLaDLnq+V2BUPJTLglg
s3a3FJGXSr2Q6Bp1O/M6MIvpYdXlNB4C+nk6WRKnLC1M3Ifm0/x2s/vQa3j0UGWxFWNznqc5jXDE
783/OhOug/cNyZ/bvMNaXau2uMHxn6n8FTijtlD0qNtY1+eiT/jpP1NtO4amlIsSgrcXytEIX0V2
XbKjnT/qwX4Gq5ZJaQQ0ghYjuGLtSmxyEv2ZUN79418MjjsiiYhPxAwjhB9NlwJPgar1GKxtyWqw
ZvitXS25uMXxyxrJcUreEylmC77mUTaTE/fmmacei4gYJ/7+Aqqv5QjCQwWIAkMu+dmFb09KP3eM
7BWWOgDbHiAQYlgkcWJ97mtuQ7UJ3Cgp46yaXdQQtegbFeYOIOIJfx2qELP19gr4fQky5mWVj3xx
0D0NLanjNcYrri5ROmHUbTcU72ea7NCOXdeDsEuAlNbj8Zvw9zwDsXkIjtvOZ7F8cFwg8ubXnRXq
SqWs712utoBl7jL/2ncTA9PSTXGa+xYz01cmmZ0RTt5ImWB2YxMiyuIMwNOBWJ2DMYeOvGA4/Xgs
zbTGFTakxQNkzhkrKSSHeSpleBh0C7X/MoUjhUZ48IPuTlA+KLftDvnTT1jcbWJF1kHlJp6GAGdm
pb+4bkyWB5VmJZalDmITvWtU+icSPIXk9qH9cUI82wifN3k3FllvfL2QR1EBdhLXevAi45oA1GWf
gw6TRzpbBarNe9qRjx2Ktg/JyBvKYP9tzUFhIpo/EoIQm5HL+9wcQ/M13Jez3q+Rdfa4VWcumUI/
igl3e7bN3wWNNbj4aVEzdK6QKrb2Sih8fdPqPjOGyNYx88/xxfyTeOE/PylTqAtRNMXQscjaLeXw
OLqjtHiufoFvJzq5qcLwaH/g50rIhH/wUJXAla0nGLDAkSspj/VMzMUfwacWtz7ggHVqzi9QkbNG
6IiPv9l8L63rUuopUmmVImkQWcYmqP/2WrJXIHoyIcHV/kEh2vc4QSCvHU+mRaw5f883pVGGhzzQ
OteH9t9IYJTUwRg7tKitN1qaViWW4drtHg9MwVqmVToAmOoyprZ4mNSsQ9exGftUpjW3exWcw7h/
maQilHUjeN6Dloz1qA1LZ5JbSMQRKrxeEKQdZmtea5lI5U+cVZjkBI/3/4VvQoAne0H/yPehOCdi
tuip3IVsvbBA6HsrUKayAfUs1rv9ZOEw7KwySwv+iBBY6PNgHOsJre6fzvDZlXvw6RacwkJomIxn
HzwcOY5K6DvUhj/1a9b/H9/OIazcCpNsn2bWQw/ZVPxSxcNgdiF7CkbhstQXX/AFZqXfdxvMqzqw
lTOGBr38UJH0Ajk6230ufWH8qKE1oNqVmAbNzULHUthgZ6liNgruGp+KwPKnJglwJmBLSF3sL2GR
HU5rRwP7AkvUZ7N2YjS66a2b4ke3zMN34AykJ8Ntd4d318aCEDWjT8OP0CJPzxGISstu99HWDogs
80VF8ThChNDniq8FYShxjJ5e3uXq082pJqqwz5lw72UFnBY6ajjLzwT2MzS73o4jHjOPk7iXlHUP
Egc7aCDjEaOoa80sOtVGUsEcvHgndf+wP+Vk/37vMIUDoPMyK6+jmEn8Q6jSb+Fi/R2w9DmmVaCB
Kbl6adduWPhcwrp4DGS3VcxCZi91CfH1VLcOPAB0idK+QBRZXOVnq+dsKfEPd0EwH4Py9wYT3W6D
IxUCNqGlBNoQsW0cFQsunkTeO5jTsbk+plRZXDHelAXxDkTmXZaIlbdY7M3rVrbKuPp4AJ6AlJW2
ZTLDNwV61IDlAqkYiJo2wcC3FxPc9Mh7hWCXqxcXbSw9Niraw8+7/o8RXQEjxp4le99QOezeL6a1
OqOGMxJA/Bml+S6ws+DnLo18PMFs7y2Eyv77OzxfVPm6ShVfPVz1bZKppXXFLWj7xxS0s/mHm6kf
5Z9lTF0xz7ugwumhPGCtGF1+7WuhRxjN3zVk8eP6qZSGveJeJGGwoaseJxb4upwOhkUgFPd7s9Dv
+R88Vn4waV9UhI0762bkcO9aLtWv5tGjZTGY5EF4583HCTm6PXdLdjJzjKQGHqnj32efwwUVlQCj
tB/jN/ZvT06GOkZHkeGADbZ9u0ylQQx+KTVS0M2SEOH+Z5aUqi0BnHfhcFyeX9rkHWkEJfNKCKTW
QXGrb/8/Qs55Us+xPgqU2CBDXLlTIOdzThZiVM/0MkxkYr+7PvWp9WMEVY9LW7YM7A+ugHX6Unol
5VL7S1gcnc/7VP/M+IHzLWHl4JcYTTHlvtPBsbd03WhW+dG4Ce7prjPR4eHVSK8zWWA9kaUamFhO
LQRdyvPCoIFciiMAn//7R2U8/c1eRGJTp0UZdM7DY3tBBLWh6lLDSZ4M9lMC8r/tfK8SS6bl+9Uc
ybD5+gb3zFTbSGWTNuocFgWFuvTLnTU/Fb2cl9nFtcILcyGvuodRSpYHaia+wDlGmprArkMVF35o
+SBDdJTloEEEs4CBC0AM7gbfcXUkGQQQ1e6EaBoprKAK86dy65SqCgFzy6hknRsidkV29sX0et8b
EUfSbdUzCHambRQPVZ9LslNWg0EmVGN0gmbOdVIGq2FwwQaCZyG+TiqDwyMOBSTt4M4Qf9iGbPJK
kvZS8eQgvAAw3TzAlqKwZasEQj9EZ6tuq9vModU+xd0pQWFIgWwAStGEaCenjbH/mkubuIuJbOxe
m62xDDItlBs+ExXXNbOXVqCcGj8K3wP23L3Ncir5P7+wSI57etXXZb2IbNJrsnD9lxpCtqK8ZBra
XPu5I61A+BkekYY1irz2vcZw4DYnWv9BIsr1pV4x7SxXqfrrCjtSDf3MOpiKMBZPuayM1qMBRI6S
NBzpeQ8VBZ8xhVL9jCsrfdv9+ijWeW+lNtfIQyA3HeStg+DWN59IdwUrla7NRPBB83NMvY46FWdI
rKbdZsQBkq8/60VGgJTtwEsMOUR2K3qfeEgh6CeIw9agz3AZSSHYAMBfhzk7gcpoDYKoQGPJJ791
kjx8109+RQzZZ6C+jBz4q2gjLxa6PpQieYDN+2PqCoVmS8BmVvbVbg7aWKC0vV/pwEiIy3JlNe0Y
Y9bkRbrmu4N6fqYydumd6nVeqptMfEjN2NIl8a8lHh1J/oF6HD3exp7YJNQ8w0CHyyLt4mB77/UA
N0Lbi+0rHHMkxgP7eUAPopyOaey/lYwiwzEncKZW/v4vwjLDH3xC8+Sgi/G6E3Soed6pWz8Iwptx
tT4N9BnNOjt0ljHl8vDEtOzpNG/Y55D7atmFxfdyaDXkS/jDNHpXjm+tr2nCHbUiofj4gxwFPXk7
IgshLssN4MNwk4InqwJspzKJH/K3AW1+Frdipb+RMfGNLBg4WMbxul+nE0l+I1v8CqyloW0D4PIS
MirLOAtyRG+E4cPAPEhqgEwM51rueZK5VUqnRoobOoFlEFrB908wi3WLXo8j/P2Xrd5iICPoWDKS
uxVQwJHngTNexgcJiwbcZkOFIIuHBBdNB8qN2HYO+jkOCK3CKPXQaDlxvtQeXN7zfUY7ZFIOknJL
impvAP2Sl0uAUHSUtNNFrzw/do2lUanlG58uOwHhzng7raYKse/peS227vkLhZkru9rc1aPJbqml
uW3GDHDYX2SW1SbLDhCUhPoOskzErhLZDZi91ygkSHRm+zbgAot+cIp/qfcUUeSf7Jy4Z6/XrMhA
ipswst+ZUovNrUPDGo83mH+DqWG+wsXvq0TIMp6ccjPuNavM8d8mYudGj2/u9kDPDh/PtPZePkee
rXnX2mofGAyO9ZW6+LWmQwXxnw0TdEbTO4h1gbyYtrbaCGfTYeYn+fDNIxnHb0lF31dK5aRZazF1
zJcSB8iCrpWHYQ/NywXi5cjLm9tyG3J0WsHrmtLFQrtFzX+dIenPQTepEHiPW9GAPb0UmPTLt6Pi
sSdRNWite6IXzL0BUO0i+64leOLZP4HfRgLY4ezPm7GKdVGfXle7/N330HJ2r/XVhzdnq20Pe2au
gK0/NfFvg4QfbYp1O5SLBHP6Pqcz7m/30bTCGVuSM6sLCL3l8rGwNHJ5/5dWWjzzuZgPiPRc0Lyd
MJ6dt21gCt2u1gCMP36a49cPx+OetmZVtZCHP1DMSHd6eq+1nKYjIo2JFnwV6kIV679Q2FqJD2aw
zYQ9s29+JBeePprt0tsTnprRp6B4FUD/5YfrWDxl39W6SurbH5ojXWTsTmETMs/RHFhp/pW5o2QE
0naCvVDavv84Yxovk/YO4njfu8Zu8eN0bLHfVB/VxPM2tvcSlPqufoepSAE8IYBqJZdL7jLYMe0y
Gt7ZSvZpZMILvJTXDfYEPn6VZ50lhl8T4J5AMvGM4aIbSXiG+6eULSFB/aijjFtPNpKhe1pDNnrp
i6u4CPJRDm/ufHWD+HvAN9nYtgf82G0FR9Wtx+OCw5eH2hGSnqVz1jtwtbd6hnaUEvWs6LLicchI
LvcBo08rfD/Tm1nWOcB7rYTYeDQd9+3A0L4PYFluslr4Y5eGNBvROb0032C2VTEj2e9uOL/T+W/G
giURSDS27e/fpusESsSqLGtdzNxt5B6Y89EjofZiw7udDSkU5I2K2m5IoZsre+Tc4/AZ7kb73oyl
/OduJUEjDYnx+vczw4k3voHfv8buv1k72XJ1tbfosWyYKUTvJGbkLk63evh1E4Widb2kAwNHAUMV
Q3tbA+4iwsfIXhYjj2MYuxNktI0FMGL/Xil4bdNFZtLFupCdrHSfiOf6DVdo5A4hgLDuF4rDgrs+
F0nLMmyz+kdJhGNXGa9fLC4CW5RGICRT1Lo2G7QaivCpR7Wm2NfpKoqFC6+Sx1OXp2C5BEAC6iC8
tB3fHOSBwapZqByl1bxRfzgzmA1lAjbIPicWMDi17Gat3VEZj4peV7rVsaF7PRKgJ036J2s0XHiB
z66HOkkUvDVs2UQhuxcWwbX6uPQYsYEqPUKy62tJ0aQOyEX+4aBPUDnRf8Fa3UVY5vnyYrnxlVdr
lRjlyZAX2BhCO+JPTvfbr1xjFIKAwuxYb4vhHGlppt4bTG7/9wZWpJBRP5ggimE8V7nE4rbTlxwW
kj39M93IfHc71SKomzuftBZLQ8Rd8dGe/+cFd5zv5/L8ald4jRTI6eA3sJFv92QIX4v2DvgVIN4N
chgIehMsZZu42W9WrtSdvHykctmVppQoGxNI3tKcMRmUqOjFvP6UVolsE0eCt0e/rbO3ff3amg+0
eynlkpVetSBe1Sc47CrKmuO1HFGR55F6tjTgGmg3QEt8XuRpGqduzCP6jCV0euEUKy3qi4T9Y0+M
ORpWP5pTcTj1hOCxHbYcvUhGp4huxFSWxdi/255h+m37SuK65wiWbMXZ7gaFvVOJKn3TYNZaySOZ
VxXLUBahv47KeuQWnHoIesDykPt8e47SIVIvPoS+6H6FYlRdwgIf/H82KBa0JKkf+BFMc8IEQoqM
CWCSVXgMyIrSRIUsDJv/9rVwxjbvAbNJVTbiZ8ANcNxXzSaVC7iWh9Vn0D5szLnWwtYzA9zPwWsu
ITvwTqGDYxH+pfDORIKzEQBj+g6KI6AHHlrcLGcLTBZBGNsxr4OG7x8uSIJTUr0H/CJ9dr+GOLAm
2oVweQEOHVXfl2ys6V27wjsd9pHnlammzDItYyogODVg/Cu2LHpnku1I2ulAKiy8ngKwvh7bst1V
ULdHIZ9Xao/zog0pK1ntV1LS6cdRV8ACR1UE0LAO7WNH72EB8zCCE9HP1PVK9ziHR7p0rvsNglq2
uKD64u1benoCNRwnj4EGkny4R6zJAVcW5b+pzRIK3u73FNbL2LEOStOhhNVrvRhJ9HZY8E1sWbZU
f931a1XjFSHNwFx16TMGEdxB+1xyd28Nydz5PxkobODOWYB8rXOnz3wnWAyQxTfR9jN6fcGCHSAJ
MlBYLYL1idxkBRV596xLV0cGIeG+yZZE4A96VafUC0P7fSTjvnFSViu0Z0pCfukRCAaebl7Qitmg
1O0Y6yiSKPO80WrmLVfcg6die6VDMY93m24EvSgg/I31BqNM3kqKObXNYnpstX7Cv9LlZcasXQej
C8UJiXNjfYwS/Fbb9ayHguRAUNjy9+oOPUbhI/Q2N8cFIKU14Vn8Cfkn8z9vHJepjcs7ZXwdnIUR
9wjPmgCkStnJRgwf4IXzEsZy14vrUKDJNt+8+Tt0UdURou9nFBGc6V08sJ+wVHCQSsZcWOHUTAaV
pTBE0U349jHJkcvfC4pocC/agwcvranPtugZOVxXxLmhNAmk2FxMBxhNnhyp41NQ7xwyHwrMHyQU
7Jl/qdvcvR+ydByZetUhwGdXqdBSkzZlnuVK4te7S/fzTMqTnQ2mMisQZGxGnnbKTIHdhKaiK6Bp
euR7H9Ww/gn9RKALhrmtFD4JOqURLTEawOAJilDVud2j9rWNgEIrckiB2yy5NHDxX8GYUDmrt4Z0
w744aOQsP9aneq9V/eNj1qWrsBtqQlIaRB0NWuryemJZOhTruKbMoAVF8g41m//AXd17gqdWanAU
D6MdJgHV0ebyi3U6dEe7JBb/P4mua/2vGhlfGaOgYMKVBn8YdMXGEOdERsi8bu9krYtKgmTyNYg0
UsmTZ4i1fSvlRQmHWD6xvfjpOzyX8Z5lRyC1fRFh+6n+7U2FKLZJQS7i5/Qt8M6ZDassXcwzZcxt
mEDNOOeq3ctgGp3VGUICzn5RwzySgqeEUCNNB/5wGc4sbIbY9rPkaVd9R1Bx79NEmgAn1TRLhVRX
aiuIYLbs5sSYqb3ZEY3t+L1lNVtFt8az4wDR1wGALFNybk2aNisagWCID6BwtXcd5KxCU89/XTfD
EiMRSAIAOm2kfh09xrf9bjygOqwvrnV+JC4GsttmL95YCNbRYnkEkqwz8dvKn+sYnGAtR8+fNVDo
C65ycUllIw5XeUMRJnxOUqrPCbJQRCDIE0kri596iLIN18PHkapm/hV46ZQRlQTWsxMq6eJRcNiT
o0XIzRaSCGKNL97bYBqIeJOPeruByjJyweCDhPqWUaJP92uHvPKLB2zF1y37lqoXd3TSsmNdTKJp
i7HaWj4TUJ93qXsdDTeKDH1vSahTlFbpFeIs36j3ep3hQsxZ8lp32BPaXsHL7yfOLl+abhGdK4dp
ndjzSTpAQTP92Y6esKu/VJokIqyoC+k2mmsVtSbOf28iWm9W7fhu+CFai5mwz8jVoHsbvMdAOjD7
z/2153mz4N+qUu2M6e8z6ZTzG5puwuPV0MU97byHQPIppKcA2jwUB2yI5tMzwhTA1xT2MkbARGXl
1i1k417XtnWkkd5mWRWTXUlgbOM18Nqv9w/0u5ShO0s+1xjFn/3MYCT6IMGGGwD0V+881D5iDsq4
5GScBmcdSpRWdehjE0TCBLeQgAab2IykKpw5VCZsbsk0b+dwAbM2Gb6s8g5S0k0KZR668XmghpbD
iDF5Bt1pM6sgSbSqbTYI5r8+UsY8Afs2S21qO+8ViCB4nrU4//ysq18k9AfPZeqxoLk/wtY8LQqQ
AnIh8TTWBCqxQsM9Fl+o4lGWGk1UzlKeWT6gl2IL31utGMHGeJNMj+W87ipIITRFt+94jfRHQLzm
pG+c4eEdk2WveLWwNayrhbL/ANfAuhIvVaAlXoO/GZW7AW3dRnIegt2HYqHqGYQtgw8Wn6HtBLut
In+FFnCFuD7cJw/1y+wRvQ/yC2rybpiumAuM2cJrflYUfSJS4fPU9ByGWnFze2wAzMmjneljPLkG
N+Jj/6C+4hfOUDuF3NlxnjiNpkW1kxeyZsNePiEG3GaJsXmzBJL9+o7UZHZXB9QTXv2nS1YfMoxi
tEFy0BwlG/r1rgEiD5SLxxRNZfL+nkGP9ARgzqKjRaWkdeT3XxahowbYeMJI6yZnQRncZXiOn64P
KCaOgnioAYJpdu12p26R7YgNHiWSm5+SVSf/m12c3ZMmpUWOIkeLbQp6KJpvhvKurPwd+mnNiwvN
2KSH+daEcENoqO+W4dIPpJ43u66la7ihQKbbWGypeNkZV0aIkO51RAZX2Rb8v9MU23oVXF7iSf4/
4GgAhtbgeArb1d1hoR/QyxpHvNUMcFdCnTiVwDLj/sHbnNXEBbxl4iAK28XHbMr0J4wUN/jlripS
kK65OSnXna0ZTHMstB2NFQEB71TOEIv3omxulVx9N2hWKGd4golfEGC/XNSAJU666BZ4eMx1kkq9
KHLb555CNPvJMN/uPVATUQ9ey/0XLvq6nST0+xJpLsai2hooXvNqLP8Nz+IxaXmQVbVp/V4MRTQP
QgF+NXZ+vI4ON4XLuAIJH2wf6KZyyQ2/mF9SNpznfrOydAkKDqQCCmj0/FNX4IRfRGebb71y189m
MF5SCr7K3q7RyF6fnJ5Wq/iXgI9n8bvB07ijzc8c0zo1MWmT35Fl2UDC7Tmv/ywaPpiuXo/797ZX
CpfNKCJUWOBynNewCFjj/ZxPCuA9JexecSbTM2yskztESSpWUJsYNAYNeg6iHMtr4Kjs54rwfoGb
FoUmrfe/HZXZSel4mTj6Zy6AA08D4yuyPNxX3Ml8VKpZZ7+u7MwXEQx+mwdUqVGocHp7AoWw7GL5
aR64OMax+2Jf5Fye1fD/emO5T0sRVBr11z73av83RYzRNSPnoJnf9pkTW1mXmwWwhhlI1zX0wGWn
W0oIjGjgNcax78aRHM26xKXdnJv6xHe1JRUZYyXLjpKwwgyQkcea9cNYPNIKT79CyMumia/tU0il
utsRcZizFCGMpSefMMFFA56LW/D22ACDopP0qDXiu/oL186mDbluPeTN8YZBcy9+BW5g1MN338Ch
p2fiS4A+YULXR8aX0gcFizm5mxut7xFTTnJQW27sBbB53pjyZVl+883uSPXHih+HatgQa/5TUUwL
zaPKVjYNs8yyrnBoiSPr2EijXfeIGRFBipvFcUfdM8Ha+pDppAAND0lylB7y/v7bTnA0H4FtysJD
IL9WNkFfgGErC4jQ3Q1US8B3dYGUmgtgttWgxroHgznlsM2GxS+BUbPtsfuAkUcJTbyokrqeCqF7
dx4JXYbjzHgbhKl2BivuxFagCsNzCuL1CymQ4PDiuGnVzTWtf8ArVToAckH5ZnWMS3pEl/Tx4XJw
TPDj7c4pNwP+tQEeewooYOc7WufYbqCocU51Kc2McASPeIWmq59N7Qnz+lNXcHGxTjhv3znZV7JY
TMN38k5/Nl+MMc0OvP3GNfO6pE330uNYH4ahYdwUwWTph+IDo0S9Winr86O6TY4UHk/IuKdPweLG
YCmIQbWFbCMlGnxJP9CL3kl0eXV6rMMo1JG3hnggY6OIBd1eR5TPhWeZsFcqxU4RYiTjLssYMsQM
i5Nl8e3G0Sl2CBuEfFfW6XPM8NoDpaz15kFyOYrzjtrEFuw+llWdB92VifaAT+Vk2t2tL+/tEKhi
Hrub/Rd32cAQGrqgHHB3xnyttpv8Xs/XyGHvOlWnBtrd69/6Aag0kbx9i+bltgPfxzx7MqwR2V8E
K+HdSUUUJtB0YhK7Fxd01BpmYLDEQvVqXbsWCcAT1MdVo+VWAJtIKgh7KvT9J4o6NsQyX7wvTcrP
UgF6l1Oc05CHxOYb9nIVwCNOWkEOEQtIaMTvGiV5epLvVYD0McRrd6njhc98Cn6GmMe/mAkYpGxF
B2yHIOTxjXjD/LAE0VkE86Ls+dObFvTwSnFSM4xPn+Nlhbo4Lmyc23YCXNMEl+aoVDhg5mLNngPr
oCztV0WBxqe6UnTgLxvyWa9qrsBjFeqFN9c4YB6HCkkhUtX8bByJZ50Aox6CKBAReYFmSqJbGL9d
vhFCs+ANwwKS+Ge11nfkh4JciwDUtA1NAyTr1YHf/wqQtboQWZT5PdR6hEr7f4f8ijJauXkSnath
0/5fSCcU8MyHqqQ8FfCTkUgwwPLQPPOXroM/CzexvSe8wqVvZan56/HH3SHZjotll/NkNMmxbWK5
tMPA8+cq32M+UfCsIhnftvUVd65RZKrGTB8qHXQbxw1ent1u3T6GIzrt6bqkEdNzj6wk9LZOjxvQ
ulmNbV+XJrmXxgSMTEZVSgwz49ysQnasfYGsia7BfheFXR0pAcqORO1ICjUymTKVKvmtqSZT/HMJ
ACZXH7KgMj87mqL4O9biLbPOQnVK29l9Clc+NPANW3Jo0EG98WmMS0hebUwWRzAIxkeVVDG9fYSQ
ywUtltOm1xrPGwKHCJz5MepUh3xmZOVbobYf/fJX3v36U4rHzYaBd6dPOv6uN1AQ3KHofvmtr6Vi
ZJOQ3gTaGMvrzANUmP0EaVMg4QiLZS5a3oWRSHXZB4FzdrLhxeS61gY0a7vvQfTre57Jz+ZqadAN
iyBn3bx9FJl6dO9f3oS9fTzmDrKyGXePk1L9PSYjrt4Essuc8n3mfpE4KIjL2gUcE05D4gBI2lU8
nw01KXhyMug1wJvK8XTAWq66KF5BMBq8/SyMY36JwTwrmsbarO2IzJ64PAMzHvAWynPiHPf+dSmO
WxUujyRl2VIRSlYkicwC9hmTQl54ExKD5d9BQVmS0g1EltnosMhQWVAHwxef5uRelFgayW/zuXbp
LWLqsRPZmZi1t1fWveU4xfB8oAXKrqkPlCKMRPCLReGkHn04FL/7rK9JGmsGOy81AmoF8dHbAWM+
jTc8J6QRUV64AgjCk7a8TpFY4BK8McRJvLWimKEFLyRRu6UgxAPkdvD2WadOG7zbcal4avxhSnwW
pj2SFOsI4Qp3EMWSDQuz6qmGZ6SEK3iL5ICSuG7HcmAiylovfg7dkD+A0cAMCeZN1D7L/tFBe29h
ULEX7qhYKisBEVsU1f0GgqeNWqGqyzgv3ezyqFuRgjQgLxsNIYtDVgGTTBfZRjxOU83ErTZWzAaI
Swq/DT1DCfoaq54yynllvCmc8kcXnDgU1v4MpoldjbwHIqBzO9xq3TpZFpaw/w4LElUFV7lVSgvF
/l8/OdQJ/eopRc7IK7uzp1KAyPk3zp8IEpqp4JEfmdcqXmC35WZ7grpALgMFMoGtRxxxRecivNJ7
wPbNyyBeGBZlTflcY5R6QJmeBMowZPYOAQmt7Ymv1fHK183F9iZeZktq74oIWO0Ra62N6SXCGa2+
df/r68I9kKL+g2B3BJ+Gk/CffIQqZDCQtCYjZjlR9Lk3fPW2bF1IXPj9X9Bg4UOQ95b4aRUDTfxk
r/BrOhPFTp14voMfRyraiGjFu0ByFFqJJLf16j9Yf45IsAmbff9b98Q8x7wd26viOWAivRCXzSoc
1oW4Td9CYnZnXZZqmKfqj8VKni+LT9xtqKZmdwaBGjaOoYDdf/2mjHeZ5CmQF7f5u7/Ygj5faCWY
564y14lj8rOs/PclO3kHtofg5cxJT9wP0LlqdCJkxN5m8KDyaPWaZSOQ6sEMdXdZqK/TJDvJ13w1
/S/nKyIB1Zqzb4vb2DBqd7GJb72tE2QX3nNs/woGg0wCSgBe0edITSCYNX/y7+NmMcW3AEN0/8c7
e+AORK0GKb1g1doqQ2qyechzJcFihs+Vb7zD5vhaha7oMeJO4CHovXZihMyaO7glw3KJZzN0bLSz
55SxArHMggeWIpiwclMikmeDHcilLuIk4p4HgIotW6YCmdHgJvscGMGR52G92AuwK7UDX3+5GJ5L
RybHhC6hhKe9JZd6+KTV+58wDc97elhUsy7OGhNUyB0pxTW3XdrBur5za2UpAvIT9bArHBy+8Goi
+OAau8H41yn1lYKJc4z9GCrim+eMnLrgaz8zPkgajt7cEFjQcofpC6ca3CRMn8i8PkyT5ZF0/HgG
46Z/xvVq4NNYZnTcHWoi9ajFwbXQg/gf7zczm6cwKiaLLfbmpdbkWx5a5F/M1luLWg07lc3JVs/s
FS9V7bu94VY88aV+b28jjho8kQjvVPN8UB/9Yd0kl5nlwv6C/d4IHYcxgFJo0JzBn25IyabxjQDr
QM0TggCe91DE3gHW81AbIcAlV3YtYX+oPVLXib8kEmKZQdUK5CTigwBggQtxg7j0k/z59afh6RvW
1UY1UACZWZwgyf+fEBmIv6rYHRVfBf2Yspr7zkfaQ1yN4VNXaEHc0YdGo65DObt28lvsCz1nEFab
UEgtWxQOz7KwEdjIZfC3e6K3LJ0zU2tUaTFrOqMC2W8/5UjrFjUTg1oANvjzqaPFn4UoLox/MyBT
pYCNQxiePIgEH97KLWmTCq0krwUs/pzTp40ErKlB3Ch/el7yBgqjTl+5yJZPTBOi2Wk5ps4lpKNp
GntmKdjamrRYIX7WGgiHmFBqi6p9XgQzPMWDR3MeoS0Y0gRt03dAxXTFqsQ0MP85gYsk0y1w5Jow
wfxxurO0ezAJcetkWbkye0HlwVFl5OFWOYsXHyQr5VG7Q7g+Rs9aZkUcnC4Btr2ceuhTRuRqySxD
vGUws+LoIQnS1ipXq1gQ5YI15t+/IZdV1/tCGj2dIlrrkip9mZdtvyIl/zf+Bgfh/VM8asNWl60h
ma1vv7wjxFjeYumaDz30i3eM4e92uPXfveYoNFOA0WyNs9WuFWkwiEeJQeJ40q9jntr5/XnFMOLj
SxEndu5avZNg7m0ieaw/Ft7F63Q00wn4GZoQNISb+xKiwen6wl8dF9FUHkRbm/h00FcoFObn6hhu
/A7MX8f8vlqe1vXwyQN0HQqnquR2fE+8IIlrZmOrQuV/EENFwGnnHniKV+5moiMUbAPrZHIytf4j
+s8d5LIe/DD0b9kSDPCZBLt4AxG+c2R1lzGWP2573rfsmvxpPM6XkW+DKTvt1j8JSbAqcOo7otGB
vs4Euab5h7NlgtcRkHRq+wreCvwhRXbgM1t9zK87/KzMdGBTjCFFe2YW2somvQl6ZQm+9ldy+IkV
qkemAp5WT/Ap3a1AuJ+yDF8UZfj32QivKAoKOFwpHNiSBSfR60Lc8SCh/LL4FqGJ8abJSMrEmAOA
J/3CEfUYrEa1blOB3JMe13KIdvG+BRQs6ahE6dX/mWpdcxcEXBquWp2XKGa2HIOzMrt3rmSVwMP3
q2vu0GyURE4TxB78gz4SYwuyjULLDqQxSceHfncABpcuwUAzr3KBu9gBSAAa+kdCUy9bfm+mvq6c
dYLK9e5UESKKZw1Destk2Xqv+aGjPVrq3Sn6Altfsi1i8jpuvFLg6HPLlmlQQYi7sn6ACBBXTAbP
XzFFr1cb/Gj0Q5iyUyIOaqIAjFIUZb5jXx3wxQaQBPVcXAa6mf+V5E+0AYqgYMlJZeeOt2Q3HYYA
5XpZhRcHcz+zzFhjovwiFKTwrRENN1+zk+qQj/uvH7HRBi+wubKGfo5dlVqq0516LKr9ZHfZNMRw
LFXu/vu0t6n3EsSYo8ppU29HkCI0Ra3Te3utsjiQf8Px9NgbTDIJCgHCC49Qz8672ngSxrkKXD9M
Nhih2z9EfZFBSEOR4o/gZGt6dPHpfpxoFAj86TmcH/vQPdKhrq60vFV7cgnaMOF31ZpA7SNMg+Pb
8R10z9KvKXaS61+33fI9Aj4+2Y3PnaTTo3gAncADKhJpGKoiWlrEzGV4XyYPdqqHFddPmpt1vrww
tTPZXfEjzyj2G725so4Mh4RaHfeyqZU7si9bZj3E+gMvrieY8jP8rpXy+GFXlZGUCoMe6qBaAkIr
4YtbFkq1/44FQgt3mRx8jp+nHTWz4Li57LXNWydXC2TaxxGcxqMkyYWQfPTnULme6L6DQOOjDbDN
EUY2dwkmwuX1Qq7PWRMW5Py1gqgZC4tTE4qXwv5xVyX3JFyzmT4TTXkIXw7CP6qjf0A2D3iYr5Nv
0mk5lTI4xMShpeF3J5FWykyeqn0OaXrPls+o1qK5y0JO7oKspJoyu3jVh8YMeJSZYRI5Iw59xhXs
OxzWdrE1nGTn/udEFj9WKbeUw2mYex1ivvrrKEJ/jMeI8jkyFzy0FFEOn8sx2vtPE/kygRYt/3z4
c0Iyhoa5x8qZnD7SvF0l7JfjMMVegxiZ/yTVybiYRIHBOQBjG0uwAumLpWlbewGmWUcsVyJFzb5p
KbK26YbgwJI+/JOJYVC3CJlDwnwVgeSM/jA+n+K57iYdvbllP2gKrVq3u6lSNyjHR5siyBjjbgOC
A2dImvp47Xh7/Dp+d/C3c6SJUrcLDVV+lgaTDRUHYsWrXW6wOYSKL8sCqjO3w10YvVfo1756ud8A
uR2rHnG8hHaQvi4hiQjxiK4h2Dt40pLLA7e4i3vgUK0YIHpxJudwKe+tY6kKTDWinLKN5rBKq1Ln
x766wQDbea4nSA2W1nTpPsfCwKEqN0sFcs7WlaSsSEFs/6hxvII7EjU4QNpOhVlSW3YnAXZS9R5p
f7tOixn9XczSKpbEl+Ye9aN+wPgHp4r+yfAwhPoDI9kP+6gzeXf7nEZ/AeAWryMWfSTkOtDbMBqu
gfR5hMbyLTPXlvPSQRI2B/3VSz26cq+S35E0gVk9nIqi2xk1oxEvJOEvfLhhDNC6Jv37uW0IZcbb
UltMlMqm22eFbMOsVYYRsQ4ZA0DzgXrZmrdeliA6Ml972aVAhbkXIla15aDdK+p3nTOFL3htsWSa
nSyXAfEtHBH4h13tMMtH63a0Fcoa2fC6rz3P+L/+LrW+oQhHRjVmwQXQ+efj81E0eVcBa6SsYZi8
RrKE85zEjeY4EYdPEr7BsxzL+e8xjVfabMBuFlXgeI1GBDqWHv1yT8GPg6gmO75LAgRHBook8TRd
AOtem4zh5KMmLS345S2RRhmCFtFsurxgpHwjMgUsDZwo48cKen0I8CioSaM4rAW/t/xZ8p+fI0mK
MEeeoaNPTHvSru2EUlfhwZPrsfyKU5lFOyefTxaMQao/+olI/bwWg4KGVNGX1K+qQpWhMuso2x89
L6V7/3WwxOaKS1lgo9cB8tWfTEV9Fw/OMusNlijrkL5rTuOeTh9Zyuuz6HApk0HAVdSNgKH/wc4/
BEAjb/JIOg2WQHSb87Q/UbjA/dfkuHFliZxCBSJUCBUeFoE12HDe1HpsBLcHlrUb0mssIKHACTA+
0ZLQLNI9pH9zTgnnmWqrSTA8A9NJ2yZOUGNaOQ0KIT55+lUhikNi5HAKFYsNPRFsLJWcY3ljK0si
39pXmulnmwSLOgLOugVhptW5jExyYrhUQSOcHsH2Yb/Ud53PKQJOk9RRkAKgR2ItFpVFinVc7Yay
n3xqqSrzr+AC3vkpTQU8MYwrS1Nk2AXo8TgG4Vhqlge0iRBMYX0rjLxeocsrQVOlk2uNXFBqWtYP
lDp9EztIqmWASsZxV+lpKiU/x1yG9Zkw+AWFZfFJ06jAZ54Pw1U5It0K4nQylAOqmQCE/MNDX6GG
er0TOK7/Q4+I5lJZeglT6jg5fIKcXOPQsEVs34h6foqvpuTlvkR6B1boa3pg7rlWw4C8VEi1lXPX
sxLxgkEN6HXukQn2B1rsCF47eJQt9zuRv1hWcEcBnGXgE/kxdr9pkUff+ZgTHmC1tdrikTmK2t71
RleIUzPnRNP2LB0X0lm2kxxsUJOHUrsYkQiCnUGCZR1J7zKXX/pS55z0TGC9KW5g/HKHaWRb9cQV
nRJjacCLd6qEpg+g9qpn6Fi5+GMh9jtQDX0BBvu+REXsTCzZWXsNRtNAX731Jm0DYyYDeOiqXDTX
zRiIQ3ur9yYot34lke6Kdela97gdUA2GGsjz3lP5sMuzLdOELo6xt/QFFZc7ko1ltI+CEBql4Ea4
OtobkYHKusGh9ABMurOUM7mn0drU7LMrOoWxfV0ZG5VvhdmJJrm6SPQ7XGG+UzsDw53itNpxoPtG
vkDDzmbPR10KbblVFYFTRbmYavIrdvhBwq9VkyEG1om1jUJgMz/nepJ4MWy39dYzL1SCnBdiiF/G
w9LZe/uqbL5sfEdTaRw/xJPzFBt9SgfQ2EDCD2QM6339IeuIh9PiCuZR2uyvHq09jaI9lrXsGjcF
bUng855VXbzxvyhMmLW0DKr7BzksgSk5a7260iW1Z27U/sFi1ewy4+DJ1FWRIYMGMl9u34ziQG4i
gJZBg9FePTL/DBKSrr7+MF/a8+hAL5yWhk4ERi6Ccd/8z2NJZCgB5zIie6zTGLcOCLiM/J7Q48Qu
He8kCO5kDuJq+3b9z856MwlaC/KV/XfINo7CS3SK4VO2od1Zb1JaLHX4EzooIJESO9L5a7M+agRI
5lQMIV99YKiRz9YKC0U/hcAZl1VziCTwp4rWpN+6skhvFf0pabf6qC0kIFwWXtQipYXDU4lNYXr5
H6qyYlbhy9ngfOBV3TueiKtgHGXyCArH1sdynib9asi/4d9ZMkpC9EOwm1fLqnpysR/Q0kBHcO2A
Oc16YkUkiJtnxTOqnI5Rwm7pO3qRGXDpOrZVx3Lr2j8kkP750gI5h9KjeIGHvU8zciMdMifk1H6h
RfanoxQ/AHnAJvSgNVNbBkbYMEGcBV15DPrkCpYv4wUsK2ATjMuB1OzkNoElNooWIQPfpZPO+UCd
EUCdN8qZIankDLUwhiiWlP6onCCNbCl2mClujnbCtZyaMMO5/4HXV+sP7+9xkSuYzwVn326FeujU
6xDiIJd3Ocg/BwF9LyoWP+2CkA/YZnwoSMlfFgZS3cklROMZ2UQ+DnRQEDehAyTiPOzkhMX3VPhE
ngdjyT5qmItcS25L61DWkxwkVF3WRPGoKYunt5xflp9WBjPx7Qz5uwvKd93IdDNtOdMpTMBvba+1
mrJABdth2YFkhVp0KB+Sd8iYYKkuSReYRK8QzwhbWbNHKbbFldo68C68ns0hgYRT1voKOW6NoQVX
6FH9vAFeApQYAKx4qUoync+tlsH0+tOmTSCPMzkAS7Er4ol23p1WpLCbMCm7RBalhN1cxl+Y2av7
OyBKDevI9+l0waKRM3M9UBYOT+XoxAOOEIdUpDAvbs063HmKBP+e1GQ4ei7X6aBjAnpc301xUiaV
K7mHRpouMk34m7w76Be5N4IkK4BiIsL6cTT1m+Yd9Kmk7X0ZgjdAjqoPEmDGTaTQdpQIIIymObtv
/SegYmQ9GFNHhuC4dObJoBd+rfQ1oKX5TAspV7v5gEnRUNv7gun66J/jDsEXFgyGAA8MyHvdcSio
Z2M3L1FuonWZ0vFyy50b3EunIqDGce0/8qO7X9oXyzAZAoTPJV4bcHkccZa3IGsrOC0Lj176H92r
VCeOPowsBJVqMn6U5CqqFbnzll78UTwpJKJZMjfgWvG8270hDrtor665fULLfwU+RJAXJlMH02Eu
GGz/5biGLygTYtjzLt3RC49KxqO6vJkTtdCEkKXTQ5bJXUM0TSViaYT83q/BfZw0dqceuSdEg0d2
Vj5upiKYIbFOlx6SZhkuc02NPGrNmR2oGxUTi3gaideFDH+3Ixq+AZdp8Nh9ECAAhjIvaeqD4/96
ZyWNwZQnxYEm2Ib2qJhZgMY+NLCeNywmfbQ66un6c4zML2E04qRsK6rEoOoiEmcaN4htxznTuly4
WVPKpLErD0NRcpUlo9t8bFCOgqM+ozS1ikNlYoutv6nOypOKO/JZrVTYBLNF1D9937At46QxUnr3
DUfHebT7NQBhz0xnzbbT50Euypt5uqwzW+aDQRbbJbvHQWluKfhykYE2RQOvTReQSVJUvYfR/csb
y+XDxlkWlabKvKUPDy2FIbm6DoyxZhUMbmBsfdmgJSHhjNNjeNdOjtLj4ruBIrrL5RlqN4rjNIDG
ZAG9uHqTRutgCbpzUJSiVtKYX49ZV/a7SiXbzJXhNmottB/iStAtTtAMyXONDP5rfcIjJc8sCMS+
v5GqO4kC7USKoiojHdYafp26v30qZ6hsF3P+2j++XfdRsDFTFDsW3j0Y3abTrFj2tz0L/fa1+ZaJ
EDdzCJy0FCxqiMbXEoWUqE9BizHk6w6I93nTEy7uk2XL5+SEHY0xqvJpVD4tGRvDIuezyvrll/Gq
tUgq2QOIWs5ipyJULBIWz/vF/uuJGb+Gidiq6Fe4K0kbNMeKtDkitQhx+oFGhA81fL6+UYJY9JJP
nq/El6EaWTCSRiJO/rAshZ1zf/FStUVA5G3dztc4JTSw7CuB5/t5cAJtSIiG8oTFflzfJO6o2+DB
CdhpNtq6BrDM2SDRFixwDxQaqBsC7/aGsm8+fxZZOKU7R0OsLlXlZHc+d5ni8buuZLH2zOj9SWqE
c/mjQgfvbd1inWNxkMnl0E5F+GYZX0m4OUAbpJ4/KVnfhvXuROdN7lGlvwtfhs83tOagYY14egIe
bnAaOTxlGGQphH0fG3YJ4t/7yVURE5OESOEtOs9ft5sbcjSJ/n37aCeDRj2cqLBQqP2klXEzaKkJ
VYoLwcJY/TzgWDcNy0flH41RrxeehFNf7YLVYnaqLTKHcKKZRw5BGbQhOLBgwzhpK5i0mRPVas0w
c2Z9DQXOSllTVF4sA3SuhYQiJnTSEeiyY0yJTFMzytYyPsThPaebt2gdFFM5dF0yUfHfpMLpou7C
ykgrLw9HMtunmT/8TiqmHDTybjEHSBXkGo8EGnh+fyQ7C+9DVSnkTQHKYVD8SGS8XGdHWzbQntak
gqcYuPQIFPCPBK6Wr1q6TewXH3iypNMmazQa16tdWACivZluNdQoeM33eI1JTym8NOhOP07wkNx7
kfZUDGkndDi+uHiJ0gMzUt6l5s08oqIfZMZXDyG4ngHRoxbhlc+SmOunXkqa9r0Ngd8UD+hADpDv
mJQGFZucNCl3QuLyTDsX4MAxELI6Pzjpu54YfBXgNyCGUO5SXD8GjCxj/LU+fVDfQdyq3LKhzYFl
3MSoGofL9pUn8yPzzBf/5VrSYLU5XqkWpP0jic9y6lcEkTeHABV5ZfsH4fDNUyP9ewo+y+OGI4DW
dXyMrnPouAgVfdGTjFHjz2Cwl0LsuNrzugxerSi8KCI4FZr6T/kLQBbS8XBeW+gETaxqkZF3hqmO
AxoYUbiut3y7LuV1FVlQLN/HpNHIYGlCOmmNF4RzjlnDeH235mATpRRiH8cbf3gdRhvWY0sJ/28d
/a5waYhevQxBImZrbj+qjv7etuklD0y6dN9xlr+1imEg5Jalsiolwp9MxH2lcZCM6mzYJZVejWWP
2hd9JtCt8UCOSn0LebAdEtM8QLwfYwNjTKdsYViP+MuqAhih3BCPUxySf5MwYAz4SRxl1HRhGGXE
CD6+/SW3JBj2Yn+1qBEm7rHI8Dlz2leG1hf2ElfaJCpVcWUiq8FSimiauTQksykBqfjYpvEsMZct
pObG2s2lkQ+r54furxq9U6cf922OnBfa4rgjsp0ApXbwA4BU9f3wUVkMHjf9ifnX2EtWq0mVHC/q
LFqeHxPwyI0u3mlkMcggAtCaZ4OO9NtTh3/H56k7DtYMwGM6Ne2CwfhVilbwmdyqkgmHeAJgQmCQ
LclhPwwtprZAU5UdXyizmCEGuxX09TYLKj3zMXc5YKYRB+ZWrRCxtXv+DCm2xpEXThUoVl1aWNKH
r5gF1WjH6lV5Wx/VKsm83zxi7eha3JvrEJUcd74ZdzetIQfdUFqwa4ULLsInnFHtxKy7GElQAr3j
ANWdxbcEcAmBZ/J3rB+kJC3AFybgzsvLkOZGmG6gXLanLBS9RgRo7NrJ+hUTPzi7jY+73fkVcno/
JV66XTl5nwAvIpy/jGU9TKXlrVurz3JZ/DMQqCnNym3uPR1xOmvdEb5cexDboe5mWsk5vFGAqtgR
8DJzbeo8u0pfo6nzzK7i7WTXwmuiAoQ2PTAQQrXFIxK3Xr23Vlfy1CU6M0SnzQcAtAikiS55TQ7P
10tfsKZaprZWPGWcvd14rCSa28Gmt/ICRBQBzGwybAuD7UtTHKPcnjdmVEhQWVZzRiOzuRrk5ZQL
lQycbtVs5QidAy/0bEHWq3E0qfwPM0zFc8L0UbdsREexxUJykUtUg1hhuK4X7ce8ai3XrtTd7Zgv
1RT5jLCP0bKS2gTGEE3QDBNUQkxm6JrxW2tZWpZ3Er9WwjFjuNNhuyUY1y3YCr0A8pSX1xwFZha/
R2KSGZsxM9A7fB3d9F3zTkEXfdgIaII38/RIgc85Hq9NLG4qgRcRp30X4l/iUdV7tu+UpRUfavmk
KchyDzbGmucu6xcu1Q2ZJYkZ13sNJ3FQBE0cOsY0HeAoAiXmP/RRBxnEKnUEklCu+fAmHHtGiyZl
vfnzq/2MJ99Ei6j/6Brykn6Rw/+xgbRyvvFdrZno1zhULGKmXoahWjbQ91aFyxbLlguEnG+rLDO2
oOOzMU1MJCfw43NkV5hDrSm/sEv73cRHH5ca3d95vtRoGn2DusD/K6Sitj5gI31JLNdRAFVV40vb
p3HljmOHoEK2ZdKV7wPzMwdmvXC4cVmmRParNdpHAZdRGBKLTLlQLxA9sFQCZUxXZLr8xXRXNxJM
Ye9MYSwyjuAqc062hJT/QuZN4AvWMXZzmkJPZfkvmv+QsOoa9Fkq4FCPG86qb5w3AlaHCMAEvNqc
zGhGzeZEODYw1WVS7RyMSDOVDIxIuVIoMBxg/QzoSaWLeORLPF91KYXffBFTPwh0mrXwD5o15YOj
KBYkupzpqfSnZFUoGk1pDxVLlv9E5OB0uLv3iRRhYt3lfIyLlk+bFJIc+ufH+nhduVGJ5Ps7SKJi
EHtETaeVWcO1V3uCR1Tt0yMeQpec/4xDIewxHvN97Jq8L4VLLudGfvtGi9V00UPh43znfcH3RVKk
jEwYLjaDnhQxA5NdStP3zWGivr/N417YZoQ62VlVwaKEunGsYYQZ9i4/o6L5NlXkT/rZ3/u39dCB
6CBaHnPW75qHulOemiSXB0CdI+ionkRNolawcDwehO8pkZDcuc9ruyjT8WAv2FiiCeLTT7ZyHt/K
RLkbpiP7bxuzTGH0EVgNmAIfTlhNfqXIiGSbupJL0pf+JGNl/H32Suv/+2VU0ogoDDqvR6Sg/rPd
V/2gYaZmlABYBrcTMJ/ghOZeb1xdkPOFDiKqfYA3GqLM8B6pazHpFXxbBTj9KPMkHf2NeRMN9K+f
qzh1NbHsRR6OfK3ZZJqQdBRQu1KUTmjxULB8A7x7rfC5rNxZzwcFzBEDmZymsudqoIBJVgaGlU4Y
X4ueOGucat41S9/GTmIdkn5Nu2ZtddZm7BJukPYasCs9A0maGJtvKW6dvHwC+KfDc0e1KBZCUvrY
eIkzhyRSwY9pXBVsrcta+DmW+xk1BBdh6k/RDj7/PPamibWkXykLfhP2Xx2En9Riz8M5LNovFbDJ
6GyE8RgwAZ5fFfhb5Gt0VOlfh2RHYYU8ifzEe0DsdPObGpCuzxTNbs0/9sSmbA6ikmu5ny7s8CWI
8eqCdLjNRTBjxcdfdeVPPBMJUZCJ+ewoC/+VQfVxCy71JpJ9TVzmPFhN2EVt29sAOyTcNtVDRD0S
wy+LcusQjHsJF5EOwPuc5/uiVOGTApM6UXXkPDigYtss5A+KM/N3HewzrHXIg1O6maAXEsRI3TXQ
VSOq3I8HYkkIt9IWfasEWLkoBty54XIwmKuv7MojDuZ4k5fai11+31jk/+wjzcrjf4mM0cABgZ+X
e/xn0aPz5UNN8mg8wy+8dxib8ABQPMHY6YBe8X5sl6L7tJMIod2xea6ZwLXC78Nm3m68ogcKELzm
T691m0KjeGbbw3Tn7n7rbXgzhJt5jiBSRrIu29leczSYGf4pmjXTITwTkiPQI55dPEgAhw3YQEfc
n0eBfQG1B9nzMXMZwT4RZkqM858lRm4ek0Y//xDtmsGAGNS2iAzKRe2rJIBw2xQinjE6G1ZnMpnh
ao+sdtdGYiVUwUE+TJf4SF4qA0S6FI/lE4xMFVxIug83kFbzI0YB1P8u5a1gilND1jOlHXgmPgCG
eJOJ233thZNOvJ1OnBHlhXjADqkGnEPoCFleu0P+VV1kTbhFmQN184CPWkFE4qzoNNLEmY2gVUrL
x+qBCcnjbn2IXl0qZmSH3EWfssujsuUH/hLbopCV7Ekj6xoCv8F2JJ+wdfdnk2HiVWVmT1VDzuy3
6tNNPM7SN/vAIqzvOryvaRvzSe+rarqPPZ0IeQ3qU0blFKGrNYbT39aeIUmscDgVLDVc0Rk1A3Pa
/iG1Q1xu/8Bysu2RzlJfxGdvkWJGiPL3Ihngf/JYEKDnJ4OeT3aZE+TvvS0b4ZaU6g+K2CpiAcsP
1NezcLFLJWLCdjR95ZVUCFbkNgi/8y14Wasp/Md4DRiw6Yq5OuaPiBk3FMZCzqupUvSYnaCQ2zvw
l7HMbgY5xyYbjyezzNbcBI94Y4qgM2JcdFuxRY85EDMQObsmozlPJq/Ffm/U4v27UWznViOxEw5D
2H9E2ZS6ZvXQcohlHPjnBC24Ef5acaHBV2ht88bgB5AwnzBlCe9UtRst54lFLwZJphImuklQolCv
IMfbi/yFieu83z9EuzQ3w2Y8wK1/Ux+zIm/rhtyjnO1gmVTFDdLboUxDmQ1hfwjtlmuOano/E/Q4
II9OAwufksYAekdDwP5+Zu93MVHiPt0jmYVPwwmiuRVIG1F+GjZ7kvtz04HlDf7KK0MVxatdd7kP
tIygTbbp/b3TUdS9yxLOgrYAzqisvr8SEqifNDOuO4RmFvM30AA4Z01EE8DJaItSU1c7qePrmLIV
LCd8jNu56F/F9nVLmiC+J2X06LVU/s5J9TtuJ90vjHlFzvAO6t9865CTgmBpwXcG8PhNzSYV27WJ
En3SPhNZIovJIHnxjBUFGwvrtBEluKUs8HByM7cEJ8DoJwDkYzLgLPpGhSB+fvnf5EVrp4mrbo+y
KoPHn5sAFhl0vllbn5oE4eOWpknaixh+pY6F/dMQn8AyUFUPBFJpZhprxpycMHRp6ymBlkXH5NCn
34sEk+UjHUluZHH7Q550fK6eid/fOnVpVgfGiZkz7OZAWUDt/ml3b9sQfN5rehpJ833bLOXLSS84
a0ah2b1RY1YjVfzNmgMvRToMwbjier5MwUN/Xv1FP4MYMXuFEzqrU0RNYNc0NyFNScNEFJsbdcWx
2OBUPT62BDNAEdvd7byVAiUlErIuJxVfXHn3JB30mkMg9eD9IYmul/qHXatpqc343QL6uSQAj+TU
j+tfvVJ/ZVr086lTz8MH1MOJXsnaFeTFmMzoeU4t+7OnveNkDF4gwqnxTGiyQKjg8eO/EPPlyUwF
C1FRr1SCmzE0GrhFsFng1GMDkWOza3zxirdBaa8i/i4EQiyJGP8TSt0UUscd5YaamdoUuGXZOMPi
IJBnwicCUuZULeLXq3x2iO9Sa9caap6DhdcwBQ62pzN2K280NtFfXjWCvSFa7Ll0LfIIHYTlzB7C
QLYx4tUTzXtI0fpkBIhmdxscqcmP0JTg696XdhiArxHDc8reYi7ODgb9iraNloqSfoCqmZRA4cpU
qjhGpCwdZ06XitHMu2/+M9hGBSqlaE5vx8FYjM6+ekgBbbhrTje8NHRgz9OlUh94CrHRuMFNLs0Q
BcRBx9iyOe7m0/J3I7GWiH+ABeQ3QXxnXt3zLYjkfohO3w1Fi1cbbe/KniKT3yObnW6hJrzeWnwp
SfnOOctyHSjkQLjEGj5yVZeTf3PwM9+O1lKLY80vimGfd3DTP0MCzznMF0BIKLO647hzpejxK9bc
7tNd/1Tf+i5Lr46S+JNvA87CqcvhqsFWR5xne3J8nHZWL5K1YJtRr0UvK1ecNrDiuCGGBtS21Uqq
3f9QOJQobfVtrlirXxNvgiYSMCrZj0FiIDuQlvIHQzuuZFMCDxfE4sfv5JvvluHrqZimmH+SRbcQ
km8Wtn8ae5Aoxu1Xqeu31pp/sUruFW4E5C8uVMYch3jaEX9MoXEt5XJAC7j0gz/tqcNWGxud77Cf
VE3o/tyPUbzFgKpklHdq00/uBDHDnxsV+6RPs0Y6Ko+G6e1+BBicqFeZSt/UNjywASzWPzq238fz
0kKLiBEdRgavp+eZd5FyBU6Fky7Q3xo+kiUhtYYKTUM4PJZLnvyLxjrFCKehql/FeCsdt/1DB/+4
jXwomTQprBTd0V3khW7omPqY9AosvK2h5J1VEooYmmZ07kxHdLqE+cFF00vR8dpbg+Zv26EhfVid
q/Y2y5n2smo9SxwSEgvOoFiPWW6CK9lbdHE14AXGMXn62weDmbU5OHtMHuROpYuXV4A2C8k30dP2
ndJ/8qIzXPreODe+DSDJVcHlUAA7fvgGvsuvKmOvLmpTJv3veP+4vymF7CtTora2rpd3a5ogHINu
x6BRl8/pjMiy/uG5uWgNy3HtBtxUuQtZjv34e8gTA/zUYUQxvwbhpHDJ4mtOgeIwL4yYtzGrLleQ
ikJzl1FplqSBQ7nVgapoBFmPebMGjBIusNUAGakTOd7BqPjWd78lBdS7WVCqpdrYEXsnt7bm32Mq
2sP486tUgCyphUpNPLgc3YtAGBX0HVsh9llNDiP32/nbj70HpihU4xKZ2wRpF6mDipHKKZ69YYyw
I4p9NiSolNOZSd0343DhWiqSBFSZkw18Jn6hje2E4H/WYSDXQY5JXv42Z7+MQOO5jHGFBP1vwKBA
W5+QPA6g8rskpUF3Ca1QdTHxxbqaEkDT5HCspWlKRTFhZs3pykN9byLH/U1B0CBLr4TfNh7gDg80
9gaay3kMgHxoTXsZXz+ttl2gfqLvYHAhwwQH7PtgsMfOuRBDN/Gt/Hm81fcEYgIaNCf+5G1AjKrD
MnFpE4wLrNncVDHTwaFDTucD7dpsKg0/GyosDylVCqPnTX/BgD91VSSzikU54dnjwMkC7j6VGHzm
v/4qheRCf0wSAS3zcenR0GeDedyERy5Mub2Wiu5YkXlbxe11xdw8ThL6VdnAOdPIhyO9z2JBiQaE
P98xtLwUnI7mfW6EDvMmv5JPh6urStTZFbrCX8Iy6bKO7bm3zqBkYbogGfHaZHeeF/oS7ufFXuLC
HVNMumZ0OeDrjGabBO6/dQS2qjxjGS6wBNx7ZRbpwRFQgXnT5dR4zlefiRU8t0GOFKb0vXK/0VKs
5h13D3YH9AM4iRHcMgN+vGhnBHbhmqz9Bv+BtlgWEmiq03MnHCQoKRfjhWU2I4MSOON/T6GLdvOn
HF7IbQEX8rbSME1ydtmnGlAP0AkAmiu7t7i5R9S34xkhw4evZPqm+vYy5tp+pfiTNWErCYNoXPap
LQxqgbP0zWTKLTANcBx/CKXDnpRzvm7bx5lAPDZB6E1wwlQr5nMoyENtBTbYNARXOKIBmtPVBTwN
4madzASVseolGjDbtDsDGYCeJF4PYTMQlwDzhYIb3BM9VjEVB2TCkwQASYDKG9/rsEJCtakhgBNL
rrc65g12aak9NUAFxPSAWd1lgCOe1rOwNloKu39ecbMr4ToXx78ygTz3MgtmRhSEZ4caJUYSCKHu
Ze3hqo9K5qyrNXTzTx5lIko1S2SjPp/dhIWiLoraKPn5oAyLjUAoG76tqYuBYunIkzcxCHA0icZ6
9KHwjW870AV71SMxtUpkR6V3KuFaoHpy2STyXZJ7pJOOYBzMU1zhhfkmFBuFDGmKjwDb11GW2rkv
mIvcjWSr3vDkFtbeTve3T/JRt0K17db/Idmy5n//nIjYfeM7BR0FpwpyiU1l70XM+h+6hAvq6cb7
SqBsmK5i3xT+S6nlRk6/N6e/AhbKlPbScXCfsIAkpD8pfQ2ewxkyc/9KsKmqmD5vO35TaJqOUOZ8
H6c/FxLgUN2FKqb4gvBQag8Jiq3O61TBhVc5YpRGw/cpta6oxOIz+ed4F+4w9mviatTYi6fAOmAt
UGyrE78n6EREDRi0TqE21Ft+CwT7v4tHZz7oqxcsAGEGngQb/5OLD1MCdJ1NpNPbVdJLgcVInEWH
KZyMPel2u8A46sa6Up7+nZkHLBJt6v1Imgh7pjQraWqmO+8DxpNaGkFGNpJP4JItSio1oH7lXZEl
roX5gDWsn+5dQXnFWDr5TNXL/GG3dVrzUWa4jEF4QRLTRD5HuSjIYyGli4KoewRsvM3kZvaoI3T4
PLorMwa9i1sO5HTOOZVVFo2miMz/7cC6nZwAbBC6EDNARQBFlrXhODV6MyzBz3RJKwRiMXWGZVoi
jf8OwGTJhEHvYXyv6XAYFBNC6B8T+3GT8kUHrylX8+0gaC/D+4yPzF9uHeQwuwJ50f2U7saRyDI6
1JVkHz3vL2JLO/E9jK3HjkG59MA2O70ibibm15kBm/vE6RVfkfS6AwjflW12dgUBriJkVXkOrN5V
90+VcLkE9XEP/iQBqPNR4PXnUrODWRCRI+wmc80nve7pfxwbKy9rqbKrmjJ78S4/qSWlkrERGJ0v
BTKi6iusdlHfjoJlgg5WvMRhMXpgbnLmPZc+OR4V3xZb+sIhOC9BhhOiJKNEQaMW4KmlALytEPnE
DP/0VmkH02ry+jRTSmurZMMWqETqT4WJwXEIsjaKQDxGK04hYApuukGkChQAIOePPoKmC90M2jxK
fcClpJDVxBJPTDWsR/BThtrW3CvxLmuzvm+yr0aQ2nk/peESTTfu3A/bTLtnzf+ugb0pnq5qs0s9
BD6AucWMX6RXn3BpJSrJx9oY/OEr6Y9Hvlqu6SQPataXiiMDBd0mD+7OhO/LkcNqaTxVe5HJpYyc
lCXCUo8JUPglRw477NdUMu+XrzX/gNXjyMbus8KvWDnCWv6oh/3VrCj/9ZyeefZ0TPfCiI0KqO4H
sDcQlPxfoLKcxiUrkcRJ2svR1n5bRp2xNpUstpS5higRjroj/ZW0SeWWSAM0DomOfCqsXrfNvhD0
+RgJHwnw3gem65kCJfeegm0v00Fb5/r8oivFfJF4k7Ui0LUG4lHwn9uoEFtwJU3AdGIlH4A/QLxL
x/2AiZ8VYnK4LUeHdXANW9wBn9vxrnWUQdjiuNMQxcvpKDSdHdgzxV6C7sANm9Okc40U7nvhnqEB
kiDFnXbV0uMq/JZYUhoozya8KoDld4LXin36WsfPumRm+oN3MPCyo0MzhjW+JvIhKaPE/l17WzCp
lB9tWM7YtyOhlB8Uhi7hcz4ie8w8apB5RHoRAfjdoFemo/n84BCYEbHOCVkwsk5Dl+RGnz5GrZlh
VsJZFSGYqE8iHORho1KIs0/Sni26NcTGqpGU3B1cdb9l3zhrJRP/YDQt3DtXzvLxD6M4Cbwhovqa
qfagZBejHfsxw3hD+UeMeimB38MOqEDbIVquxQBCe74MUbuftNidV4p4cCbsF8z3ubc/R3ANF2rk
h29yYzVXlTjFc9VdCyUxXZTxtQExh7irYvCEU5iy7HkTGDr+Jk8HJD7khqC5CVxBXrMt2w99Shvz
hXVfjnLqAnUt1QP7ZVY2sTMnu3lmW8RPy3nQIudWldyLkW3/YAQh/yVMOASAnmCjmoQ7bZ1BHnhd
F7K703J2NncZI1zrKC1LB50vMNEJvk+vpKDf4ou7+4i6e3FiRpp3TnaagAaRZ4Nz9JHkxeh7ZN+S
Q8XXAp8LEe60NDAM/70UVinb6UNDFFObMK2DdgSabLKDW2dtmJ2rU75SUSgr72aa4szymfSk83mz
zZP/Iz8OjR090zh6r1+kXoCdy0bObXwkjzgfZJQQr1V1Hh3tqY4BMaSuSctT0FnP2jF8fBXIW8a1
20z1Pdi4PkySU9zvhUSp+iwfdywzClEjXVGER4l0SlAYJHYGBcCGTqA4TAv2BI6dfSbMDCjW1K+d
zrBhXPJiIyVGaLT9LV8ZydiL3LsZidi7FY9r+aNlmVZAgdMXupzlfh2mOVi879ZEhEFBiIZMJXW9
Fm/ePTA2JmqTgnDqI6vEF30Oa4f5sCm2ezx2lkfwpeG27BvupzrDbT/p42bNscKs4/eyVHNuBnJI
8UHq9HMTA9qokwhF6wvsoIgwFHRCd37m1P71scIogvQYPQrp0J+TuIDwGENTi638dFoYeXtpAsko
S109X/d8GQB56tPdV1gD3NyzlYjKlpiX9K5j/ei9SLh87z7GCTpzy4048CprDodFdZW1X+tnFQ5a
oUf7zXthxLA6YRyOXwBVc1YIZJIYpzSiyYfhnAyYAPqy2fxlBqT4yH7htwbrqI8NaNK3f7jPfebP
w/IGwPe/iwEd15AQ1JV6vVnD+9XIIrVz9u0jHEC++Zaj1XcryUZcjC6ApbaToos1jf8bAsBiPQTD
2MMGji+rGJnbCTCaZFeSQpOkNu7L+mWqiE3RwcrWlRMJCewokTQt2nSi4thC9TelTDtHxY1BRyfr
2y5/kRAHcLQcxWR8Ze5cVFMCDr4qmXQ74LUDQe4XPDLBc/K9esnHIpHimhl+CnzL4rlSpbGDRTnA
AatL2DsFJGyOjC1cV5trVJxNi2xrrhUIMZzeEiAnWlYXCnU837gOrLQrVG8IXMzainsInQttDdFB
NvhvmE7QqeWP3mp34gOirvhxGCqE7fR+tJbDQLFlGh1Gme/wmS8SpcBk4rTgYSCAOR10DQwn1oFf
X+kIGy1gp2Vc64UFtWI0dGlFNqybWxgvoScgJbUieFvPNE/hSry/wo/ckqGqT6G3KRWFVI2JB+cF
ho5plkIdnq4iXR+KBRkT64+k3LEwVSHZ9JaOdg8akcqBydUXx7rYXvG4c82yOAQFz5pYx/o2foBR
uze9SHLAuD3cIKwXd2IBv0Ds77mEXl8znxfLLhsuRs/7EM7K8qKuqJMY7El6p4KBBwQcY68sq7DA
MOTqbUH7J7PZfKvTUUtbgDPRn4xSZiJTe26aMXY8vzuWfMuTv5h/sK0qKW2A3lfaSkeBr3kikrHu
sY/R4oult7yaA786Wm7jc8ffdxlhRC8B4Op3B9MQ3S4pX6tNzbq+BLl96t5DJTg2WdzAIeYFJqSj
4RlsP8TCeOhRcpd5C7cm1GaGGkec4FwgZJocqlKfAi8UWKKbg5auqBKsShiTAep71yxZHKg93n8l
kraCBkF6wSOu3kb2NR26voA/YskXiv1haM1IPnaDxMfF2bSZAl0uUsh9d2TvLfAkIQ2iD4EI9eDK
gpWrPB1pW+bkyqWm+Ixqt82u4EfGqJK/C9yZp7nb6U61LNlsg8Sjh8lzAwZ0hSswri4kYau8X2YE
MFIY+eb8nLZJqWoE46Kz0oMM1tWPO24CbWEWknqsQN+Qy3g+kkENTduFqe+g87Tp24e+eq/9ZcyE
6h+i4RBSu/fOl4nDeL+hVMMYr0s7uwuQbFTVcZftfx/boty7JrhiIpgroUPa7KlwQMCCHJF9OzQc
UGk++MlRSuXd+TZGTQnNzATdjmjRVeByH6DArDqFZR5JRoTUenBWJgsQsk2d2a93S1wMbV5K5iT1
+1j7wceqkLMGtF659Ipemlfg3fL5n+aKO+Tss622T14v4NFXS8Jcu7w3AsFg9OCWnL2PnMNTOA3W
uGhQ3rLGXs9wXwZXF2cpMbRNgaw3ea3wr2sM8PjqJsCXTtiMwlJjFtagGmfLa/nsO6Ua/wCDzMnR
wtyBaGaVPPmvvpQ7941v7hfAfhiaNqGVCEHtBTO8A85IH/U97JwyOz3v+a5hb1kNK25YKq8Atf/f
Xy7dQjCFqYDvy6vdkAZGFQJXlFlvh7MCGIGH1zSPgmf2WGhxNzJD0K4JJZRHRQJiqeP2OynJ5Bs7
vFHSGhlHTLMWNecG1EX76qfPGyyL7HFC3CSI/CxJdYlO52sEQqVPcgXcYaqhFEDnDsguuPCl9NDm
eEpzqYZFAAKuiypnbT+W0r4AXbb5enTs/32myMXfLnJNU34QAN8c1rX3TUFcD+4AGXPqFddyON15
7oCqgPabXOgzNxK7VwS+GXARPdX5EwBG/xkeKI39a0wq6jE0ZOxaQ8AsQ8CgP16P4dGrpQr/qz6b
osUsj5b4bsa1sr7pRxOH1p9wP50ekq2vnWl2uaSvRkrIg4Vm02SODN899RJoQ4AVYBKs5RPucLF7
N6tAE7GVAWruAcsgnjxz5zkD3LA0RNW/OQzXZlY4z66o4V3faSpsHxq7TVbBT2DfxwcA0TfDuZe/
zMBP3f1HIV4tdgg740YHY+y95Z4J0MGQSI9o8rDvFOc4H5go83wx20QCaWfR0v/p+5ZtUnahqhwa
YQjqd8SmVbOWqXQn3ShdCw4Xa1sO+CffuebbiWybFPCIUSo35uholQ6YOfqhnwRlnoJSbTIGGRwY
zZkY3MNpX1NKUBp0Qx9bCm79Dwoo8m2laUgTKKMAnVHHqqWAa+rKQ+3OLKxbJh4zJ56ltTQZ4hfi
iLoHJ1DvsY1Zzk3H7SCsC7zlj/tM1NvCRBmAvLUg0KgmZxap+Voej92I51DEG1jHZpZv2nHVOfvl
5BawTmdVX6TtVWD7+kcA/9E0LMfYONPR+K1vATwOlBOf5W/ZIjPvFe3o2U1OGX4CwDhOvSD+92Ax
f1TFDInC3OvO5ybajXL9uiWB2562Fa/vDwYv5LX5CWs8fc8DIPKFbayPmFnfLABviOgRLe4iv5L1
TCmB22mB8vNYwjJGOgV0FmuIKQWJa9J0hyzoFolfSAY4ppgoyM8EEOQpiLmlpdqqrrMqLm5FjOM8
bwGqiKC22hm0KdtyAWHUCoTYN1idJqjwD22gyZnjD+oe1Z4OJ8jFdfrrNyvoEJLgzt93UbYLYIeJ
KItpJHOs/B8bpInDmoRiDeMB113zCKAIE5heH0k2ibY3zwStv0hov+vlOCjN9Wvp+KyNC7bIJueC
6ed+dpKqHylXGJpskJtYULTLzxMxDiYlAQBIGSYWBc9H3E502eQ/WcJ9U1awITPkb74/oScdUi2D
aUK+3KgFQB7bOlOU/yOQ1GNLUo8kD4w/2RXhiMHX87tZ7Qzvi2vKdqr/2rhQG/sxuGtTWC8hpDZp
DxTMHMJACF/tgeUz5fvEfk/TLsz5ybzcfn9k/bIqRChrs9y281s+srCxolNq79eaRX4JJ9/8ReRN
P11Aj7+SDUsEO1hcF/1zCbbIU6yVUZwi+oGyWMpLMGl2fKNQRwOdqv+xMXWjzTdBaWL9RZifw6lz
LauW9n4PecgT1vUtWHNjwqS7sRlmGU7OKv4hvizCrK/ByEmKilTGG0hZmWtH/mhWLLZa6yQYIcTO
NM+4MUNbevUseb26CsbIZupYWS3IDC/7DvNRslcXZ7UhVHTTrY+PrUdIWu7p/7+ugroZfFGXu1q2
7ukXv5G7NdCSfl00StWQqD2hepFscjQETnxsC94BLDzVuPTlHZQr0paqBfa8MZ7raEQ3oGRZT/AX
YjHGHw/6BpZwENlG8RhDacILcMWvCKIqhkjOYMkL5ZdVgsvCJQhKHPuD0jByH7uPDMS6bz7JJB+I
x5S712sSqL3r1eFABZ/RSUpNyDGAIGHPAbQ42xqMKx48U+Cwv0hgP9DQqvS0Q85G68uRG3pPyFpr
cxx55RdhpN2nD0kHLHlyZZkTOX3uRNHv3xgh65AowfLZAxw5nK32mQ4iKqjO7kv9OaMwVewweJq4
HnpmaZhf7Y5rshfgq0xswhsZvodX2J20hinu8I7Bbyy34dGlf7/t+35/XZ2Rd/G4857acQ0RAn/+
The74SqOgW5N7tA37mo3XzvpaXXW8YQqm4lU4cso/rrgtxhMwC1iXy+tElHHosB4vIqFTqVQJ3qu
LFTTDI3Ck7XZ4GI+Q7DGJSg3y1Oukw0xUMhyEEeLXCgjJZVF9nitijTZ3lWpmu3l1yTCd5HxgyuO
C+vloIwq7VJp1tXlvrKSAJuy2KXOXGXaHFN75XUgLmcQKlD7uvbnsYo8p115LoaV5E/pd69g0E/P
lV+2BtEb5kEoMDu7E5U80e587qjdcwpXf/gZ2lZRVHGZyry59DhVzZ2ajmJ1tP+YbKnF3mmPH1cG
SOi6VQcR6MsGqLX9bXyB8NN2gixQB1pjF71RC3Pl1S/ifxCLYlXomPgWp6datBCszz9ZE1dL6KBA
QK+AzGe6ZmjRUOR3QSznqUpKOquPCFpd3ul0UxIb/8oRZbnosOoaeZpyRSG1osZCsUijMxDz/HRE
oL9O7jNT25TV0XK3fjdgNZoVgO0h2/+Ev+RTAl9nKCqVuhJallSeYfA4YNiFKKMmbv23XGHxv2i7
A0EpqsLz8eLd01nJCDU50gYH44LukKvBv18tL6SHyVJxMfcosfwo4PHa/P+G33SuVI01PtTRPMHH
qPbLV3ZNNWFzZdlDiLKNjQW8dUw4Bt4+Zbn3bQvAL9345L7LMRhoVnREfDZs/IH560mTxCBbe7L8
sHkjOyO5BLGwkU72z8E7ZMUAJrfaDy+H9iCt4HovjJ3XqY/zRPNWyZw7oqcNZzGzK55udnq9+uAI
JG4bT4HeKX3ngbZ6jBqlTH10NPcpu89XlVWCdR4814xRb6Iemv0Y3JaYdYeE+4XzQVyAPH2hvPMq
2nVsZPj/kCg/MGS947Xej6XcFcO1c7QZA1pyYvEdt4MDgUHz7QVZK574EoNx70Pgk74K0ay67OOQ
HWIktL4GVhwfC7PQ94xhgoLqc4Vr7Q0V0RvyZx5NAqugnnzg7XdCDHll+BaH3wSWLSHignS0Bil9
GKaWgHKVkPLXWCHZshgOutbYuQjsxIkSE+Mleatbn/2wM+5ktcCnWdVWX0ZTUVICptxh4iRZOB31
70bVxc46D0ObtEdMWj3LAaMetwNM8BlduOlNzKYgpLL9H1SWsHELSZHQillyS5/f8GfoAlBjEjCl
1sBwJzxV4hD/NGu9SydMSKCzxbf6ezoo2l+eJni+kf8YkObZLNnDcw17MVohoGUOQz7dAD2YDyfL
O2lGsp/UqaoHv3CEN8FXXOQYcmD4OW8kWBHiuF7l+eb3v4apYqfoRRVE9pIUsBAoGsa1Dp/2ktJI
rhPAn4RKtP1GVO0qzY9CXEsD6TOy9UlCaOrAANqN52hN+NiVkUW74/4NADO6mJe7LSvvK6Nec6xf
GQUxJU9CVBLLSlq2VP9riK5rfQ9S4LHn/9NRLdxVB+JzapLn5mByfdmeaEB4vYaZbcB7ssS85wsX
7Oss5VgOXezfiehYDoKgXOuVSQLgGxBbX/ezMIcck7UIsH0WT8VRX18Ul1hrOQvy2J06JVedkozB
HHdkNspOA1hxFXX6sJDwVz0itj7wiab/qcIpLHFvG5+lZ9S/DUjr7aYcflmh0cmGfztslArOLHLW
EuJj4yVlDajUgqkEK1VzBU4Jj9DkwgIRHhXptvJxm32MzUPTdyEhIai8it6WbNUNxpRK2gPVbcNv
WpBhoELIc2pJgbhFxbI5q5DVkFkCIqcWLHGd6p2shCX3eBf8grZjADcLBLYVv3+fyvgMghM5KB55
MBDVbXltRbMMMnfFKJdqdyKrFNtHDZJq5Vlg9SdteXvLc8zZId/2D0aY3jtw4Lg5B871UmmfOiS/
0tyQVzRLIx8VVd1WMewgk8MDOEKKDc2cLjulvWCC+hD9ksZVns8knU4ISqw3ieW7XEW2dQeGcMtG
rZhy+86OCEs7sz1Z0PB2SDg0HQZ/MV9zIYAdxrhvwd65EFWBpcYSl0FUpsnSUFgsreSeBidg1lRQ
ZsZEeH5x6Ip5JBwfBCKy9v+F5byQyN2L6/VtC8RdEb56W6ohU1zHVifJHUc3Thp+1bL7KNpJYyS/
pfJib+iWFofPJjQ08VoZIO2nNsB+dBpQh99bpBPrM+XIL38Fb6dnWXqGVdYyAXsOBfLfnbMvtBYd
dfbfmy2j6j6aGQN+2V5RuDywuPEBccGIhEbuK2JVEOAAdEMHDP5VEq/Kem0tXP76dqkX5ZBOI2ll
UkfExLVVcHtzrw8djDMdx57Wkw8fuk8wIZvoCpZghMQOmHZRkRkPeN2/v/5QJ9phfzS4pGEhOWx7
J20VdmtnbYMl0XRDeLghFTrqDRyItggh6FNaAt6jcmVXLc3jzRG7GpDC/0TKq3SuP6DUxO3wC3G4
o9Mco+7Jo5Xa004ET5PXspZDctKlMSm83P9FJYbZLME7is0wkqjBrC3e+dTuCpSblu1heylc4+QX
bENTD9kJr//yrwyCrg+SHTtYcEMleMLHv9f4cPo24pk0bZaEGlH+VstjdJiSOP9g3oS4RphBN5yY
SAH1CFnpbPm9ZSalgiOl9ec8TRNRb/YiGk3SPYxt0dXHN+5sD0midkcQ31zwMx0ZRA1FNpNNLuyw
nR69oBkh7UkY84om5HdIDarUo2OS/gLVllYW4j73rmqVA437VXjNemV4QhWPm/jk9LKacatH+8Cu
umsmIOic5x4VkI7U91rMZzVH6H8PyRDlrhYmm0vzr7bfxyeX8ofEWlY69IiRCsK96a7AdiN0zNa7
27vsIBz1z/CnLpG3kPVkR/ZV6xcY9RzNK7dm2I+jbaoX2Y5JSLOhDzhaoBagRyZQ7hZSZ1M4hZbn
R+/CtjMUOQWBu89oXgXlw+V5WtKJ5+o9jOztBo+Di5cv5ZJQMgb9radiASjVcth/DGUGd7EoHBuX
XEqyi4fUhP1KphjqBuK92RenT95V+xqdmyQhYR5MtE7HBKd2m7PF2JQbArggzczjeresHFrjQRe5
gdkUoyQcZzq+lpM3kY/SzyEoOzYaRSBHM8oaQsdnJROWKQJ9ZRsPYPTcRbIlVzkjMOxhU/tSvJs8
BZqYWBMLoME8N741E7EgZNX/U1aTe1wRiZPfduDy3e1HbN2LcrKUbHQOuTJzfnSD6wa/yuzPV/Vh
QhAVjqA7qeD9aI7WTZkC6Egxwg0xROI3m5cNDnyDk5kX3qSTSVANRYjfV65gy+8NBh0KioT28ZV0
nx2g/Qq8ZskL+8R/Cc8FRIHFPvH82eOOBgMYtUUzBSY7HUv43BEa1UgG+Y71lPTDY+K4AdBDQ/Yd
LcsAXjKvI6LYBEk3yVjKHSizwVA9EDiS8FrBC1rxqJBV7QjMLaRwjRIZk/WmZgf39INTzGxcH1zy
v26+ejWsdCq0pzL2dleuKtQlaGZ6ztgCXKtQxQocXPdFP7atZAO1a84yO07qIevrDxWZ1tXLsTJc
8ZWx90MV4fU+w3TkwSDLnfg2WmpQ3E2xOKRqqIrk/D9Mt+K2aEF0kaeG0kCkFz9GoDU1My1JXmse
V1e2FURxAVxRGxBdzyvVSAvSnloTOXBP8WrRkM6BcsrmI55NkZ63bOyVqoOYgbtdd/EkwsqOYzE4
bo2oW7PMnGGDGYEsaGHGwme1xRXDwoxmBW4vqQ/4VnyJQrHbQY7hhbhXOvQtF6SEIl0YWUysLc3c
tKZHvedEPCI9s+QZ4mdc5SDeBVxofB2JxI0ZNqT3kPwwi/zgA3ScY6v1leJNEOdDTiWvpPz2fDly
GMESJIfizgbVUjZRS+jhtsurDImyq9Om8wU7ap3CZO20WPgw16cHg4O9vENiCAr3Q/YSL5f8OoK9
UqK0L05MmDOIfhdptWFXljLiG8lXOhpvuGNqJI+vhCatPPgbEuyz4te5PU6fvjN4FTWeGpU9FvQN
XfxFo5FSDIMjMRcijHvAUh/uC9IWStBkkjBJZjsiRWxHH0WdhBrv2VtU+wYTPkYQUz0aZOet1OMQ
0bkXuYx1ZSJ1LE2zFhUjQax6TECKNpQMrftCbqi+OZYGQEdoUj4zJ924QIm2f2KLiocTX2LXxc29
IWnzC0KvvfGbHw9/X/4/P39qhyUEJ547vg8swA/qLzCyUWFHbJGGFb+860k6SIS7hBOB6pwMDP2D
Y1yaHJ742OoCVJGvbvr7EjAF3fpxeDQpbF6FqLqEGWQ05xtA9I+wcF9r/1qyH70rIhU0qsliOCWI
xV+QrEswE2g42rezbbJI5znSGw0AQ7oNOiMFlw8hQ3RBZzMBq0xx9WhJ7sw+MJCW1MhnGvgDm5FJ
qa6Saro2r0CXoHsKrJRFGwrBuiAiQXGntEP76ZE6nL4aSrPI1ZPutRq6TQw2vzzfq0OmwslAmbrq
zNp1GUHqyn6gShXzgp5HBBzzJ24JLBnSV4GcCgYSDGqiROJQh7/OQDN5hTk7MuKfKDcvSOyQKImj
zVahUbIRduXtM6acosepQ7X5bOfWM4mibrbbiqSbu50dg6mnRDCsyeWaSzxDLcJervmdR01P7ggw
zA5EfeNtF4kXOm5VmBCEPonD9C0BzIZId7cSntUFateNheCgi+k7HWFalWXqjTz9jRTikbALYSgQ
nX+O0AGXuAsR7hW0zvOGZWoFWpz1fAD6x0T4i0W24bnQyMjxIehZkdfshus9oxgEed4+iZ0RfGzU
boQy8XwB8WJ6qbhDZPHluU+MKnYfsvaP7X6BxjrafXoEXsx5Eh/b7eGneAEHjhwBaBpAKNp+YK/x
huZWE0kZow+zzdosDhZj1IoJCehhivVdJWbWvjdZd84TClFW6kRWrtNhTkgXxlXZdjDnn0QqO7qk
hGuPSF3QKSe3sfQsGuyyVCsL2SHD7mGheUKuS+53g80EEE4q1eaOLFFHVSUpqTUv03JJOAzZhHEW
H6flXW1kXiaMUdYGy9VjZtYukHZwSVljmxRuzE13yA7qrlYwYsEuqjE22O/sbDD2rsnjl6qH8daN
LoNw/PAsvzZJgOYD9vwWROU125B7ou7woq0by0KVJbwTVaY7nbx0nR/TrPXsU+SKt2miNHK4rDko
0GBLUvdmwCQJSwtslc7lmR0PrQEluqpOAC1SLERpxG67Vkl+zT+r8Ub0f89y2uD3DxIv0EdKs97U
bmnzdOLbvNPm+ZYjNJ6w+ak+vXrBD8jdMIsHFfYsvPsX8ZDDEt4wVTDgIv1IiSk1fU3SwFhoJn2M
mELNkZnaucXPELZEW2tkq2ldURQJY/GRnS/BxNzr3Pfq5m43twCYyYA2RjCL9n+6moc6R9moyaYG
KDaBGl4GVOkrPx7CnLCOgNWd+OuCc8RCojR/ygvEcEfY+ESdeOjY5pR/LuvDl02/zG6xot88xWOq
O6QbEDoI4PTGZoci2d1TqUEDZJ2w6s+Bhv1bL9HpmerweA5fOcadEntABjKprn0zxbRn+f+pdQxn
1Uv1eYA9y9scm8kZPf0iF0s6cRvppFhNIhXU+CCcUpqQhV7bKP7fR5XqKtQQrqP2Eb+BxywKOHbL
ELkV+xsQ5aw7jg2wTax3hPxsM/hx96jXtwtBQgpEg4wx3SZBGQDLedQho2coS6vIvevZaoQ/liJA
+PhxZFnIqTYg2tu77WpuEgQ2PwUR32oKNpFpByVyT6oQTJzOta/y20P4y3/rKspeuggJ1Vhx8pR7
q05IYdxLw/v7R+Bpcct7SnVg9S2wR6XRFrzEXie9Zw9sz7b0w1Pti2JdtOKkeJcyNEveYhjK7VWR
sF8Vi3fl4LVdGbGxeZssdEjdVvmVsv11Sc9j6zct8pXfnqC1IsxiKMLUCEoMX1P8YrBj4KBIAquO
U0o5P5QQaGrksZ8uqBcZVv1RF5E3txUaQ9EppyVhOBpYe9F/SjqOS/2q5xcRFBTDkEMGvBGabcqv
iGzvCyGe4tA/tSouO/kdX98lWkk9N3g5KmcnTJBTqJSB+MFbDKYaeUlfN2sCb7EGE6oPpx+gTYYN
yYfu1WpiV8sSTkP3jLYfMLSPlMFs8QK8YMhDi+Q0t/+KEAjYe9vSpu3sCsly43R0DlHuYPlFOu/I
yaBLnszgGyjo9X2k5mvfPCu9yoNGvlDyh5sx/tioujtLfXo2fx+XW+9WvkzmaF6vhVzjk587tGNe
VVaraViQCfQI7r8tBPfReRgWSI2HjxMcBwbI8VtR59lIJXZzD/PyDkr9Ez5AcB6v+9lAR2jPQo9i
FJJizcqXhKFRtAcb2O78993ixdDWvZOwgE6nHt/C+hpOhQiAjWZv+1rCYJ9LNoHWAMUPVXmibSOO
HO2661W9mA+EuJYOFUqeyQOAUpWFw3SXGUFo9UpLzzpBTawOpNvzefXSZdNyOaVh9ghwbrS8Mb/d
zVjpe0QQVNWsuN2f/g7PuYXTvrLBtw2Gcm04SdbDZssA17pnRafgEVQWE3XbNQFAAZC01iqXPzWi
i+BQjV38v/3Rn+L8PS5cTyRgr0afb7DAAZAypa4C6Cxh0F0OOet0jF6oPOffrEr8EmJAkkYmYPjj
847KL80Nw5z6Qeez4O0rO6pAUGCSFzPmSAAj3T8stBEL+ZyZjo9vKz6ww/Sk0KNTzIF+lSQzl863
+v09cZ1+dTy94jCq4hLkhS1wruT4scU85yYo7fkOXdG5vNgJJnw6pTaWi6TTPOqfrR76bTA6v23T
Q4kzA3pZa4JvwNiUW0EK6Adkt8+CpvDgNR9JyivHlH1rRxapOTNZc0KcdrBDEGCzu8KeKS9yvaQa
eQfAJVNgEoGKuwzOx30+1ER4sONtY3T+7NOh9pC3j+F57mJ0b2WA9e2WQGoS6qnteH3Vx5yHlt+G
AEsOs1uVAp6PLhf9d6zoZ8zY8RMOcaCHeepLTLaRSSunFNbYH7w5AXiLiuVNntOX4W/+8Ub1lLi6
2+1L6G8MLP2Gw23nlWlgSlODPH5hKnk/tk9ycHREs4bI7/0y+xn6MisCbkuxiBIXdJ1dYowAtEJf
LkBb1qLXTPRzfWPlzBo0hWl+9UKPehJCWtaaAVzaW3MeYSPF9mR13AGQXdBWzyDcDVJ3TkM+eC/d
Lqz1nFAPMVk5v72aKxZa+S42e+aYysD4IRo3CQqdEcBkbYypO262cab2kRfKahx37dj78nyeg3ur
s6Kc86gpiEwgx1kCglKZrWuPLuEE2xEF3fq/d4E4zX920RGiUCq0bAPlKPYXiiTcsZQvkX2P4HFD
RgVflfSXCn84GDnk3gP+EL+d4Rhhr27oNQjnBVmWtwWsbje34tElqvsGYGXfKR/NUlji+El2283E
FsqctXai4afNIR/On+3Yo87jweNY7345Yu4OOYRkza3rykXRoZKB0uIUrE5n4jTDqfNQCiv4ocLq
LhDqVBWr09UqCDuxJma/WAfWDNcYoIILsUAYTiaa9KLiUrOKLEMOBC2KVok/V6dRbscJpMPZG2hA
xORegRxxIMX0C5PiIQm530NYDykhr1XRU93nk8nXr4RV///yiKW48/bVX0cPMXih1kuhFZqonT4g
I7hU+k3He/HCWt4nvYYmiyRUIw0mIEMaxyFDjc5iILYxmbGttRboc76xfqbO2ah88dajIMH6e4M0
4JWLMLGsx3Fg6wyr01XTDS8vt+pazX6+lSOGmOoOvVmV42oWOlGLDR2Pk/ew6NdhZviZVhz4AhYs
JALcCaHSdk7xBA69lulipveGwZgbBmdK4L/3gEkJYZT+L7X2PIvbaBBabhE7wm1uYw/XbxO/RMnF
YvH3vJ/62ohmNcrYfQcgfjWfeHKzgNq7azt+lw+ihIsYVH8ixjdMrc621GsuXjPdMasEyD+CX5UI
uYBhxJbnAsZw5E/6ck0XoqjTt69Ez+9op6nL/D3lwUVSNHr3NsSk8jKdur+uU+t7rJ4TxjIi7zlR
eG11HJejWA5fwWW/PPfWoGG0noKdE8B/7yGGJ2oXAnJN7ZElRbpSUnq85HyI+oOW6z0Hr0xFJmo0
7bC7MbF3LXPomWWXDvFB+2ka2wXmzFIvADZ6lGeGCI6BF70qRCEBABNnO3SWlAYDpcGghydBi7ws
hYKYFbeYGgn5Ooy047GKqcMEZrmidg8KDkQ/k2IQnfa7EvKydCguSYQLpYpo1A9haOme8YkirVWC
LIYjvu37/M+gEKnekD6YpWmiofes7MlJvCPLWaU3xPswJS/mYKX2lV6/UzniRHHqtltHSIy9Rsuo
9jic97AP10ef59t0S9Q9KB/3r3EZky5f7mz3vHk1UkvfHiuifJf3Vrorb6Fi5tMapj8lvL6IXdvi
jn/o0UatFkzxQIPXK1zrRniL43XURe6rNxZ3X4s/i6efLjIqmyzoWJVlBJYtFBXgkRccO8rjhVbt
kc15z+p1S9ygWvsYt7DwTQqOp5i2eVlu1qPc78131DEw+yrT9Qa+ztWnx3URW+BbvEobArFoAEpu
bnqmVizV6kM0s35/kjxs2a7cTT31zSqTuMSue6Fxph0IrLDgdZnJwRhnMKAC+NxngacVTKGtaSQ8
E7JOOtQw1v2yfEjqaqSHE1L3b5z6yZA2Wba6mBXf6nBsdyThq8QwAIaFWSJz7kokot4gujzqJ6lG
FnY9O8fscIYCmTYFGI75MTJpEEt/I6lqfkkbQCsGswIyY1jEqTTV7C3Uu27XxSmBztROxVkauTDt
JV3guvNGQHylPl+rBmNZys8tpYdpmKOPd+VGEuNceVwcsutflP8dKOk2drfnX786dccno5H0N+Dd
cTdAjTcl5UjnOoDqgCor1RN/nG8BxvDSF+G/KhYLlCK5awPeEyscpEgfFF01JOxSRcb8m8xt3hep
U5aO7TahOciD1c3jQ+ON4diQMHd0G9usBDlK8SJny6I7MP7hqlf/jRGTfrZtAQ1gvjBLwMUbbVIk
oZ47OxVIbeIqPmjM+rydT1gDNCaYxCjro5EEx/mLeOhYnAFzXYbaOAsMxicrcQyZoyR9wH81QcCe
LFlisj+Tg94cEZia3F7Co8FHIsShoxB+KeJP1qgG7YLCoD50KDMOcinwI4W3hFqwxqA1RHGGG6Xa
l67dk6zDUPvas+49iaSc4fB82gLttVMakaZN08olAsXtn0WCmMzTBOnYtfRM26eWiEjA9vNZNqBO
paIu5iGjj035t08r9dgcThnRr/qwq6qPiLzi4HgC3jiIZ4gz2aAGw6kJWdXBpR+UtVzyPnBgnDlH
ar3tFPC3jOUSrqm/+EOYa4/fkbeO7MRl4Wtm1LwoA/unwhP5TZzbuDqf/HywDOZ1nl7nML90byfi
d9V/UsB3h13xbKeWb6LQ7V1mCCTZkg4oE4lCfdSkI0SxdksH3irWuKoFNTuVeG9pbjan5erqiFH8
GHe/rV27ayNxL9G1Sjt0eVzbVDexxszGslfvTXyxbOEuRTfvWiR0PEFuilhPEyMEvhniWohhdnjY
ojrUxZbY2LRUubQ/Si4Jjulg1ln5Bfb6QctF6Bi7fIF2f2fPHRhH5AbIaF5Th9pISFprj5FQJncp
zEMFcthUtTtOdYCk/0QG+e9mdjDqJcyaG4wPYb0Q8VhEmGvwu0y++sSW9uHks6Bq3hRanpo7qEzP
6JqKc4GFJjXqyUWU7LTS5Y4NKiNbdDyuAp5VQf5qeoaU9hDjVDWbz+kY0+MjM+2w4+kQHJyBN4+W
bI4F9EG32+KUqpsA5EJKqviVOKIXD8qVbp4xqS+l4DwMiAuwIfy10kDYwoD7KSRWf+i40mXuC5jm
Vu56f88xXcmHwWLUWVSbtBi03WJwp5NyIS8YTJLTZeMRWW1nnxKtGqOi2OYsFaOURVm5qVaQ//zj
+Ce3JK5aGcaZVaoG/RsAKsgp/ZCbsBKowiECvrxxNEbob+jF1erSQne7iDFYatgWnSNvtkUNn7F9
TSlq/N56lql0lh2/Esw2VE7CQ/DmyenRu8khL1AGg9IXfAn6xRRRA7ZHRxVP5x84wVH/nF/3Fxg3
v50dbmcRji68QdVKTYia6QpBXDebfmte5TGdlIuWeo/OSckV+Xyon1ZC/VDxbCLkI4LdNRoRIMwQ
fJYm2HMRV93O3rdUyCx4pYodxrAji6FUQxzZB52PC70BcJzqkLmsX7nt4eFQBfpxy2ujmMv3qcvP
o+7JHjfUGoRkzNgw/P8kKn4/qjYBccEJXxn5dPNgpYf2S9DpHmlaI/JK3Oods2RZQCLrS2i4/HAr
zim3NZRDhvntU7GFfnGIreUT4Cdnfv170o0+bYBuONWTyfUVx1dm9LuK6Mp7jr+cVRl5Q45fuPEo
M9yhbcNHBFRboAA8JwgFXZZO7SfcJptYCwszGPnPuZhh4HBlYuxLpar5buakJRhhm3sjKnJBEOHT
zkN8dUuuCm0IPJXAS4xhU74NOCFvPvZmmtlWQhdQRDz+rpxtfC4wDpT5eTAMivDdj//C6IlVdkCg
6v5DKaZRXgX8CTKryXfr1dx9sYAoPzhXsoqvMGfY1qfUpGHJ/fwPhPazo1Pg3WgN9vioF4Q7DVQU
I/y+stWZzgmYB9h63SEZwzN78TMnulo1XLv91HRcn9B9uQIlQH935j1ONFGrpduRTrgZu4Yin5S0
u+rQQxpzgCgUNdhzLr21TVtSDuIwPnBmoH2yKl0cnm/1UQGnoMgtnJQAyFLZkDQlXbjugyloteSM
Tm1lZPCcj6Av9wT7dY+MlnixjiFcKYNTqU17qQBy44roPC9OEWglmrJy8Bo0o6baewR6sPQBdgfq
C7kizvWbO4LtGDnlBWq8eg/08lw3aCntkbWk5YOa4QyX3AnFyOx2p2B0d9zk9Pq+kqrysmuV74k8
cZu8GY89Lhz4l1rBKXc0HETK2//sCW9fJNfeLMH0yo1YuBWKBpdJ6FU13tnPtdhAuKbeZaE/mp31
A6XoLyQtNxr2gDl/EDMR0hX0ODPsxRiFSlvwIiS/pEaWRa8KvjyUjLzxkkrIyDZeyBB4q168A8qN
mYt5sXSI1p9jk6d1gFhahfahOIy3ZGXw2oGj2+F3ImBn0JOsmrqQn/aJJ2x0X5uOfy0tiEis/7dX
ohMwcQEHKY5SztUDc2W5KBWrRShgD8OaLJVbbZkuPZVb5vpVTOzpBxXXW1f+kX2vunN43lDlj8I6
mQ4b28OqIkLCSfqjGzJQCKpdbLa6YZoF4vVaV3/4KnoWInyR78J7PXWuX0AcZl+JvYQfGKyn5hNV
ltgDAntJqTwRjpUsn8rxMOTHlUEj1luqcz11/Se9jOo21hsvlwtsB4EW9ORJxalHVEgl/Icbcly9
FOAon58YTn2ddwQQrKsQ8uuheBwJex1aKh2z2nj4qhtEKB2G1s4k5Fewsh43jorO3CSjdMSAmZnV
TYFowHGiNGUUIxeAJh7pGU6gHR0lUnqlsSh799I9Q816vGDQt8a0XWGk7Bj/aSej6kVzz8CKhjeO
gsC3Cea7ceePWaDYmgj+VJRvy8S8LM0ZVtvnhi1Apa5GJOUmtOfXUMbnsdtaTBWiKVZ7OCqLtP8D
W/LbYSfWeJ02ukePAem7cDGOWdBpYj0rt2CdyAmTJ6He0vm4wuHh1aFQJW/bSBuc00Z8dv+trz3J
jSmfiwRKTiCft8HKTQxJLxMoTa3PGyQkdjAaiJ9BseYBxp5v3MT2Eb3hWXxmqtSAjLF6v9AKdEXf
SzBVyqo3bSNGKH/mosoI+6640t1Yh/7DyBFU/96fQ8A+AblE6/LshelktvRef6UAaazB56q7YZKn
n1bBA64FpGOzB0KdRAR8+ygbk/BBWhfjtmVJ4ZbF9jJq6zf6NJBMyEP9cayblGNODfucd6yB2LKP
bAY40sNCrhFvz98rcaM6Wu6tJ9B8IWe2wpqgvvscRRLJ1CrualGR/rHGSwWbU+5dY6zoqrP0DUNm
0vUnxi0byHoFvOS9R4FbVevN9fethNcvrTj1G1QZt+hMvHwFxStFacrTqj2P9wU4J0rrZv6LZggr
CfVt1pQoY3NPISfM1qYc8If6Y/z+Jqe/v06Zg2DjgeW950haiM9f/KcFcxx6XiuTZOQ6D3ZR8St8
b2OLLUxPx8F9o7H5dJVs2HGciIMg78EgGkvJlT+CuIhxtagMraC6MGZpLGcvnZulf1fMCCArmKCF
v/YAlqDPXXRySDmbJSzlixBznBaQCBNLrqWjKP/UvJcTNYEBD7F9fefPOdRWqOkGly/QrWZybHE7
CyPIKM3Sa2cZM/oDYOA06zC1okePcsvZkVmhqe4OMnvYhGNvbJU4WxbThYFVVxvYnfLDu+SqBQTf
jFCj4ZF+ZYcGYBpzAuHhMOjlVsmwFIi4IKvsT0xCaWTBGuSiKDbnWCSEQCDVDskst2ze0YCZ8VgK
ryUGLTZXx52Pe/C1QRdWCqBeenSo6Yi5/jAzroYijNX4or6KG+nYuvYDfL+TEpjErzkEvAWZofbH
qGUL+0D7OQQ9yc4p1WWEI96qgQwFCcN/CfJr1RtXw4Bxxzfjy9HavBNdXXm1B3Mj1forS4d8gI2B
noITAQPEhoJiVtVYsZxo2G847mQI/YtZiZjzmv502ekICO54VnZGpNfFHT+CW0AZzjl6jam88lGj
+U6SRwHcr71jqBcDohRqSoddV6ipXyNeRi9wfmwOkdEjB8fIoFFsyeIPCbEV1ELIlkRDuOeVVH/F
/PJ19Bi8iSL+lOZor+ZnIyX97UkEsKmeakNqN6+Qz8PLR2KldQxz7Ei0A8HyOklLdvgEKOFDleGC
KBpn3GS2E67tBs8YnjMUaVyUE0kb5ma3a73g4nBge9g3ICO78wYj5ZrB2p0O4ggRSeGzJ34UXxjb
RFdM4kKv/WUMN47vLU8LiYjoO37WFFaUzani90jOfpGTNi9Xb6TivEkZ5hWVEyXxb4La/EeCo7RZ
nShBVEhsDpYVi6b5tA8VTs82WGYltYvpVnNDUsgsMYYe2E5tpK02syZVi9fPgPf+DA0hngMBQJEy
pXtMDGYFnETQ4tfgvjHsfu1mdW6U/gprtDq4YaIAFa4Y4Fb8qJq7SR27r3Y2eseor1/JEOHFcqim
l+ut02Af2+/8+tfeGQHlAejY5Bqmt0clRAKxQv4RUNinswMvtW/ZFhLHRCj6eNkp1gFCc9OY/OFX
BWqUXP9oWaEkBkF7gwi3OLaV+QPOWOfEh+rzKQLHBKhx2Ru72jzGIOpUDYCtit2MkpR9EDrqBBeb
wS6avIduBWzZmB5yC8rVYdirVNzu2qwFbOg5acJnbnbvyaw8w5Bv2Rtcq7wyfJvvYRyWF3qTQUEI
VHsBBaq8FN6qQhQigoGAP/+mL1mmlAg8BiN953HvP54bdvQfy12/wlwrhUg3tkiUsWpsykslIlCf
rKXHKJW06g6v9WSSQuPVBA5M3LcDcwVDMYMUXd4v4Idoma8LIa2jiDj6UBvZfYPttrfBSoJTMts8
wVoXgU3KOBT4x3Dc8hD7mYfywK4hHEO8lehuXuNISzRwGALRHKKP/hSCaTipAvCmDztpYivbOVq5
N+eWLfcp3Tc2b27bgprB+Pl4ICR8oIHpeG08rmsLO1JhR2RPnmRKQajlG0qo7GcyoHt6c5aP8X2j
Lf23nh0yFWTAUU9Umcf+HbmDAU3jKLSIxgZrzq37a3NIv7MUYAokoOAq43y3q+oChiXlobNaygSZ
aYrfpf0TatEfuhMRFuDw96cQce7ndxgUMTGXHKQLmr4kanxVOG0AiS1JOnzXIhM4y9nQnHOoShRr
tMhAoZErBKVm6lD/fWf3203wjGGMOyWAK8J9zriZj5Xgt42i2lBmcbacPt/rge7nRCuZULpkeB32
lQ5HbXdcVBNSoCofjOM224XcVptQE4izHKgnCgWLuKbdeLWTW1lUZGjdT0zuFd40yIIkFs0xDMn8
7z4jUKABYpZAbrO+p+5J/3bmW8J+8x856NA9jGvfZfha02oPK3P+O/7xx5Tkl7ldk/ua+r62MvRB
DNpRbeYtm4GO9CsJUi6cohQ2YIEZt/FEQ6X3G52IJisvyZoax6rTGGUcm2mddYYoCcfOaK/bI3em
0+SN4CYiR21Hp08FbLQBjRv8upoaWQTHaVOH5JfgqTCYS03sRGao3f1I5OYZJXxrFBc7IJtA2Olb
ewzDEbnF+pB9iuF3ojXY8LL8Al4uylbNw6+zTYa0qLygQ/YNwbhBuVkWJypUbpsSRcyCxoJq9n9y
o8Az5zsgWe1TZCzxZlVPDHCNC+CJEjHAPgzmAWPhGiH3/UDZkY4w8+RUn9RS/ykVHd7ssfUd7taP
kf97K+fl+nFUPwyIwJ043BjvEjBdisUoS4+PmMhVWaIGozPTr0N+UnlHJGiACqxzXj5r9GGRh74u
QXAWw2SOSpdVA77LVQ5i6PxYTFSUVWLHTmleu6wKEqNm/7OG9pYLYaPf/p+98um+Zp70sccx9RqQ
4CBjLMt/C9DdeVQ3XGkovf85x/Xt+iGoV7x1FAl+pmS5Q0uXIu9SyTOPlh+ZqHkXX/Mn6xq97TS0
sZN6tLUPQdia5IrM8nm5qGkwnEjoJm7NIZqWQvsVa3MPR6jXQ0BKcQ8ShLvzZJigprRXWfn83mIq
+yfuttw5n19BBY6EDxV6JxBdewng9c4Nd8BHmCVtmTI8eSS8X31386ApboHw+GVrAbxnZcM3br4D
lrom+UJHc+fY9FnR8nZfH0prs8yThHqg8UKaBVWESzTAguK2jvA+UsZA9pdQLGC0rErQwA/Ehq+T
Wayl47PPTMJdJCmt3r0H4i8rLWtwQXTqz/yJsfBExwePU2kg3U3abQ2fw7t2CCR9QtgVEQJ8KYSc
PRpQMIUnMqndxFfqOzFJELkznndPIenfyzcUSL8M6hXgIBYc87JhUcwjcDEBTdm9iucdYeiDRB09
DGoN0Jv7SuJnayx091uvg30sJfbhY+1tzlF1dMXwIkfNsJqMIHWIdsAryjrOK7fSJI4be7bLQYq2
T5Snqb2UnWAtOj4pfKDUXC7YdTinXKHWYzAwv+qsfkurGsHjYDkuv8cVsfhI2rXH9CZlvMqvD/aO
LiLf9De70K1jv67MYd0dUfnE6kB0cNJZDgF1OZwMGzV7E9muZdduLSgRcgpJMLCBZHY2p3H7YWY0
9WOmSSRJDoVMm0xgQY6D3oSRHiHzUyMXIu6UB2aYnA0S1XMZxRKJti9SkhgDjFiK1TEdm59sK1YB
p5o41A4K33hkLpxtW3sepKfjRw6D6ZxlFtIAEecXhwybXbtAOd+WVHwrXOLMpY+/RSe6Z4bHhVgU
6/wDyeFl/1mcxi3E4PUCnIIrVwZf3CQaUvuqir5ahOFE6poZA3HorH50FpEAznsclKyOQWniTbbY
mO9d/dUtxiHBCaa7EcpVDCM3YMnf+A+GAnXE68n5KTx1uewTxL7pOvWfA6Iqb8DOEDfXNjnDkCYi
egx6fCMB2EWbYf1qmp4RYEmJAvqoDIO/RlXhtSTan/oU3QoLi1QWKSIklu8ZrkW6iqhVTIi0N/ze
/338LE+mxWVG89fyEkHHRjYf6EqrnBZod9JeAxeqKmSbiB7OqkjaXv2E+wxW2RJTcYceAjHnsU3o
Ggm6Ou9Sa0Z2fuFW4/lFFUCEzEW23T7HUK61qaTR3mTDVdBN2RES1FufFci0kWSndGtvi0+tuTbK
n2WPNzA0yNGMkKagGRxOtYirr496IgeWAlN6oXj5fsuYqGTYEPm2uqdOyB+Zw5jCQ0h78z/rzsvW
X663iTOzBl0VFvtlK1902bEJ2f5mwXz297VUho1VnCjTfbLJDBvZIDezDhOnF0+8ZQQKHCqbHzzI
nqHCVch+HYNALhiTPz/nuk+pwu+uoK8vB9WmgH2HfVK/ev/0UTB7O3P3ey+FtwryxZs9Ql2evuh0
MrruP/cttUh7PYaN9dHbSCmg33WFxPpb9R28HWOtynpdTf6an71W26sUBlRUn+iNef1wD8dzFZMf
1y65NZbfiNEvfwG3PE4AmqYxjNqPcNyKUdX4FM2YIha1cnbFY01bO1g6fwTbnkGqZd9vZ4zDqL/5
lCChRlv6Eqkxx2lrj5NtWDo23JnCt3h+hIXXx/5dcfZhkXKqKB82tbBVLhb7EJgoFRxnhVuGJtHe
uNPAF26bRA1QKO0Ivy2Mf/jJCXCiQlVodVPPaD/RSKtqJD2hnGac0nMKzvB3viRaA+OU7nq8lKYF
H7ITLZnHH5il2alNP7m0SaUKxcII/N6Fzdc6H/EyM5nPPFt5/iNvkqqSzOyiWvyl/HflAZp3cYT9
Z+assxk/7D4iXvKRc58/RnVIMWE2rKZ81vcQYumC7b53ypzldAlUREX3IyXgQqGiKGXCRIxmyUuA
8TEavtZ8soXIR90cu2bADZnkVaUe1NanGScHm2Ba1TAd/6uEdHEbINeZbDfuV9OCof8EiLp6810J
1ls7xagqYXMLBH8V3lN6UlmNSlDp5zecA4w4Z9zRFr+vbiVjIvuQjqn10nPiCRiMozePLpM7YRm/
HAilG7VqyE5t9qqnSrba0tpiCb6XSjR4sGLlg4W1USrgoL0cre8mjEq7OENvzQnYKlMQZe6AMa9+
UxQ11nVuxiLiBOsnwBg+mnSB0LQwjeiLjJwmQsSpuFCurJ2Zo0DetAZayXWW2si+xwma8HbQg9v8
BMovSWsJulO9yT7F0Anu5lvnNjopKgfQSY3uvSi4MvqsaQkDoS4hxRys6qRttG8dZsPG+ts899iA
9jMgmwc+ihQn00XjUpZW9cHikI0+y+TbGdZGge4K92VqL3+RARfyIwjn/z+ocEHl2onUAh+tyVFB
RwHTdMz0yhUr0o3FheSVvI5qIeninRTRsl5aDY+6X4izI8MSOtA36hlvn6DpuLVB2vt1AXEWtfbr
xvouxO4t2bDVly+SrzHGPLLRvmM6Js4jENAxXYvpB5onnjop0WMwXEe/g8/XECjVF1fpz2wjTLbX
5imqvy6BvOykbqWDMy5oYGgoZk06zWdWD93dkAfCkhsw2jHbLDSm2hMwvqQZT3x3T7gK1tvLJu1D
RzKe+woL61EkQGt1WPqeKNNC4wM6UP99kdnhxwsGQ/1EgY0ia6gjOlxrkZ9tmd4ZW8tt73VsNUAG
kQ3bJSx+PZgl2RuOzM4K+m0hIQBbOtxmOt/NCQ93p6dCXVicvYz5Y3d+SMpkixKSfKqjXd+yzPRD
ZNgk5xHgxj/zEo657+VIE9j1CBZeF2Sc/zUsm7gohneTkEy1imWwHoLJEea34XgBtSje6Nt1AFdN
uUxDheZyU4Tyt7gCpallldVwqt6YBlX8KOPrauEiwLNv6cBYVFCNnHmkNXnv7ZZWtkdtmS7oWypo
ube3BPz6rVz9CBvMtpNJu8fimngPz4HtYt95frA+wrwzoVO1L+qWMLgqsBTXo9Wo2W2x9z5r+5aG
PSP6RwwE6IBrBccXdFZtfg1gvjw1RKxfOuZe5cPULiNwdLaYktRggIGrGK4H16kG9gAfv78jrlxX
H3i7F3YWdudrt5NctTFKY8++uWoKBchn1eyEu0Vfa2H3w09S+/wMhhj4lOD3ePiCmDHuPdifNhzy
k95pd8UnxBN/hygTVFygXUYUBcJg5Vij+tr+iwojIZLIoH4cQW1cd0vYWWchCZT53Lbf0pfS3o73
YNwV1LU67J9TjhdGqZwb4SAI31k3rooYAPDYpSsI9XR7FNkWKYP6V2CJGG/tYG+r32lxAKL6DkIO
2tmDOgbUCBB0qZ3V15yL8tSbsEPPogYkN2l7Mrls6sJ4TvQlNqP7nEFxzQXk+895Hx+34eEjX0RF
pak5xO19zRU72Z1Z0ajzPq/aYVLgChk1G8f6pyRcKRvbBxgWVqfRvRHzIOadKJzINM37QOG/1Ra3
GAdsSVSSa32Gt5KPmsedqNVuKlscT6ggwm4RgaIHpZLMajOUNiWyhsW21MFfQICH5OCnMtM/5/JE
Rl+58Yx3BnBkzq2bAzF3qcDSeXHaM8yZjXWBHHwsF/ab84cctMj34Rk4uwBstBO55hqlVcTMT5qO
nkZDwSCwvFEanJJgxMntvB1ONxwzI+663bRvpa+JKRra0S5UxLcc1CKCbMViuF285OUAyrgRb+HM
ofeZ+e8h5Xm+vgd7LKG4ap6BaXIEgt752wFOEmDQ9GQntEhk73kdzezZTIw3rzG/+OCDPFpV7etv
6OxBGwEK3ZUYl1lQD4DpSrFEKEVLjbGGg8cwp1odJ0mqr1FQwBzoL+WEE5NJNF6T3Ao3nALBm0xn
k5fAhXf/U93h7HQoKtr9Dff3Px4fPJhTzfqth/3owH2NF8EVuo7O8Ma8sMr4EtEnAV6TawcdXWre
VWsKLA63G6dYrxcLmd/1KkVolr7qtVfVPdJ9PcIZreTA/Hcf8Ji/Jsb2Rngc/6uMVPPiE6Jp7ajE
UqdRMogs0Er3r66v0rD3OpUHrql88ljNclqHcJOXl7k6kiACCLm3k9fEWjdnBgpGHA/MZfvGBXGD
5ZaxUMz4srPFVIJh9h2gBEuR3A9sOw91w0y42KLsm9gzwuQIGL5M6f2XQiX8C+ie3EKlg7IWwgKU
qDOeGD1ed2sTar57eojgF28BDOWxmHex+K3OHEAV+G7Om9MQZbsYmAeFq0DraHjel9Feh6NBg8Fs
1G3LpHzpQp0AfLIzJGiLmMg8mIVhx+iIpMFGG1AT1Pyxhvsc7PH1q7phouzAbx6b0/BZwPq7hEAI
l5m2tUVHZ1qxIC+qGJuBPkN9uIBKsZ6X66KyyY0Po7p8cnWpY9fCTY5zK0UEWG7y2SyUb2gIqfAW
qnokfmHpEAmEdDzLM679fnGZKWOxnfO0qz1Ge47iMm9qZsAS/j8uDFsBmYXzLzvl7nAhnfmPrf6Z
xapZSaN7AyrPOedTQ06wu2Koi4xnLm3ip6lr+gFH/sdHdjgW1VUa4muh1JSzM1H1KQa7gBihZu/k
1hEhtqASzkOJvfNM8ZkYDJneq4w3aQsocWX0q2rakKuHNq+X/1KBIVOJrw2hYHrjH06NRuWfnPR/
FwrvZlPrMPgXjJC08qbTJvN+ykvgNGUyT0J8SnpEBysAep46/4TX/4OeaAXXEG+CfYqcDHFMjZQN
2Zna4h6rVviTtQyfNBssbfRMOdHA4uOmQKFCNQHhFeJPdAgBe3CXuKcu1xmKluu7IIR0PON4r0kx
ZxaF19R2t17bIqnnsgzjT8AZX6RhtEJIg51y2VmsbhNmVosHlC9+BbNonaOCgrmWLiybjru7R64k
q6emY1DSDi/UOUGFzPr706mK7m1IGebD8V9S/OxXYIHoh0kLe24qW8VIY49yDDNFl6vn1inB6OiO
Fc5xMyjXMfhHU6OSLDOu3QORNAXE0pERhCnOKso8RUy+DqkUoCDCFMd1G9pPgJgHs+3Hg+ajxUVu
Q42peiM8xAatupBZaeIr+HLWIZdZUWRT0nOCRjePSbe60bXRv06gIm8vo4JUAz/wS+5+D/OFznOb
cSN6KHL9IeSbaU40+zKjRvL4eRHn6xcZeZAzMHLTKyQLOwkPk8MWmPJU0Hb+Zv1sdC6htzmVhrjA
VnAnwB58oL2E1TvHcIZdR4x+XDdpGHg+Jsnkw27H/StJrxF1OlEpSXm9QNIwLJqwCtfC4gFJf2uV
2aNj3aRzZyEkb9Bhk528K3xj0CpyOoUM2xT4NMq46L+xSBH2b6Y8fwxLpQJHnWKJL2SkRIrAxkuh
Xpd/kCAlqOfedVPDnaNYZhxsqrAoqR181Pgkn0qhZf5mCWhd1NxPegf/XoYfMO366r4vu2dlZvqd
CEpl92ZXwlwh6X6bFFvpFUrTvMe0lZB9EQTVRD6QCIsJIPGMHQmzESFxcpZXGeYv1nWNDkJGePiR
4IxCHJXhdv7dAlGIwYg29azLaf0YiwOYeM7XJnweLKHjJ563gyLb9b3I30av8EDrxJ5xucUp1EHT
XYdXqRkxSlOmP8k0t7CjAhFH4K3TDBTIBkIta5AzID0EDEgLjX1ytAeCc7C032tkEKIpDgqvsgiV
esbnCGdF1PBAZOlg6u2UEo+3JPUxU4LvpqrPy5PGvsr6W9st8U5DLqsnjkve2oGlxurSJ+TlxSbz
vjfwJ76Sn1ELlJU2D3NbTi6RRYnaDrwrnrwcvA7KTjwOVKrXkiHRamiUvJ0hpINoIjw+K1+g+XVL
sEgOp8WU76fTQ23ZUtId9CYIMtq91XGrNvnIcwcNkuUSAq43W4RUkpPT0c98WFrlp7l11rRMYJxX
PEf8xtcQq5dGDtjSHFNsWXlZBMp2BUA64eU+UfZ/jRaERQNG5/o3fFFyC/QGhAXImFBX/JlI5OYx
vEdyi7PHSBnuf/Yl/Jdp37essOfxvJ/hVMopd0bVLDFbJO7Lnkx7bBDCxxpdNNX09HmbKr6DpoMO
6gCnj9jcMhQbXcE704lzr4CBYctvh61hC54R9v54MJPtHI6pMzlaW7McprSkXImF3WFAqX+kUo2s
ZSZ6PMtuW2sqhepnJicAekgehZMMvB4hLUL7YY4PEPz6XRWn/1+v4lUic6tiWKZj3nD6CgIdt+c4
92CTPHZYfQqRBjdo0DSqE81UYbG2mBi+msDIIOvmbP5on2+m0TZp2lCqMR1W3TLmCvgeQrNFIxf0
ZHIENBpvARGKCujWrNxcfuDSgfRh/gGH7Pi9NH7D9NtKhasUQQzifNC65QIs7+f35J9gXQV958Rr
aYJWa1cV17fmQBTKLrtJy1l4rLEKwF5ZYF8rHWFYVl8DUMFDh0KS5Uu/jRkoBunK1D3XUXO3yPrl
OvdvOl0A/IAQ44TW8Br4Glc0eqDUE7uB0glO1LvtzyFJoPub1/pNxhfyeitpRp7o/v6pneIOCGUv
30KitF5/Aw/RCPT2O/zu5MCK73Eem21frsgZ1wxwsmVe/xOCSzDLDJdkOMgar1FSUFzyTItzuk6r
/RXfWvBVrVmhG3ARXILsKDNbBCKxP0VeaUcx2PvEnzjOGmxxULzAjCwjX11e0auPKcq64lCTExhQ
24mhQuyLeTXFDvB15QVoZcBlprdGNlIclVD+uqSoRkVoSA5/SfaQ6ynOYLr17yBcnRrJc4+OHxmH
ANoy/ZyHCPJfK8uwTb137GpvZ8z/ZcdGg6M873Q9e5DraWoVKYVdKozhApeziyErqeUYkF5BgR8D
ZAP9rl00xqKRl8ExNez2ekOegBfBWOqy9lLMqlB4NUeVzs7yUSQRAkGSlNn7SpJxcFTw/rvNI/UG
9unclnulNMkVsFW/e4LojJ6JfKlWe7hsa0DbGq/o+eyHobrCRbgZ9vETJeLpCMMd4kAXweNXUV7T
EbaQytFSSKIavlssrntYDbVyM8UPoomK9jbymWltxsEnmq/+eEH8BghG0XlgRpBoF+xu/DcDYY7t
mkbOeABEEa545BJy3e6JQxhX84VTZp74GSd4AkSlzg4V8hA1IzCHCKRo4lsB7jx0xY6FNXwuQ0XP
DVhTv7fUKyTEcpwvPeQV2B3aj7/yk+EgEEI1D7MnwyFP191Qei9bBDmDxn4L1MB8tpmE66w8slT4
8wexJjF7UMgmw9B4Ocj2lPVc987FUYfH+B8u98+/c8lbZhqQ2PpXeR4t+1b8lhsmfBqZRXzcXZZW
ofakTteP8qOZ1N6tW+OhjCzlbsR9BIilD1e7saSQkzYAMegbuZ1jLjWpM7NBFSpQ1DPJEJcpIKRO
oFnWJxn3sGqvOtGYflyiAvZEBJOkOQW3n4urIEY8yVTLYLKserlgD623fjg0Dka5xeM2GSX30bsX
tdC5ur4FKQZbreOcHyPnAQu8ZgXO9b6/ACH6GkUOJlQ3fB4NAfm5cmjSG7fZl+jplIql75ApLdWb
cjRH79/3Zsw1Wta1gNZ5MRAQhImViILUKO7yNse4jt2BBXZtgZ3ksuUz3LXgyjSDs1au4y6Cg7sZ
wHNK4FgFSLNZ3RyKxChhymtf3qh8BBXl83JLkLY+uCX9E+Vf3sG20JgugJJqt+ysN2PIQB9N8+hX
yi+Lj+maBZBQce0PvMpgB2x3md9C9bfGMfYk1rgcLuADwRXES/6RpACAcrhYeIJ4k+6LZmoTP47F
bEo4CXnd6mtvIOX71cXjV1OV8v+vpXoNBM3mqar0eaM7Nb3ccELk09r/YwRXfSQB8qvwrfZkj6fa
mgmDYiGjyZTtk1BNl0huhjO7MrDDlihQ+sKMchTWHyiGGhTSORfACpDf4fKeED9/ZsVYXzb2dpDh
rmDdVpY9F8VI922CeQgu2uQLHRRJ7pldsIP2C3D4HQnNh/wvxGplqJhaNq6bgB03uKK99nBcNEs4
PltVWvJHvAgoObcvYn6Try01nvAtES+wbSkikl+bvwfwRUsvfOKSmtD18E/BAQeeEycBqU8KQSch
msSgo7jYLhsOJoEdMp1J3lCxvSCJn9ZmVEYsIH4doSIJZsat3skpSS2J1YU7hcqQsPUaBjqQjH4M
dMoZ4rLafD95Mumhw+ksyhi09O25m1jFtF1DCKxiZrRloXYasSL+j7ruY7jWZjRffTkGQItrn8y5
GndH1h/fRAjAkGJlMUzGREbjDV/QzpQQI32D1XubiFU+OzU3MFyLYW63Ajn4fISkhG2+9wQ0hr2h
sDrc2ZyqZxkLVUTEbFAj33TaV+PadBv9Lbo9aU6z1wdM37FQnuH7wsoT4VfJNZjz+76T1oziqYLl
h7uiSZ6meZ0AyKfpJiUZm5P1HdM8riZFsH4Flb+lWoQXVf7jp/VxXp6GD3KIA3wM2SaPmte5sjsZ
QSzEGq1Axe9i+6uzJXYSx1dRVdwN51LpYqZT4LA4/mhkenTGQ7maFQ/G72um4MTi+CEqLW+fJ0Db
0fTWenhZQwF56+KcrYU8n5+N364lIas2mgkrjO4U8mVqftgyaQGjVs7DdDo6FOyFABk1ASnnVuVb
qDVi2AwuK8vGXddkG+oK20OtBIWGqDSmir0hNUVT+UclF5T2oRuB5P2l643onkEijHTuG33sxLeL
9YBSwecsgCNEpj8lzzEYFQa53ZSyPquS2IHrhTABossAvxt+HCgoBDBgt4DXgOoc9lyfiErepnZb
2gFtenAoXiZIjj989cJXxjnQuG6jTY9bREK4BrAizLpsVR+8auBPOtYmo+ImtahrT4ssq7JoQKBs
97kiHGackK+92Y0dAGJuACB9Qyl/v/9URhX5C9BGtibsG8baZwPm0+GeRSUcvtEc1/z5uKMRs3St
lkkNz4p3vUY33aYCZaN7jHWMPZkWKNzEZd5QmBl4zlIb4DhDP/0atPbqwS27ZYgnDLwim9kez2B8
7QttXWpODc1KeJfEGSZqXPF6kBQ6yh2GHPa+p0eAscU+d4vtXhjYZQKsjraUrvZbOU+rXaHxk1xJ
qwBgLBurgT4LwAxTJ5VB4tWUlHa7jVc3crnrV7ejdUs+LJ14xb623/K4EHvI34UkXz5SAzFSilNJ
ISrfJcGQF7dSm1eLvw2+iUp6dR1qy6EnelUgxLrUmEztYtoqYYn7CxWXiTcF1vSWXFnvtPrmBVRs
ANxxbOizyjKK7wjfDx1Cd127xNIa3GtucpX3aiJG/P2u+Zq81tITTij+EI5FwBUhQYHk7dhgwCKL
YJC5dYqNI/X6HRbKPwIsFlr157ZJsg+QdVl8FA4MgMQADRQMcmVs01B36/f9kvvMfX0V++/H96Ks
TJTMxgrLqz1ourxf77qYZgdecrd/WhdPZkJpQouXjK1zBjmlmVxY8qaQI5kLaC5L5SfPe3LqbSeb
FTd8K8xSGuSAFywDAyHNmrTMMTYtWKvOBwOWFGBhrQWBS38tfC9IcIBk65J0tSQTwqpPzqdTGdJh
kyLmOFImm8DQ1EofNfcbJ27srUYZryQul/jKvyqTJQKBEO18AjsqwWH71lVgBzAfO0/IyjmyVd4r
AWeTOXvYBVkSV5hADgdrFX2CLvqM23MoWxKFEcP0MJQMDyiZZaX9ICRP/hCJflKPVa5NoyzABGu/
b7rdWRpD5wOy3wimxBLryfCpz+W/vb11ZFCORcpmEcwZcbdVpVsrnl7etwzIV7efYOuvtLvi3ezC
2cYplZP5NBtQTeAn4XXInttjRzneWlfxqygIydzu/xy6AmX7/xyGC8+XnxtE9rDchQ+Mmr8meYSc
NUAQRe8IgE6Z+9/dI4xBhKt+4nw20SG9eJ55Ta3F9UCam3k18ZcWaw/weO2gNntbcfR+VGmXWb2o
6sGPr0eF1Vq4/di7FQc+ssHaJwKYG7EuBpuB9vmPgtfp20XJ27KUbz2n1LZ32XUYPQo+SOxaa5bY
pgOFD1o4ti4JMEBfTAxpJB1TZmdgIJvVKgWIcBKsRlXFCD/KZqh5OL1W3XBpAZ6DDyVmbVTCz3z5
sFy1eZKGqYmuTNATLYkcbKTR8ZWTesEKSeLt3PwjUnpU5282Y7h4+8+01ELt0rQyog3JjCTCnZgz
ErHnTyY8t8CpBxA3FmzOlpLxq7Ew49SLgxqfNEzuHGxjvHzVwKh2EV34Y9O6BDfysrEnX8tOJBSE
T1KGH2caKmP017urG5++NsrH+os7c9m21VBsVhErpRlcG0tzNS3HWH8+iReEqS0NxHfL7K8KCsop
f1ZFuwFU7gHnar/VFUi4TRE8MaTPFdl60ER88cVJ7y1ZvT1zqZYah6dVvB9Rl0xQ2XtreXpicqk9
zw25yoqtxJyK1gtzXAxuVdGdLvymabsW81KR6oBSQZQt17XFUEYsuuzSP7YQp7G6rqcYdcnsN//0
82DWY3JB+wMZ4b8Tda05sRTcEtTN9EeDNcQ87OQceRp2bykUlEKpZLA6fwJqa806tOzF1Iw6UnKc
/JyA0J6oaXRbQuMW1vftvs88XuMXETIgEuUn9JRGtAxtuxlJ2iLX/Nq7C+KJssB2rLXwXIWwdW54
Ej1/Uzt15bfyNYFVj3h6CWQ+xtrenk9gooi1qj3I/FQfjPODqyDNBeCicchhmVBk3HrPLV5CVc5D
BUjvn8k94kbnri2Ta48DtphxqPFqoGhkBc3O1IDbklWDahc56bBx4felmz6F16B4xm/i08hiXV9r
5IDYkdz+J9pBjoHhAAScpyI/fmLQtglsI/bNRVS9sAjYhHMba2ECT7HPIX2zXjBWZQtmIa5MyLeZ
K8InKTrRSIUUTM6ijIPEjfWBEEqV4fwzKllJ4lDt7JZLutNHjij9BCqdTprvtRBaY4afF96KIKF1
UIpLC4wMx7JmGE2+c4E5+nsZ1VUBIC8kcoMy8dvlGt1m8DOb8FHloCkbG/kbaIFBBcGKcMWr55uU
+3cqSZ5uWM4s5V1RXmpbifwy54oYEIotb/pSZhioolL1P56sm4viV8DGoRIg6rVRM1qcfvOoEiPs
FPmF5iUQH6abqWtdixk46Ig8MY7p4nj8h+rEeadXppgIkE2vS7QPHc+ef+ETaqptVlgJxsVqlEoz
JAkdNYdDs7PC8JJPpk8P512AgaKGGJg9yrQ+FheT89c7XdGpqdkrPdvalFaXj1ZPeNagLDkNEy/X
x/wmZN5Rp9xirtsmzLeIMJp4moxQXSLMtEB3eD6we4eOKjEUFZvD4m6xy4eM7IWBmJesU5UN8I1w
1QlHJTBHpWSzt9xy/tU6vLAi7Vrxiq6VaXTxXuswS1EpYLCSh5/QWyK6PHqFUP1HKN92Zxng55hC
+x4+d9E9fzMEH6XKkqZqQZYYGAQBkwvg1isGKQbkuGd5pvVpyymYYW7ZFZYmYQ//2YDJBJ+IwT0K
54tyLnfk3qnncnEu1SSpBQBF3QBza73DbKMBjuWyCTUkQ6CsKKenqjiXtW48F7K8mgCqlqNZFqlH
5Pz1FTiRCFIEp1UcwnPWgSaEMjh87vd7TwcsNz4/g8waUDLPKVyv/JmjqGmA1y/rt4hEoAqzkWzp
FKMhjEt7IZwO7SpIxpDOuxaVXZQdFW0vq1UKicZIhYPTEq+MDiQZBq8XegdAzaQTSMHKysg3yZEs
+iVHvz7z5Rp1wGskJmzDIrdgiJSysnf9HZNs7fRz2oVRT84Sxi/wUpNqOIJqY13/87LxxmBqtsr4
bHjm8DoUB5dBB1mFTP3qLj/5sSyEYuE0TzYMPDcnARklws4HDrFB3QLbt6iysFeMoz+h2PjK/dVK
xG7V+FJIExiTBZi6q26oGMT65vrjC2Pd08F0S38ZBP0vbMuD1A0XzTqUJ5R4GW15ElATAro6kzjE
3wA4ZX8BL82CLyE9M7Y4SlTe3/nuFexrWSpCWt58mM6pkVREgRJBETjpVg5xoyPofT3/7K1L7FyU
hbhdLk+QOy63L3XrezQK10v6EiYAIkFbGxAZg4Y+kQxnZMYzvB0kBbeKFsK9TMj90dIE98w5JY0y
W1EfYyq2vtbQePvIME9e4xUKxPLKXETQzzcr1/lg+0Gp8uu2G+uaKWWFrBqt44HPbw5QP/De4Pse
dz+chhTAuH63Pl1p7GNosbXllBjXFnsxjOogI5vxf+9MEVMwmOlDeLYyjpD7l0MiS0ySuRjcHBEV
nLsm3A/PK8+D4QLll1ykOHUgOqMNqOuGElBfGhJWYKq4NlCQyzT+JaRVFdlrOUBEihokOIa+xGci
/LMi6yRjGvRzxR8ddU6GId9EfzMW7X8rpfHPcoUgjkJZ4WPAFHbbBfQhjUC/fqCdQcItSVh1ufBs
ZDn9ycwlvI9ZiPl9Zx4mPZFPCc4rCVYpNDZa8Fbl4sXcvRZvzGEhEdkGrvIPdR6hC792EK/q/4DN
mRi/UcLcBoVp5eaOj0I2mORrENx5/jxAit5wmaEDA4X28swWJa9giB9BG3ji1nHswgi6T5hZSLeY
CUJymswI5xKUoUUsf4wTS43KVt9/xx+HsvYIpIi1TRb0wyj8MeoqrMRjxkJ1XXFzq+KMF9R7KNmI
nFfz1z/bhAvQdzybZNOk0PApF4dWl284wOL4gk/CPMsnCx/mcfMkYOep+DuOIRBqaYpxC3u8y2fY
wy9WsJd6UFNVcwTQzote1/nNH3SwEBGt94FFn4XlPhynaxM86fJb0XEuRH05XzqnrtCFB9fxTplp
XBKeWkLiM8NmicNveWGLIvyc2WOob/GexVjwCDlzX7hvvzhLBLjgImQdnBsMWSDA9Zqtx13x15Nv
r1ydI/tvwub3VadbUYGK3C872xDb2J6jypA3qtT1G02olW4awFETnXpaJPIvXUo5rlbRTnbxUnUW
wr4hyhBcLFg7ipyfhUNQUHiMX2VG3TrlXjoNbnfNYnBhhrLFRsGKZMQKLgGNPbfj7YKgaMSoIVay
dVOUvYFEHcGope97BzBmXD0GkoQ4uENT4O6dWM5EnbKTcnrNrmO5NQvUF6S5mHa54sQuTuksDkvp
0f4261zmE0rHiDK3QHq0gTFQi9d6fNM0VJmnZ0CtzTLOCql4fgBcpI8xKSZhOxuObBUh1+dkjbpn
Yi2qc074falvoZH1OkwSYPvL9Q+zAkw0PYfBE/ErpWX2u8yMHXYXszYe5eS3nDD7bPSlOT+zkEUB
QAdT4AeJdY+TSHMJYQitpPMRVyNuzaiJ6WjXpy12avftkGI5M7mXlu2aIfcHeP1wN52I4a8c+sMF
O/FbB8fCzgicH2tZJ/O/yT5IjLQdobw42jKH1+H0MAQgynC8WqXxLUZpa/5eXkmpoWUCJ9Q1G5rg
rO/92vRRnsY/kpMI4/YxUbhcm4rGjj3JDor1n42RzmPKRX/DJStc7Lys6jxc14vaTvXEQQUeUPBb
bFwILhWWpkpMpJ59TNpmh+3SnWEoN4r9YyacBw0VoTk+fdlZwF61p8uBKzSHaPnsDjWB/8NYAGku
JFxLjpIFJRAbXq/+HRNye+DumR3ctFHXHcdSpVS8wv2Pre88imiV1h2ViPEa1mae5CfnTlsMP9ZC
+CE4wJc19ozbSe3t+n1gdYR8wXFoHZT5K7UctDqK8jMfhRzO7T2EXLh1n+QMRy+76F2+G/D+gbkA
PcD3Y10kNVZLZDl7KDTp52NgK6rYFXyS74OBHjT1gMpg8YvE3ObfF5FQqxQtE12kdsfQnl3enpCt
d9R79a10S6vGrygbyHDXiZDtVATbRJ3BL/4WKfMFBmrnprKCAymm2dy6K9QLWjLOujueF93ssnva
aN9uBtoxmmUEEkovfJMepAkUhbTqeMz/fFzvKIUznWV3royPRWZ3oeptS+kGm38klGi43wt3sEdx
Ul1Ku/qqhqsK7b0SgAAYfpZ6OfBj9wko/D0XFqheI/lp40fy2AXV0vjvzPSC57FgiX5Vo7hj397T
2PKTctBeHgbt4wuf35h2WobkZfI+MxefI4oONLBcsmGQZ3Edyr2oqyoTRsbFFZirPaiNLyILnOmi
1zVLqKsJ4chEruHiCbm5c+GiRRkFyPoKlBamczjppjkudR1ufuLaN/lPs/+NUKs/rz6lnfQpCYn6
7SSK5dsR+Koi6cV6MmS/fUOY47tYvRFWgFyApqEu1uusDqhkXroHmXY91yuY5WE7of8PBBoVoSP2
sYYzYrjHHCSkVxiNOvzG3fbvGFNrf29iddT58bYxpQiOVFY+prHM9X3iefAGsWQa8j5HQOCREsZu
6Jnmo7/6q57KwgO/J5lT9Kr7ALkwzMaQtPDRmamgWQShhGQyoB7Q8sqlEi6e3TQZq5itAm3cMmwB
o/6c8B2QXN8qT93Ib5013twFKHeNPZ7SLjFbxcIHUf7RlqybINlsk1gymhOOpRhy8oa/RQBAe9Z2
UNmmqaLQYMqtjB4z2qdurSmXA/8YFI5xX1mmymaOZUciGSZUPXDq0N8AmC5u4nQbZzpSpaVBBywS
/VGJvoppjGqJagNBmcskSdjkgH+0BZfrbkFdBmnQ/V5KHGOUGYFP7HHDF0WHRb3nvRS66UrJBgiY
nZu2kgr/l/JDQ9egbiwF2YMNaZ8Yxr/c5hy8gu10++sYmCIFApb43y22r7YsGuIMf4O3NUECVHZq
3JHw/YoXuWUTYl+FRQpvmqzlAgbYr4Lwj5K07ARyUDQpE3gHaUROriMXXVZZ6viN2FeTZ2FkYOf+
EGNJ8Sb5k8vXOTtCxU33y6frKSUwlSTEuDHkvOW9OAHOIKFUlcK/rbkVweBKirR8fuPnDDqmVb4O
vKMqyOBjLDKXeDbIfhkAC7pHo9U1NwXpfgBU+Nti6Bb6R3M3x/xaW5C93ZpOJdLoMdNLjj+WfZQe
bXYOqW71MJztTItEtlPpsxID7P2B8kocpfTgmwY2m999cKSmPlfkggtd3W9D+rPP6sDd0uub/RCm
Q/1ijFSfEXqk0Z/djW8i9XHVzLQNMUsaahK6kSWSzg+G9Kv7zSuVo5iueTzEF7XaDCDouiJMGR7l
7K+3/2OaphhfmK/4QOUuD/lpD+d6eWYSf9kfZRx90nzdq3i+1tIVNWp4zh6zw8IF2MWBpfxRKg00
tffyIIY/oOjpxnVZhObgpBfbpCFc4IfZY6zpqp+9hXnazyO3BJvcPG/EOommhzeFPlWk9DSAlytG
AIqidjujHPBTz9B4Xprx3/IgRKAk8PjcgAuD3Zv2pifO0rT25P2tPs+YRW24tjC6ycVsbmgihIAd
PndL3SeLTWsElxFF45tpwgwFnzQyRTVfaJ7sM9CsIQ2pIdQ6qD8Hij7crNW+GywFgLs3oaBTPnxi
WvsKbCEv5yB4GFKmtqey7LhcLd6kphNjYogrDVnR9zIw4l9X59CoKFGFfaLO7qdXet0FFTQbOD+u
fjshzxdDa1C5P1ksdYbuPwsRgzdAK01GA0MUfjGLQkWDOV66jPLl+/gduQQSjq0opBDJLXOWxxxh
FboeEO1OKU38SWVJm+NMmDELpJP/sDffRkS8PsH7c4bbZoDcf3EZsM/39OZG/jIPPWvw1HgfSZJL
RwpgwMua2Cp0MnaALfurf15c7NiRppnzAqX4d92Rp6W73zzlr5H9ivBPXt1lBkL2ELINU1N8bgHf
whtLrWEZtdDtYQ7mpNh0dW4iekP+vth/aPqJQ0dP7TfS4rpCYEihSebw6/uv2o9C+ZoazfayzEK1
ISt0yozY4DTPtvi/ctW2vIXiq8LIDl4LEysEtCG795v4hA7mFugG9xDtQtPtxxhlcnM6+j/Fk5Fo
BPUuSa3PAj6tHQvOH/tbXGn4FadnBm1656sADnZnHZvZgG+JZhCzlpR5ueJW6roN0ue5qYaA3LrG
3x0bo2ttLYxp8KaQbWPenhUpnFws9zWc0wJhdbtBhrvLSF0phA9aLgjfuyYeSHuG3gvtaW/pQJHP
KH384BOo9+n3ctpm8nBxxL+7g1UH411GPF1CMBYFBgFLReGVMjktgGPqFNSaY8OSt4Ffi66J2rLH
kof4C1uAn2jAaSBwzIy/Wqf5ajLYwGbYOXzFeK7mYWNHoxzkZTTCsEWt27N6Q2/39IMBoTQzJyek
BVv2RNOobdrnxK7xYv9JvhkAyRr/SwEcREPE/NtX9wN5B5ntFNjztngaOZSskJphaNihvNv3wwLH
d492e2Zy4i6x/3L3/iR0wm89j0rop9N9MDVtDugKBEkxqU9p2FXZLqfWy3OhKcqIrSxCsfLSzvO+
7VSuL7psiLWgFi2r7cXH5G3B8qOAnaeeO6ZgvQ97WRyZ4U8rsrd5s9nrWNOweKOhyaOYijMdm8kD
ejVKWfvkSYX9KOdurt4fVLy30sJbS9XnvdUoC+mSIh6oaCcQBTZP2x4zxsFdXMEbNe2X0/mAhJqD
pLrTaEVnQaDDnYBoI7EXaSkPN5f7MMKOwM4ataT7JmUX0s6yOqdmgGgo22MT2yjjgvPrLAgnosJb
61Xau39H2xOsyBiKfEWkfcQwbKLYLY6ddMkC3MokiMq7wYn0m9GQsV5I/Fg97bF9rB5JOptgzqvT
imOIrMV3xVt1fhShlhi+qlIGwGGFZ6dYXEkteBST86Bkx2w22cuNBg9Ibdma9Qr8i08yUPt2BJJT
Hax8P+ZUYAVO6mtDFfvJv10ybvMFnFGPVSRs8X2d/qgMEiZbM4wWA4ONSVSNo8uAzG82Skh4DRHA
1Tsa1BILp9vvscEbBSSFrxVlW8I6AduGSUb+3CyK968OmGRuN1nuTY+vvCNApx0DrtnSus4byAF7
oqOXm7L54pzW1vCvHb1hyn2VK0FSIWEOP2T4ArporsSXEGXqQibLaMPC6WjI/LSl8Op6GBuHFNdj
zjYdCnh7VgvEifi6k717I0nXHnqwF0x3dOqIQC1/6ape31dhhz55ye9/BmXdaFIGizO6O+agFw5E
c7XSsZbctvavhacNpRyw3B7PGwHBbIBxazomlXBsLUB+09uJwQf/8Mheo08qWLM2+RdxcJcbSBTJ
7H68Xg/6Priay0Xt+5r7Ck+9oCuWPqVnjVEBhRYFA2RWbBvURPAB5Q5LZq7H2YViQos1tEtww4YO
8hWmTRitF958Vws/UoYrsvVfIpn0jnMglE7WECTIe9BtoIdaSKebMChgDgRQ3duF8c/pmgPC4WwZ
X7NOoydPVEPXZzjHCnmA46BVdK5H4vFJTpJxEcvb2XKRfuJoHtuTkFr2TXSf2aIpGItzWO3ACvph
MMKvGA/Z8+KNUjGgXvGknS8edhWpaYXWgfjQfPrB0CEVrUUJzhD3uxCk0IpvQYnS+tb1kauAoYFy
BmkkEp46nP1Vemu15XpCNNKTmqZQxdabfLh1Q1q/uJ6cEy87huhzKsASFXN6LUqI8fAZ6b+E497y
6MlrPS86OIScxjVVaRIo+thZ9DtnMD4VISN/fr78nSDwZtz5UFWr7LQikseNzAPpiZ5BpVlkOrSD
Jf6vd8j05u66bcbkvepxDVLL7egSF6XJZ4kNzF9y6FNLnqY8HF1CYEFokph8n6R5JoRyAEabvGSs
sTD6fiSo70lyeIY96qqa5rMzNSlgN5+4tL+y6UVnUUgFTT1+/EMlRif1ZN/Z481BEI68p196drcK
kjygIyPaE/7zk13sV25UpBY66T5yXMZWW5M3vnud1HOcVXi7KHpzjUr+ecMgARChcmHIOOTkOTxi
39GocJVs5jqtK0odO6wlmHslNMrGNLw8R8IOPyQmUrjnWQ/kKYg0caI/jOK2qFDFzltcQyqLrNnl
DZ9NLpAjWWyneVE9dtKGdtEHZW2MBrHfrq2xwNtD6FyrhPTsq1zHA8AzFTQjtxMFiX8dPg9Z3ePA
GJQelwt5H2N1UXUpm7wEOHZnBOb8uVFPN2WH6NBoxoDQbFOqkQOUKMiTTD8bUjCMwdNiZU19I4Hr
Ntp/XyErU9nh2tyrE+0pHBF9qANEPunro+P78BPkZNrbnu2LI2NfNw2UWz19o+yHF+avOGb92qN6
uZoMDvT2fDpEQcYRs8or3MFQyEXRPP3C5iJYLqaIZfHtiqAVV/QK+/c3wx7DV6af41n2Wm5QzKwd
0dudw579AoxHs8cum2Kn5s36M0I28IDMcXS1qornXVqI8//fY7JodAPv1+D6JTBvNgg6PecvRBU5
wt84+xtZPrevIZsWGvZ/E/KX7Ae5p4cAniRSW1X08OeNaBTKJ4UgMjTMd1Bvu7ebJrqnCRqdIQsP
Bh+4/+1L81azCD6o/I+wunaR2L1e/BRcH16OE/ZklCuh7P7kqarKQfM8zKK728RGSotNpRqp49/0
l16O6UXoXYwbkvxDfPmXHNfUVVNTvie3NNLeXOCc9qShsTDVOoHPWF4vBb9TXdzpvw43aDtUlA6B
jP26WpLbSfnfHy7NV3/bm4iVamrd/Gs41Lyu1sQrabVUZSxfaUIfkz5ihtYGvi7Ulc44HhUKEVPI
Ju6ZCtHo8xWiMPY7U5hz1S4iFxFQWevhCUn3Haiq/EiJJKPS5kHd9p4eBximEpMSlQQGOMGGBXAc
u0GGZngtqEk4m4z89Ker5b7N8ZGmVYaoeZgnT0L9Yy1j69t5rPrDkNNaR8P3znu0hNEFiYO56Q1V
/m6wfyiyIxHjmREcvs2vY0dhRloGUTClHF3jTnCU1ajIbCFYalC1n65uRuU6N53dJgQvmpAkKWij
7FPArS/j8nlDDRcL093OMt4EWm2LMplFWve5kR0GWFR9v6iqbF+2lTV1s9TOU/wRJJFlL1O+iehw
90cV+ovODt6o8iq0WSod3lrqD6ehn8/xHx0OYGdHBct8UzJ2wGFy+8Le+dnFWG2YwmEjmbhFFf3O
Iik1irKuiAdoIQYq+TSEkgQvkcLP97i74p6MqiW+gvZuTt33gfDETrCcMpZpP09P8SNN2XUi32G+
45Uyc5+ZYwqolEa6qlVdjBf2zrqwyJ/Y1VoAtwtszLGH+aiGAsP5q32/mJBNp5hTDTliJta0+Qiy
clqrsvWxPhccrAKueXloXC/zO4VN+7teTdyayXSLkM7aYHXT9vhvXaNRhOiC86MckGhbAm54stXf
iAgO+MyViD6KzAVpW0cldNFZdi3CVcEtfEQcY5upZpDzNw/yYQZgUbLEMPRZwqzquMUxf8hrWhrT
RF0aDiUEubOKiRkmsw57/b1TN1e2mLOJ7fyOJFDnEdc6ky4bEZVM5c3Adi8diVWlkiy8Lp5kQo37
T4lO/8DQ55RaNapF05nJp6BhctI/bbHvGt9mwd3UEkuuTSGbb5aawa8jCn6heV23Oj28Mm6QuWo1
Zc+gO5XwqMdeGqA/DpbaVib2T8gNCwbOy6dyFt/JAxWOo+HEo+kaQTgiCXqimYD++AJONGNEw0Qg
UzqvO+qDj1v8hQbC73A9IICwhPB1lLjrFNAR9RQ/0L22LYaGhh28oS5TC5n+G57EoF63d+hoXkYU
KBaIw0bpCsqnCS2KbVhvf9/7ArXdrLqACoLnxd6Ug4HvZVNccwSJBsw9NHuvgTpPUOfwx/SYw1xw
oA80DYnhC0jPZcK6XvfWHdVoKeOR6b69z1Rdh/OWJMkLVylQjBrE2/xnCKq+88j9H4OuhOv1JLTT
vL/s+Nx5ttxLbB8RQgIwKLVSeuFcP/MJ76r0pmvC3P+EVqj7YEbnTsUmW4s3jITqegEDOoWaxPvr
kZQ2B+WKlzlELA1H2rltiXur6+92MQIURvBPg7VqTZXGIXAXnOMTOh1Vzvsz7uRHx1uFEyQpkk9Q
BE2W/he6FlGp4KBMvkTNtdfEOX8m+MIXMNzCt0OevCZiD4632xu1/64+cAfrWturg0QXHFD1rOhj
FpPYobOovPrdJeLWROm+5SjJt8yJkbaX3qzX9s4RpXnXGHQKzG4c9Q+JVAn/ZdKzTUblcKm4eDi8
GyhWw/IqzbXKh5p7JiiiSf87qFFq5nHd6VF3r1j1yHz1RGSA7zMwSJ92Rfy65r/ubdd5NIPyHO9x
DCTPQcwA9Cwf7A0uKg27/YzYIoJOzB1tzBYImoAxc5EMyDvanilq2w7/tDh4am4rNaXjDp04HBQf
CSOPCtPI6B1/vfLw7hkwQOrBR2sVmX+4eC38KYJBpX2TpsokPIvAyCahyJIyZ0UowBe4wRg3jF0M
++TA/EGl54Y3ZQyXlDqTxJNiD/BzuDJD39sPiFHWKXCG13Es+vuJekaAmTyRHXKr022W5FaumnxA
XPwPY6BnXFwpPKBogkkPehbZRyLXEtQQbaRDWKcv5Npd5oMnPrqxxu1rYbWcrtI0jGo9z1Xd3uIq
XlnpqS/+OugVfmkU3BaLDx0ftlJLf/Ckuu58LV/T4zxhLECXAwRp0EjAVtOcfbXBFAYq+Vt56utK
A1f31H3C104zTkhJ5jnLEaCjDmYFnhU55Z7c4BTcNaYg6KNJUvGetNV3hTN5frBAnv9jinV2t5P7
qshSZw3XMTEsTT/Jwxst5aQkYCpuGNhd6iBPbCUOrxgIP61N+TfFCuPsMymiePgyRRqrJFy1DH9C
dRTQeE6ktsXy45S6wm/EKBMXo9LiFrFijm06sYURy9btUJOZnkpOuaDRtyxLAqo2aT5/44vJYvjU
ww+2o9UkuaQx4fHLYxpbh6l5USF1fgNNqnT6SNIvVLCet6Op01Mt1dBsAx+KEfu3hnkN1Sv4AIzK
UWbAegx3aMWU36xtM6tj2Qhmwi81HtI8olaz8/DRMwh0t+tewkqnyLx9McUvRiEimyQ9QVdS2ftu
Jt1vyOW10Kfet+vMA7N94ZCW6B93DJgE/xlj6BYd6SeUdCD/V3d1qqKKDGi+Wfuntejxm1F/0NfK
72lqNj7ymFUXV9lRT/1k+W24wbwK66UqxmaF8yO2PxxbhjXscbXvJiTU4wAufOGxCu1NqTvrRq/Y
WCesbABDhRhOHLIc5CFvJugokhIwc5nGRuZ4T2PJIMxNbZs785H0qvBRUTSoB1RLqNSPoMkq4vhD
A9XOJDbs+u/D6b/1lO7LZv1DNoa8dz8SUCHHTNPY/IhMsszgjI8xbyXVvEJCriWlUEm1VluB2kRl
kvymQY1kfescwYPf6JP0ldn8ObevRA3Hs9y/YMjaeD5l/ebsx+hQvb9nLnNwOEKSKk820pJVdqdn
/egxSFAzWDLY4tUA0O++5YMTtiT7j1KH/kUd+GroywlelSpMv7SV80mDuxPhyn7VbyNL3j1yJrir
mP32K4QLo0ObeaIW8Uhlr69RqmDV7N4U/m0YSmw7IN9RBODResmcqgEJuNOwmFYwWuLsugf8Owml
NgMyA6lgwnqkTmnh6LUY6L7D6irMdBzc3WLEmEGXXN0eHTcbTaGalKLNvKVXtgryM8WssQZTj1aJ
1lZVME2jR5f/5SLI+GFdR0jc86FtDwFjPiVqyXhZhJmuSv0j4gv+5IkdyAqBus8HJJJc/gbIuyZF
aVHkCBKGO347sXrtYPGDdj+2/2hbCTCQWNtCtjej5xCt2D94+sWbpzZLrZFcxIxljsoz092yE0L7
wHplf9tLVm+0wldZwXapJBbe5ZdlNeBem8XmLs78ox72C9GtJ69dWPg8HpsT78dtwg+OsVcM3KRH
iGBezpNBBWvzegviB9agIpwmo44bNMNVwMpzaSrHw/8Y1xY2MevbiYnhn2cIWEPwZtxQ5jkqM7XE
gnCQyArE0t/UlMwAJkFPvkmZl4Pfh7uwuE5dMhfcoN5Qi1TczpEXMhWK4veGT1U5QTc8/6Aad2X3
noKue2WyLUOgI3G7TxYxxSsY6jgBAoDIUQPHJnIeM0nXbfkxEP9aa52nuUb2n8Df366t7PlaU/bv
RXcybwkBkgtAxNRtiux43MJs3V0gQYhw2Jr6Gogw6dPDpzt6KsZ557QOB7cWea1i9OwR8bdKbuJs
ThLeNuU+y5WsQ7iCmENZiAsRxwVnAV2fLCNqShHpITHNQdiogu52L2DC82ccbWhxol9VYex8NYRC
OBj3wOhrygj3shz5F+uzLBn5Jtfb64u3CxcRN6UH99s40dS6n2vlTIkKGA+0Rd9RIHJ9b2JA5qKT
ug78hPQDVJGFX8+K1usFEVOia7bRYy8qPm8/3IeIaZYb0VWodzJ1iwd/Ji+e073Umogro79wS8Cs
0rh50d/6MiZWek4cTv+SlonNXX+1cDx2xXgXQphVZOSV/7e/R2OhWFZrTnPjpFbKi6g+WyFVN2AS
RztKkQMLg/rgY5KoJI93CMtRKHELTUkRY/GJeuwQKhPi7h5SeN4d2kzQJSL75J2jDOzQo5GQ5Cc+
Rm7bUmdECpbyXs8v41FKdSII7F3ndazNYwQUX2yjq0+D/RcK6kUUr21vlGbcuXbSF7ycxoa91d6W
g5pqQvWj2tBqekYiq/Qskbx7pLDgV6f19EEO7YpLqw/66zRHhf7OsUNQdaCw6ZgA1eJGzE207r2b
oClJfKelqDDNWVci0iUh6GtwkCPCX7Y9U+8QhfAiY38/5mSfowj8CYkwOmsU6xT2HcGLH3bSSsv+
cTUALLBBhmmWpsa1nxalbS4scUJodQUtA2Px5j550ABClE70eWxJa2lT7yj+HFlH9S5IFTKnrzAv
Jl6ZI9qRe/dcyjAB2HQwiLFpq+EhBLl4+i+7qccYztiw6gVSsw3lJNRApPUOyM04QbSlZW5cJpjB
z+b/T/jSvzUMvQmc/98Bsnt/kVwbyWmfIpyYKHoHl9IzPdPO5AoBlpLgERs50ZwsqC11VS0PEH6s
dN0ggUxCZ7ArwgL0KJFGEWateMWJBEpzq5zYrLUpYBl3yxdbDKAfM+IRhHvLGllSOPHsAG1x7ZZ8
+p5KK2jM36+sNd9z+gCp/l1PlN7vpc+F2wbFVh/9j7vkdCfadAaDQviBKhC7259vl/00GBD8L5ms
mj1Ht6sxbNRm2fKH/lgDodyJmK2yAPJg4CEU2D3/aGizVVveJWnJEEL8wJa0xgGwhG3niW45iqX6
lQTZrha/YVG84HYx9T8pDwtvYBQB7c61RIod3uCWGDqfx6D07nWRueM4dwMjyLhyyyi/68H9Q/aO
cEfVMMM3MKbQr8PSSVjhokkx+hQnS5PLYyuxO75d/qX1vECjoLGcJp+yuyBQcqvb32CQPdFEpQCO
ZngA29hHaOwwUmQXmKUPCyrYAzWbfWhvPYdjnR5p8k1WlCMJtOyyFPBJwiV82PJ1hPWmkeh3Ln6B
iwkKdjDWihJZsqVqTPdZWGYiFH4uKCSo182uqi/6AP2zQvnTV+ZcNDl6S5CeMILMPwElt6VwlOqq
CFByFqMeZCpBxY4K1vrWJXNRcAJs1RqJaH0B0CjfsuIX/xATWfDCj70oKH717YjPiYYLq26YwNJm
JQb6xmgwoj4zCb0KvkxS2Y0PWXG1WzDCPh+QFFg6DLl6SbxQkrw9w69AGSIsI2Fzdv5roXYkRKbl
0044XskjZRVcw8e8Zgj6bx3jCWNYDp2cPCBwp5jeFk8DUfJFhPGBzKb/ACq6u5qwiucYAF1cvGns
MU5mKd8anUZ9hwQJqUG73tyUqW3NP6B4SElLboFJ9FVJaiFzkn2/pWWoNPN9glrq+Deq1gUtI6QX
zkmQUS14e/6b8KlFhG91O+4jdvgEYU67IsRoRiMWdWAVdI5yVAjFl3fYKnTuKUoDvSXgfJf0mh1I
BjN9+QUAcubZsB7A/c4hTlcOOIDCzvyweTGHePFPlRcLbKe9XGCiCjvN8B2Q1rYjObj3kiH39vt0
x95CX3X4xRLLFX+T/Mc2NVmQw2Tco5EBS9zPDNuq7pDw0PlSTYLeQ7lxBSaoGVaxWwi+B6zS/AZK
gU/HyL7biEwWODNum7TS/YrBAfT9Q1UIDpIUjOkCMWRTX8X6q5Rcp8IDCS4CZNZ8PFF/RcRb2gPV
ZzztXCC1CgDzYnZ2kgzZuP6VVSyCoagT6Ao2RmmOWSUDFpGtbWolBqV2IEQI/N1o2dqz2xDqFEEd
37H2e8FKVNvGty10BMsbLVkmoE1U9+2QEqt3FV+lC6Sft3T9sMivNfA8PUNMDOWsFnNwjy+xFs/5
Ctuos7EPr9Ms9SJdqzESK/U1ss4n0jGJmDF9SurcSr74vu9dvzoPeyo8M3rtDbBYE2UgyJ2AQ6jJ
UHGsM0BAoSWtAROObM9LcNl5Cw15O/5xUbjr5/7JO97TYYR1QR184LNNzWSzsI0RvER0YLaOraEG
QZyV+FryZWtG96AIPX5zvH6IzxXd4Z6XF3gKvZT59U57KqKWF91sdvx9y36XMMDvro03lO32ay6K
h4DhCRon/L4h7qUKEfJSea+7IjSkAq3ho4SStFqshx+41ME4ZWbZN+XavDpNLtn0Z+6mJwgv5UPc
UbjAjNF8njXqHqJoFyW5rXerzU/ACTIaw33B1HdaiCozW6Rc6eL5pzEXm1idTrX5qg0S2p+NnJ3Q
GlxFxZgZ1RPL00PmZ4Hp8fbFR0CLafSMWrHSW0kceZFsqKfQrnv1FkvchalmOc4iWVh1QOtVq69N
BTSw90p4YzLLdzX6QfUVaGCTJ6msvb0nqYXz8pnTE+v2HTh1ECFN92B3MfzzWdrxqP3xLBxhKUim
vs3Z29kdegymAvWYORqrx/Bb7r6oXAUmH4oxlyx3GWMjvZVEs94ptRYdPYRNfnWgZfeV0e4eLSrV
9/Qd0wMAhsjcu2dGo2yDQpBcoVO3XcBkos3GcLmBp+CLcaH87e0P8R1ZxTkKVoioPkLct6/jS0Np
n5+Qe5Vlbt6xMg20En4tgVgShB4PypBncfh7gIGvT+8qVBs1nUJ6FUkYSsNgfSYgB6B3ImODlMEE
l4QCnjQpdfqozj2b7iuM5IuYa2D5YiRVQzRINKBt2k8VJrvA994IxdaQUgeBJPFRAnMO7JYcKo5y
vf6RSapB/YDFbvPXSbRdM//yX0RvSSWGQyfqD/0HkzOOt4i7OVyVFi/oJ0m4hT/nQnxxw6RfYnT4
QYDRFIKTbo29PvBe6bDfz/SrlwXGclzvPyuAkcC29QnkxYioLxiNj5zDGWg/XgNAjcXZGaHdced8
yD6lv0W+oQsXUhRFBbaceqC3TJbr3dJx8O/KsgLd/Ia3VBbPYfUlvkhIqfsWArZ0m/x3BzCsHM7r
HaY5V5QpMPvCT/w1L88YWSgVxEYnq6MVshs/SQTu6fHZn0mxWjzk9dzI+uILs6e6iTVA10k4bDPe
/O9OKTM0ZjsD+jtGRzxt8Sz512x13o31hMeRm8RxU1e3ZBnb9Dz6sZ69piaP5f16vgqtPJvec7Jd
DrRy5Hy0Xkz9h+/0mru1nwSBEdi62FsmbWEbu5GfAg98MNbmtEkMI4vcSGlCuNORAizPqKGhdD9H
CsskA75r1wAW4LAaQnHMu5fPFqXM5xIVfyxHlRyj9zlE/QHOUrxfDKsPVZSy555xv/1YJOS7246l
Qj7EEK9eUQA+jERMV4w5ROrNbe9yUi4Vo9NK2E0b2xc69A4tyAe/jwPq8IE1Zg+EoSz0hbFrfDfd
a1rioHEXC2pfgJdzrNMa94ESzZrTgxR1rQuIiqoVc2I3cFzdUDWMoaoVD8Z2MxyAfLqa2IgYb2zW
c/+zbPK5PqD7KRv0+5GYMdl0yKgavRdEZmGcfwgAmhFRDWYG6ywMvs+f/YxJJAiRD0WuuB6DezYK
Uqq2lzSKiJNDtw/zivT78NDnQTSufww/iX6u/Iwyabp1Zqk/yGjIfI9TNJ0QmkvrEzdh+OEIfMUl
QnQJiyeT5QT9Oujv0MpqpavlaO2Uu6eH4wzY4dKG7blIhy5kNTxUjHBP1bf8kAqcS7qIbUyhWIVn
qmIutpLO1SpHZGcQ9Lhe7ZWHFskVnnuh/d+0Ldlp+a5oL38UrkFfNSqwNdUh9RZYncrMKe00yHJK
3VvZGH+RlOFYRL4LzEp2hxCaj/T54tRtd9J1N0zAop+FUr98bN2gzg6PHKYbPyAwA/haRPvu8d0Y
WqqA0TCqlzqugMVJcixYHVzkt/9PEBSQ+MK1Kz8lBHybPqBqRwuR6lBiJd1nKf+VpLF5KVK8uu7H
88XZmk35UMHsOggpeCWZgAQLMRe7f6BFTemHKjuUYuzIR2m94D34QxxR2MpLpYa4U54m2lrJDI15
kzWpcYPdC++EkPrpj2Nz+132s0xGA9eZdrzmYz5DrcNs/1l2D0jnSrVjq+SsovObAxeHBNlOieLr
/AHZDcmJrQehbQuE2t/KwqHOipYF9r3gJRn8oDF3uyZktPZqHsYhM/WEPWoYJdfrGIjBbx78DzSN
oF90LEORWFsnGpsgd5mmxBwoBFd0V+mm5iYLY8A6gZJ5koOfD1FK0oOx5fOnJOCVyyA3LE7cK0bD
sevIU+e7/PUwl+qivaYOTt02Sqy7cMR1znHTzycwb3fPuhL/jc0v06rwdcXAENJEh9clc4pNWX1Q
QKyhgEj3JvIVlAauzZmI2nxkxdwEsXYnpnXTnx/TYtXR5OncaYDWLqaX5MUfrbduDH278ZtBReE3
K9JToD9D6Mn/BFYEvsRuRcQCI4tIyyP+xvfJKJb06F6h+DPWyKSgPC6nk84hBYgPpvhKPfZ/+UpB
YVxhUl4aK+2m+ECWgZow43e8driiHTdMMQeyoZ0T3C0uKTETOlyFfP8u+3S7Qh/rWTuuk46PKfTj
IBEeu1/QVumgjb4Q1xW4kR2U02/Snq8V49RrZpbQmECBjRzsjMFd4OgHtwC+Y6rEbSvpDRJ9fTbq
35AdJt4LYKgAf8rhhIUyrIfem4LF0vH5QaJSiVul6TFmBkxKbzBvuBEpEWAJGcjcOZ3cul9PM77x
1/KhLFSbxscAbe+bcdDImv/xFEf8JbMGzq08l7yFDntGHZ7wF3Cg93/AP4vrATh5EsOOtuCkTG6V
TwibiYzQ1wwUZEki0UPUV3oZb1dSIgqFOWV0WQfNhoWFdAv060Y1tp4AcYr/+cWvvGqSGcbDs+5B
foSrla+S4zFL1JPJa05N2DBzmCPDKSRMfKJdxpOB1M0oRgAw6ivaMK4D3fbUIRNp1vUqMGgH1SBS
73H0iEWMU8vq5Zk/igFH8gGJeOJoGA5ON+/7RZgulcnMkBywA8X24TXcJRvBxYZPTWiQjjgfTdy2
Auq/MG/lwSm8FXNI7TG+TLJlk2XC20UUdDuqZzXt8pbEx+uPFGI+nAYCQDJGtc+xmTvv5u2YHSn+
WmAOVM4ViPw8jcfP1T1CdBaiGHsZ3aAbdeYq/F8KYl9NYJHiWwfXlZeds8s29R/WQPfX3F2kdkxY
f3vWQUkPRpf6R/2yQdf0k7TAAqcFaiSnIr8NmZhUwmjSk3aoYKCh0ypKNzoK/C9uqDqrfUiUFwYV
phrZWNAp9bGcw+/fNUFaFKQO82aAONreb/x5br4KLQMDUXI8TRF//Um/DPEEcorpu5xyjOUL/DkF
29XUAfyEbkVNWkNRPQ6xkOvjO3p5psKGFSAU3Asa/OdkGg1JYGa8hzDuoxe6LIcMRC7BWkn4tCdT
ITPPmk+lUIQMBlwVurAn2UL2DyJauMKGNQPJx1dmi4KwuPGjFvyXqiNghYc3zRch1JgICDkQAzLe
NXr4QCtRYVCUw6S/Pywu12BgjRYPm3lsxMCIGp4Ha+0HVqquppYQ7w8kBj37fFFrs5cvZoABsFEH
50L6dsZh4Lvs4zCacm9hgrRthq3PQ9Bt7ckv3t11EtVyqi6hn6sWIxlXJnyHRN3DUhK4JH4pmFDI
HZUlJnUPceya6xsb+TzoWNcU16FrFmBD9YEsU47Yv+/y0IAvQb7vro0McVaYgzY5eEH4i0346C6F
EaNF6bKXK7F2S58Rj8kV4U4C6hhj1dGh5vdx+WsvFXK4bLDffd6VHkUFaUMcMLWGdkJpex/ZsqsA
3TN0PfPb/ud9OH6zKVabDCACel82TXxUuIKmq4N9nQ1akuuG/NKPPQOUiZJKR8aWh8Xu7Nph2T74
C6ZI3hZ+sHAXgGZabq76Vue0/q7WMUWKuhBmuybSQ1WdHEsb8+ve4kasgAweOf/dhUVD4hDZKhUI
YIqUFvVx0EKt8tfuTMGrz4oCAn7hnmIkkATQYL84H3YrnDdfK7bt8OYlXX3IL47mVlGlE8FTr6r5
OmFCIkG3MHurUwIQ56dXGfhS7SFgFawYSm2Dj/YCzn6V2zmU5TTKN70087hfpQ3J4rwzzoi9YU87
u2Fqmu0LkKoQSShas9N5uoQZNdikJ6gvmaglFfXsNNNtE4GdXNZo9ZVPEfDMyaFlUeDW5q+3wIWr
ezWTqvvRxxxZKYuNLiXX13TBJ2nQuPuuwZXQJFzA4FjjApKZne5Z8vRjHUq9efFaFCvSGIh8rzZo
kaJwIUdA+wPPtCHNra5GYvQZ27h+yFqLE/86FLalndy4+hXx46GH7DXthG8D1wnIyoaZfj249mzh
EAXY7tjasiDyktQM7fWXYRWf342fNfbiMRzzLvvuThX+l7+/WuXY5Z5J5nNevF2P+V2Rz2TGUTvZ
iTqllaiZDvtbCoUnoMSpv234HS1RyswjdvG+mQYvlgia2sec3tiXd9xn9JwpDjz0L2fxIQH1HnpC
nNvewelfW1soCMlJPM2nSPSRjlXRWmR/7w6Z2Iip4wAQsU1EeyynAMuFq4Ggdz2XKvFD+mwXpxKa
D+nMGGr6kSj59zfGpKS1fionnvAbSRCi7B4pRRgu9k802d2p0RbjKu5S4N7DJ/tQKyYrlatfQUjo
8p1+83hJ25X+nYt4QhpGlYWewDpKs8axOJSulU2BDcGJE4zN2tDKY34homfdaAM088VUqIIIhJCt
Q2rhpLFxNVlMtbVSkKQL6m44rFQWq8DMUyQgSwDTYGBpWiQzLi4TloJv65G7HH4dDeXOmwaobMQh
Q1mqjlXUOCenQuTeLfHFSEFkZCa2DDgGy4V1UAJFnXbY9LIDMdVaO3NMAB/W0m+nf0Cs7GTmb+za
ZAST9mPFrk2nSMT5KgmYVQhpAkEV6kyokibxdB7dWoJ32xmmnaKQKDEWuaU0MA5fhQfp0OuHC8FH
PlxzcMH61fuQ993cVMpWhjLarI9b+BqBzk9nq/hatv3PcXrliFbCA+eaLoTSsiffswV1G0MgRcEW
1fY/Js4j4fAqRLEJz36WB7s4+YPAvk7v7juD2+xWp053KH8PV6/bPa/yr2JZHH4x0+UQ2aNWPcXs
/8gdIzfzb3JnIuluLGnVoEGCF0R/b28rBbebZ3ES62xmnFO4LBVCfD0bNOcufYUbsVwg/PJTluZ1
koojFNroQcifng+jChaR14ToysKdunwh5wu4S3N5TPnhd1XhvyRy+K4yDfv7zOzRVV7Pzrkb5YFx
6TJy4M4ypIpfOABlLCzo+2fTVU27+IQxEDAL9iuBcF5fQETJGDm1uL4ShiJRs29s96Y0zV+OievJ
q1svIy8qrSP3a8CLuPfWWvUZZhCOxbYWpgJOUzaX576g9EK+ohXMsvV/np89rh3CgdiGxEBx6ZhW
jao59W14Nj7ClK9YeRFWm4XNmb2sM6txRZFJWQzsGxx9UiasPKX8FX1DUmLdB9g4dtpKYMsU/fba
wJmKX3gTXB12zr9Cdn6htzo9hSJMZwEN70S3A2albU5VUL+R0612phqd5OrxOWQdrXy8rOxVF6tI
2+EvQofyL23QJO1Lb8wsmpkwzOqU0tRDH3PXMCfD/Mc88xSoSN3zoopDtPt+io0ynEDL7zgIAaW2
JNwqxkGlZrw96K3y36lUtRf1oUvfeQy3qHU+w8NiJw1mWJeasaFACULNLTxjREh+Aiql4Bz7lT2U
NiReZod/X6mo/S6/Z3DAuDZgX8/BxsHCiYfvBpA6iJrtfFfR1c/7hYtf5mMo1+w9G5YBNnGVAsk/
MIIcxTahQ/nffa831UYEEZ2yrwuMrgUyBfKFQhKigFW60tdZS3hoPuFg6SGV5XvUlblLVA8I4QWH
gTX1emGw0bNXmgrg0aJRQWn//kDYkv/qk4c8qzxhiWh1Cr9x9S4fnmhUn8tSBDAE3MN3rFGj01oW
uIyS6YXqqOmpwZhLm1oVpzhvO8dQcd2Dg507vxvWyX8l65xGZvLARv5QD342ImTg272aTx6orcIY
fbV3UqcX79qNMsW9rbhaMb/31U0VsW7J7y1LBR51sCCCzW9Cy/EtdFHhNyIrAFoQIHV4BqjTrcKp
WF0ZXLseCKVDVnF6zg942C5A0sXXzhWmoQU08pXh5OOQd+mfGJiFKI1JdcIMdfvywqTV1uOTiuXD
/9Gpm/vAniaJGCmKEBRlbKx6SiomlbIgaUAsSDIEh+uB/wckR2nzEViaIwJVtJUvSUSKOkimfvR1
KXgk25zHs7GP3f+kFzqTqeGDs1JHKpnfvaF8+PlIysDIwVSPEr+54GJqzYQeU+II7stabtFmPpBl
8ifAo+W9oLKu7zI8rE1kXvx8N32gbfYsjQdJR81HmwBzBX/xQM5Yfade75WiX6nV5Y5nE9Cg58P9
28wT3woP28yy9HP11ML+F5aKYIUKc8w0IYJrnFwKrrWa/kiMsusbFlJqhf/UReNoQHhPVfnGRzc0
Qx28cdNoYhGH3mVerShl/ZgzGL5YUr+3Osyk+YGLIJhzSFv0pLWgTY+N9B6CpRuAC8JpN5MSUOac
Oc/wQgJ7uoEk0g364IIlwwMhDGtAQNBCToD3wwNr5Uh9Gc3amhwWjoRV7gsiEWUSrk+TlrUeDtUT
mmYkij5G6OBjswVAhE7EmlGLm2mEtUYLZt1zdCdF9cR90aK9iGQGE1alLkXeJzCxMyE2Jnq8TpZp
qqa2a0HGPZ7x/j1w5i0ZaivXpNsrUVHPAlduWYPkZ42L2QpYU56RphwWHRqX+HtC5W4mobbtX4zz
LQYU5ae9hXXCLxgqpLroqrTjkZMy8zRl8pyTK00OndBbXcXq+5xuU8KedZrUeN+rTK7N75W+NJbZ
mer95DhvFTyargXWGgT0bKPY4lgog305RnB8bhGBnr/N0Wu+AcAVX1epm1ZxZtaxNPUPvYq5r7pX
wcy8h1Lb70vNzPK2RLXS730iVD9VrhrbvRpZhhop2RF9EiUlKfCqMIoRxlvRuWB6Al8KS8pUw6Lp
hVvY9sryCQUkWqcE6NVuqCDrFT3Gdvuma2d9K2HOpMDdzds5UhI8jdQbi1PbnkJ20gnp0EOrt+Yk
1NSpA345wXzpkvZzKSQRwRn5kjK0TcHmY70+tOhFO7QGCuNQjwl4iTggNl+O6b+HUxr16M1/A560
Go7BxJEE6q6M7Vovdwx8ZvnyvMuoAhP5dncdGXHt1WgM9n+AX0e3C9FgQIFeT9nzZ/rbmPUJCnug
w3jAGrQXzm82D/myMqdhSNzrQ4HdIgGsxqrm53hmWrwEpQE1kY+DhJTnbY8kR9Py8N4d/ugAYROh
CV1Y4s9p9SdTq+TsfoIvtM4R5EZhTOdIp4mf8gmuFoKfsyV1y5ii21T0EdvG9RbgcEsuKVduraPO
dw7paC6us0yhtTXWcPVeqxWONTXvmpcixGq7qDFoix7xhX4pXsUQUw8wbizlzq67ES0mFDFIZtVN
1Z3rDpUmTZrYqZD0FjA76eNfSmBEMozCSmIdAD8xbrnU5T+qTflLRKRq/rGpISKDWfscF91Itcmt
RvtGSS6ar9FcAxYw21SqLf78LE3e34YZoLZXBkaMhCfBlU1PxnvSWnK9GvQiySawnyfRWIIDjFmZ
SVUDzTnwqkgVaVFdMzCmw2zFyPGA66HXSnxdws3GXDyz2JPp0gwv0ztpmX7Dx4TIgAL9lSDwYer4
UHE2QkYPy6MFhmMaBITmIlQIoYo3zys05EPffPQM9pE27jN8e4EXVOBcDzv5ez4SVFzubUdfAs1j
xoQBSBBIjh0Aug0dep1n2WLFKUVLVFcHeT23gPwB4hwgiEb9FwmvClnfckWeegnxJsZvYfThkKBq
BcL1ABDLdOu6hL8xlYvTMGW5XnrvmyY5vxF9SkXsYx7Y0qOuq07WngRbs8m3HupZi3WMDr+L0boQ
hqzBsPXhz/mP0LolZ/KKmXB0pNUqQt1vN+szLaDsKSrbpPYEpEJ8DtyI/6UWyrqGMdsqCtVMq8tu
Rd/Wg8cdkxkpQPrcCCpkJK40MssvVoVbPUpojetWxdO432YhjAhbh2nRjSuCcFMdkitLfHzpSd0q
ia3ZufyXd5vR94ctUc+8tQyIsbixZjVhZtznWMGUYJorOHnsMPLsAo41+HxctVDlQSLjr6bd0idg
O2y+DRzn7vgLCIyvyV45S6icXfwDeGh70l7MTcGEXUGSfOkymMb6ITOug8yaHB3MR7w6B03o8M8R
92eBB8J/vwglBNekbs7cWIkOps0+G8jchNAyQLRGxw6r66+EIYhqas0+6DTJGXZQRn5OgcX0VG7u
1WK3ZciMsuz9SFDxeQjPKMuPdCV6w5dzb8Qs5Diq5jwPZ32DGyUMa/nOBO1Qyv6L3Ho76zLnDl8D
hYoLxZ6zWjfEKFFb4mrGnTWLsZANuib5lvwnnGK/4BAW73BMxWMNSzM4SffAKQaCCEvySYdGPn+y
P9AloVpFRCN/ZlDDTUg6Buf1FSFbakEJnoVQJ1+t2c7t/vxOV71AXoTTOKLYFCaxZ0HaK9ikbzPL
xdxtG1zRpt+pTgVh0NyPf6RydP8QLUetZG7ISF7ccnwssUJfQ0YVOUOFXU/gVy2cfkwtQpfGs1tR
Y09W4HS9lyAf1IOj6dGkqyPWy+3nsu4jFS2BaVw5TshK1rIAxudEMqpns+63HD3NpFbtz8u277cf
egE89Vl/IiZdqBzlZeBz0039UckCUQM6ptiocYs+8tozZiXYwR8EZdcPNfTVMR1JMDtN89cbgI2C
+In9GV7+1+yVS5cwUOoJ9uC4dJE272f/KiKeGbHwfMKTeRA+oe8Yq3+yxDmcKEIzD1LelxLjL6xH
etE71n5H5KX/eGNr2ZPRWPWDR07x4g9RGTDmZgyk6pSplOn0ResKn+mkxY90Noqt1SvGmA0F/deL
97n4QDTsmSHNXjrEVPNDOk4WSia5tovWFNkDI22Yk2mjd2IF7xBW93HSt5JsaGwZ7+BQu0huzIy3
6aCgFozGM66M5zgXXNC8cwCocsmgO/CiSyLh+kuisfxgU3nxlTe6uhm1t/Ds8ZNMzL0YayaH/uBH
VyfiK6GcI+bQE15cCWFxG8oneXlk+nkDK9OPsE/AERN2fXhE6u3z+84CaJiLHjmlju3+4zUye3KB
9saT/Kiqdo+ad4s3run7I+DXdotoE1vJKTeSPdx8gFGydAUqUYkDEbtiJmDbvMqYp8AkKTpirsa5
faHNCqExSEN/hvBijfUyeRvtjeQ9UvwG2r4kB0ZEVo2yqB7RvOk9ueqRhR/8uAyCRJTJwVM/aucd
k3tzOBugCC2FjjwWv3vES41vgzyoajVgLiLGehBLJdQ0XB6xSMF4nzurhdVS3FMKkiWBDehywJ21
1kPYC66lE/zIt1E5DSl1qzMau9wO/oxg5oD65u2kBssLOewfv71e5NyxDLFfpxi3Y2G87NvvzixB
GlsUcI6WDeieTX/Qh4xOoea6Eo12w4zBGTEz5h7pVZ23RR/JYrKNLcNCyIFC7T+HN7uwu0RzuS82
BOylkUfqerBT9B+7fApbqS8ShjnA5aEjTNpzEdKTNuELz8rIwPHbTvfsyk9CIo6xvhLsuLUa8eeD
UAf563//08gHInIJUI/BEXeXXjQIbjtbZ6M2ynns7q+ozLoHKuh4Mo5gOgqLOIQu7W1XvdVk9xXh
ALitDVVADWtCeNzDJ4HVRqH13Me4HcQDYJnNqPyGZv0643Pqq+vCMylzdh8ba6AR/Mn5upEzg97w
hx2z/9U28fRuLs4wE1QioH7g+BxhX6IgOZjdhmTTu1hsQ3zA+bhQlELjhfg8BcIsK99ck55PhX+n
iNlzLKe+H6QJgv9TT4IT4Kje+ja5JCmVf8SAGd3UTSpCd5FiUefNnYkK4PRDSx8Vs6ZJigTYtl0/
k+lDo6b9OOAsGS7Gmf/ARWVbKntAyQhZp58OfWKIL1Jdq2M1+7ka6ex3wUwwTQ5zHwGniyOIXytG
OmPPqlI6EgSXudttVg3SSEFR8JD9ogRvlMwOLTraLpouNnpeqhDl5TMoR4ywCU3wkaKLLiRk5VtK
AXs+UZRCujKtEwGERi3761UuXyP0Y6TL2GMpy4wELPMaq5nEW0lTuuU9aI4nbL/caSZoVQqxVf+C
SJcCXl9z0FLJZbE6vWxRuLl2PfYJfqLzqILNPyxG+NbT/kFNvi/FP1yoC6W/XKdnP95R2J0356w7
3D4DTgBUVRYnPvlXxAYglTPBS+DJwVDcJ/W3B/HlWH2sGglPpVBzBqr8iCPAfMDf4EwB/k2HL8iM
AiFh6YJKa7IOpaIPT28xcnpMdXmInz0o4lfK6Dm390LzLI1vAgobVJgpqMJdC8AHdWQO3T9Mb0w1
TIza4SLYX7/9lgp96/HiP1EU8UUqqD3Cs/7L9lgk7eYhHwI0SDD/k8OheqMOsbHZ1F7zsNwsu7Yk
7ri1d+oyzhmT+mzL95lgUSiFdAJwzm3Ci5/ORkum//nuRpThCYJmSddUPU9K16C4GYaTQZUKVsHx
cXlpY5V2xyfOZJUJXqpyb0xmgtnkcsuO61qWcU5rwvm2bViEViUR2tIUESgvbhAUkUSEJIShIRFt
w0D0Kp+0ZCcgFeFqKgEt3cs7P6FJDHjsBTwbZX4wBwruD6ehhCCklqXLDL0zarXR4jvvyZzhfCdw
z3JtdrnrrHWzeJIkxy02dnilAuIWzaiXPbIAV+wxgEKMZXG0WILD4RkpjETWV9oiNG9bFctE5Dwj
3l+o7SY8AYpIGdnF3re/4TUeFmXehUikih+H4zGt1gxa00crnB4KIkp14mp2GeYh2XpezWeu8GoQ
g8Ayl3RKXaACaWCx3KuXrSDhPphKduDq0kD+ssSmBJRQ/EpwNUXQFc03tKplV92uOF6aHu/FBcI/
b0Y4CeXfKaDYXM8sGVGwt8zOFPfMfFiR2wpjVwhPWpOrYlK3+Djy3xGmfVApTmEEPZa1Vhi2+IFW
+C9c0N3aEfS7vAtWKIfJ6DkNdw1sG/LtFZkeiQq5bQRH16+H30RPGXdZRnqfghWR+ZYP031wsobc
Sg+3GubgswBeTAzjnyvEj7XLGfllmIVLTB6co0A1FL2CS5JvDatVi8ANV13ILldMhIysQTuLEx61
zSu0oUmT1pfjZ3U9BfsvH4jsvoRK5BUfd0ZdCsm2sAZccS8Lni9twAq+kGeGi6IMT84+W3lIW7IT
bcvmOv7GeCFS1gDbVZkRUPcpHQL8gvY2eXBTj8q2+BG+t4PgrUxrfcx9gAzCfi0+rPYOd0sbBlm+
eGgyLzAUdGXoFbPUYBq6oGlCGHM8hZcw+ti2Qy/M31ib58qkuQSxYl4zX5WXSTVsYNWz5koB84Cp
GfLwTlOCajVaXqTuACraXciLDRTsf6uvZXs55s5rL2U6I2lfdnTZOSWSNQaMlEPuuiUeg49j5yWf
GHtCWfGEeUYBh0IulcKx+Itm67NNaBKQTPdcelv1h0r6bxiEztbMvqs70dxs2ITwuA9XZdlr39Sx
x8ZjSOMpSnAr6jSM6JeZGkowDMFvk8akMLlevUYSs5eFfxdUI2+p00E3A8Q+PQv6AVlpOBepk2lA
aPwJdv+wxj9bhB2HOKXJ1HH7R95Vm+3RtIdYWhEOpUZl/bNVAhRXQobdWlfLoqNy+x3oE+Firkhd
8vbQ7J27JSG3YK5AJQejbBq4TPajUnRE1qjWsYSCNydkvemocInqZumUUXeK1ePd3Y4ui31Egl+g
tKmQGL+VGjMixJ+RdoFcSMqzOTQmYyBAXQDiq8+dv0eY9b7je812cs95xEqJ6W3CzxGvT56AlsJ2
+FBd1BTe4z2NfVflhFP64PbxvkiJ5tg238u0+1afQO2AmGXuOsU1uJnfttL6EW/MGx270QBON7qZ
kMTmTCgVICa1x+f9AX0fgDWwN4M2R+UXAisb4mUU8qAgmfrWFUcoswgWsY09cKFAJQTdDggGL6w8
vL0Sb9YWhD16pbHYmbgkpuqeNDnLrIV2C6u9VIu5/ULJdwCXTHgA6b6PAZRx/HPAGgX0qr7sShlA
4mbyauJskMopT6g7V9PIO/SULMvSGZtkMG5TQKOmtJJ8kBJzqeK3V6VAPEvri5RB5AgVhnsu8hde
wLaR1Do7oC8T/Rmb9+Itc4D7ppR42//2jbe98d9tdgWYY816NqxXg+GIfE3HaLH45fDUrP9SGFoW
eLnGBnzGfmnb1m/cnjutC40oPA8LRGUo5pOLFMwThJmfXLq8LqFLbuLlOpxfJdJFjE1XIAN9HGIq
wWsys1OkEx7RfvtQc79e4h7GNcpKHyfHwLwZQeHxOA34QJ3uJwvjY6pEIr00dJ01jwpXuyf8/F+9
QEqPeYgP08L1RzUmd3CnUQdyH3aJEjlvj5oyUxtp9kkCGxOsrnyLdCL6PFesBBQxbAcDFipwo+cb
qDY6tRpd6ET06BxSAMSkHEgul9FjvN6Kp8DSDkjtyIpFZhuM1Ni1W4brqWKA5rIygmRlRZYAWi2s
bTrtwzKpi+7RMK1N47oveL8oW35QV1WJKAbmNg+cYzrhAUlth7u510QysCD+1gTD1csIsrmmNuEl
j59BH2bfgOXtoz23Tw1zoCAqJS3xK43sbtOxKQxJEa/oa14PdZ4QMV5eH/2/fNg0ajNr1shAIXRo
7WjPAjemf6iDRLj84iVu9hpty4Nft052w4ZsdBw8COGVCeJkyUKAbA21hExQzMMAhK3Bo1FVUIwQ
04yUe3wo6G+OQ3PQlUOmULluH4y8UnDN2v+9rn2LiHg/LjGMpMSmw/3/ASWblK2Y3NZfPVv1CYBC
H2CP/J0Ml3bRC4fbOOay4crUL/k1mPwDCZts1kY+ddbI5AocujkOrNBlTXiK2XY2QSObJ2HB+pmN
DBfMxX1T6lHBt+/hHdc+HcY3AQThPg9iPUZGiDYk+IdwXz14lnrUN+6lasEmr4Mxwe4NeTkEOGai
efSIoF2KAequw13zA7MRBQ59FaguMxVb3FlWpyacSEjSScYjdqENWOpmLvyYr5STq8+B0k+gVil0
sVw45RoALPEqOdZX/SZs+3739LWMgvjU4KwpdRpiILuikqAd5X9qOHLAWLcpAF3ozX7qQ8XSofOu
WtQsoBOMjR4NkVcJ9QWxdHevnZYFfpjCI+0fpWYCZJpBNj+dyNe7FsRlKhXe+uvKU4edO2JNwDdf
X+o7EgHAhvrbgt+ldn3xRBdkLGfMXaiyRow+MYxy8Y9mfJ2t6IXvjKUKqJeU7B31ZO/yCzFP/B8S
kF3WqWm9Zd634R2QG3HxrL3kIH8KFS3Y6LqdtRbymDRoEH2iiBfVqUtmknODkP4Zmb4ipnC8QCDk
IETdo1eeiCCIjIzilQz4zT4sr08/i0yl+mppAiVf/3nGDooKLxfuDWy+1iNR+JN/hgIXO/cFoVuq
c7VzqJOnUeI9oKZOM/sEIHIeLEheyJ5X7Zf84HwPsbtURoesopNGEZLAwr1jPQf9niqHg7SJ4ny9
dIA7BISQFAiHcvrjVvVqW9bS3dSKczVWVZ40xp8jSxMr8epivoo9yA+nS0ZO8WZGVGWZrLi5ZQIt
kDcKhoNTdz3WITWA/rOfi1w5CGqMUeB+wlih3dRMihb4FOD/AdUjM9p8ZRRy2hGwDbtrV6FnpuAR
JPNUUBDkq8pmtsAjXNnSKDMN7QUJ/V2EDCcXZy6BooxosUy0s6XuzP+691N31tyIq0ZwQFJUu69j
0A5KukOF18ew85pLqM6+7xN2xqX0Bqo965Ti6AMCbvuaOwH6xFQVn0TQ2R13AMfbD0ha9TzbYTdT
Z2oRL11I8Osm4FlQRqw46G2nehPCOg71/7+OQv08Mt9YFyAeTHI3Ve4DTJeq0S9J+lbozCtjCYeG
BEH9Ul4C/kePI2NlURhySKX9PuZUeCw0JRJbEkd/9xTWKCYjzwvHeSJ+q8dBnHQRHP+n/Lpe1HHV
kmdQDAJUnhdPtAMCXmHN4jCQKv4PrRHa9kPwcw6MzH+cuYnZkzlUglco2pNMG4iRQsQ+EBjRocx8
kCSRfsR8qhUkKgLLKMrfn+vq27owlqitmVpM7W6m3EVt9r0pFNjg3slB2m2AFUEtz/t/YO5FVIOb
o0u/m7jGoCnRf4FrAV5k+shxo6DT75uEWe4IUtYPmOyNcH904gfvI6wV8EbxdEi1yj5b3YEbs/bZ
xKi7H+G6Ro7zLfcY+8MRm2co5SdcLRYaqSzzWrlki5t1jh+bRMq/dNX1OVVEQbrIGzSRsfFs8+uB
bYjiAgl3PmU9YHTAHukM1T9NnKjPru0XWHMB2r3ZA/ri2eljPIhz/DFPXTqo42bN8gsgjRjr+BWc
SBCgQ7ijNgrGTfX2tiprCfv9E3xWibdqvH9vGQWZTu8NZLSHHh++vKIn+Du7oSWHzQ4J5Y9TRc0q
6iXqUnVQDLhtTEF4k+e4Gje1T7UPwXm9u3piDbSLX48DQMdz9a4tQeWTTO+8qjCVbnMuetBggg3w
VFk5H1BE+assDCq7Fc+YvdDwZJTZ02RYBIySfHd31ibjyjKnxf/k+eHiXdeU1c+B9DkfrkCrUfSM
8vr1dMLosVwqf9O8Gii3JIt1Iy95M58UyVCnGw0hUueucPiTW1U8GYpjbcpoGr5qZLcYUnZMv9TB
HgYGn0PzpxaFzXsM0xjKRq5QE+AO8uaWTsQxJG79H4PUkEHLz9NH+pJxHo7lrRtdq7c1pBmrW8zf
aNCI3NxVA9GNZG+G4I0p0ChJvH0PJSwAh/w1SZruJWbYPrdQN7UcueioInxuZepkxzdm+zez/cZT
9TF1yqXK1NSqn66enfiTn+GyaOOGr8oUtd0io/LP9Tb38xiw96Zfrfq8YC6bWAr7XQ7XN8SBwpVK
tup8WbC4VzbVfWgIb4GaqE4jnl7adQqwrhm1+rCLVR19JW2n3zbcom8Z5zw67eq2JNpVlhnOulSI
g9+gFkGmaTcbuVLdpooMT2JT13DeSvck1lMV6do4A5M3+1v8xfBoPN7piP2drRvA3mcgDiqx3q8N
TgmLoK58OLpE2lD1wi1i3qZKwb1NcD7/myXLiz9y8Fyh+g1tWHxx2/j4vxwsKhgw6788jEa+NZYP
x+5KAHlNwdxGHOcLLkfW8BQKkxOGdYxIjebnUfnKgpEgJMHK/F8Jxaa9LnnMgBY2JVb+1ywoaSEH
eHEZ0/eafBH4YWZReW1oxEjxMfQHzYA690S+NkqCN8vNCQhmzeeURYSDsO649VSmqlQbmeN4PbGK
vaeAC1Nzm2LIA2YD/cZn9vECVlECyRo+fqxsOQH8M1bBYzcQgAEAxdrLnmdoMLfZKUsqq95uOzvj
d1DY9Ubk1R+QYmuVBFamXg8Ennb6PZKat6vfDC6WGnr1Nj4syleSqg9XW+HRX2NmtkXHbRJY1hnp
/v4yCdd3P4RZWCVqS5/ZbOVstx5anqfjE4ceZsadYNVHWmc4Y500oaaMHEq7P+x73MSSNAdBFxc8
kXdiBln+CVg6kOwtft8RGBCrstnmnnZMcJDbe3LKjhTQa3ahi2eMteeSRYqM6ij+93RQlnDwCfdA
FrxQXb3baC5mEAyZ/NQOUD0VI4v0uToFi+gybtQdd0qplrNksbVD/spRqX855D9+XHJGadjXPjxg
Oc6d5PPhSXBR+YH+naudigE6QTtJjHQ4241ao90SU9hKxH2tWxIGZ8fHQtIX32JHQ5ONJhQwGDgr
e0jrfx3d398ZyCQjTad0t8xMOMMGAzfA3TxB9vwvcgYHXCZtZXHCTpmPza5r+mWWWrq1Vm745nko
VUOqM8Eh+q/dJwrgAz0n06D/2FyN9SSz4E4fJOoYr4qbKrFcRWTUHLJBa9euGAF+J8XHBG59m76q
FygX1do1j5Fqj6s9NSWgTXggALHpc59EvfH8Q8hNBOmVY2qihVeipun1omOYk4oNZDu+/9sgfOqE
okP6AbJ1SMCJG4jI2W01TPZI457LnZoAzsd61stoY9QV04LljJGWCL4/oJ41xbGEgQGfr8axcgKI
fU4ecJYGWZCbVUIcoKldbGH55NDQ7ymknd7lVxM1uFwjiLqewGwyYiKIE8BDfm0tBWkX3DXEKf8P
3JBKRyru2T1aYTxMFSWUmCqY3UDuZE7h3Pdq8A8FvrYI/LF7SyAt9jkhb/D64xQ4gxC/jEfaPV5z
QAbVkbdRw/rlrLF3KvT8LMNIZx33YreUooH9zv4y6HUSaIp6F+q6BIkKQtqlQl5OpjvfR9BaMnjt
v9iy6drrN3lR7XgoC/7JTcRVDGm/UWvwNnes8HjnCYSymjkXH/PyXt0dfGE412EzN/dRhgFcJ8Rw
UOWS6zrntiD+de1Kh7PZAnQ31YHeFWffmG2qrm4pPCWoZxvEK3WP0+BEGZetON9rYXVnghSf3H8b
VO5UMd0Ec4i6DNOJVaZvGCxVA6or2JF3gdWLDz9pgBkhZunDYLACeNDt4BwnpY0oCrGQSck4ARVF
wyVQdmAfCPHAR5bH956uCyENVgBjiu/OwDa5tQvJoU5NmQEtHSpicHFf4T32COtpteaNvEia45Bl
p01rduvp70yQa0+4063evH0ANOBThsv4WfP8FCsVJgeS3YCa7MXXMAcXMEJC9YnDIrebHTwv6rEh
lj5Jj0+tpMD9fIhRv6m03rTuFBsHL98AX461vFousOuxyUdW3ZR9KSByhfkfcaBxOgDCipYI/DUd
FiRodxRzGa2IVRe0k/nj05/oacrLYUMw2fDlBcrNNQ1cipc5SgJAk+swiIjyXjydZNBguWGbKmnD
LkQRNZwMkUgtBzt5b+8chHZbcfnk6Rdn5gK6TgrMSksUxyc3aiPCAY7SMI4dOA5noTRAYJtMARNF
CMRWtfbNI9Np4QdNy5cFK4k1gEda85BNVsDmevdzhPS3/8FZu9uIxBL7h6YdwbX9moFo7BWzj8WQ
ncMTAhfxsDFnYHs7rDdj6eY/Mez9q/wXdJqrqHnYSLcdLiDgFszt5iS+yQzNXSHU3ZdehbduBWLQ
rJaqFMfDlmyMZ96Z4L9SoGXuhlK10SVwSAiaUl1J9HVuCYOe2qszepM3GdCh5u6TVj0kEPIYdzP1
CtfCDLw0oD6MId9yFkmiNHzjEzLbg7KTKQUhVz0Q8Dn0Vy4No0XYhj0XeplGvoSrBghMeX0W9fDx
hzEIeASZbi39cfe8MXl6Czy1ICdqvdM6UNCG6MhLJH2DT9kmFuAEX+mP0YAkIZE3LuZJhzkBVW7o
nZhq7rkMKsnbrBQ8rxpydcFuU0UF18XAf5OHFcDEkD2MwVtmJ1M0NmgAChfH9VIkNY2B/IOMvXOG
7Rg6rC4qYEAdFtuq25maRgdnMSWANvy11belE+f5yyg3je6RKtb3+DJkhm35UotruDJOQRwswgNU
nybBbum9dsBFjRaBf0E4JjHnopdt0UV7qhj3rCJjfDHPauQxSI0rPGHDL2NL5Yfv4JAfpq2JgC51
jO9yoemMqTXN1QxQ1F+m0PlU6pwzXakdw3YCXlfGomXSeDSKGgmYJT7ughrhlFqT64W22lzgOx+f
7YlKGTcFmKzVVP5ZYZKulhXG/h+Y1pKgfE03dC//HMM1iW1yciNA1Sr/Bram5NsUfnIlrj2qtUFV
RK95ZYAJfH8w9flMVb+hXik2nA0YkhJrszTS0i/HSgdx/7sSBqFPo8UGB8B+xqR6BMASAFxdtqqc
ODdmGyEia1asOlDy3dufGvQCfzxgVxe4kDgRyJ1OppuEwa0JpIw247qY3GbYJ4R8Zrfv37dBU/Ww
vXIeJqWNG9PMCNqbdkbI1jx8MNJtNHYgYkNeQFguVxHJSTCTquo5BnSBWlkVpkpWDYwpVLWERdu5
0R7CQjwE6Zaut7rH/ZhoRsM0JC4BK2x02hJj4yKugXaYRbpa70f76eUN6/vMPKYCd9kkxkOj2TY3
Ul2kN05wjl2jQC4H2XrMCiJfAS0jatbjVjo/iNoZH/F1MAvHgwffSLvJrQ+ePgCu43D6SvUYsed0
1Q6VizZFAQybDMxh/igk/1i08wl6WOcIUfckJ4c8kQl9NQ8p8XnaWvN84LtjvPCHV8Y92dUMOF9e
/psWm5FjR594xIeJsQD0zacfGnjqPoB0zqRbSQKd9QNtrHm1zv5pvX/jBPkd2pIutGihLpClkdwy
FEL1s6Dd9mRKOp+sj0V2U6+j4tCRjzY6mx9mgVzRUjlKpsgJ/Q2obxoOpyD2GJ4qYjDdum7WipVx
7Ej3uicKAnVgCFlynx0Jb8wTsIh4nZ9mfKV/11h7m6KQPPTRO4ECziv4aZ5DDUSdzmzC6PSmAf6R
ygpMfkU2sYeTVBMtTIVN2EsGhkRABS5rtn0TnIR1SRMnaaqB7ddcKAijVd42O6qXaPsHOkzmTMwT
RVttjqDeoEIGv/EYRRDcuCFBpn7yn6reCzU4wohWShOx/67YBtNMDA42Z0LTfcpVGRQILVt3kyoC
3rE2ZvfEIwB9Qp9spFkm7aOzeDZ/24MAhyyJ47e9TTL5HZqAr/3AphnNwmbdd1fbyTiGXE+QokMM
hUwliTojlHQs0AuraCxB5JyWuKG4nVOBmCYu//BttdooRdBKAA4nmQhn7NVK8oJztsBRZ2AVKtDy
Q9TdDtGXWuJ093WCnIXUiZ9rCwTvA7vbOlGsRNxxUc59PuWBpR+RRIcvjrI4I3fv0Sq1tqxbZI9f
3nHfxU1LX1rkmnR7P+cjMQvbouFFPrbEpnoLkbj1mEFDv/dFlhYhL44BE0veTVjCR6AqobsSENVF
Zi1W8XBEwWi3vlt8lKkji1YVWJmEJnXv1wXDX8oTtQgs57Irht4lthsD3OF5hdrVY6aVQkHsnPwb
9lKLm7q78948Rs7HnFbEkJ+Ryqk3lRdHZjXsG5Nhe7qLKZ+NSDSh8vWvhHF6uGmzBShTISqV0u5U
ncN4rcOALE98W5Ltg3ACe28pq/5AxTEa6MLDUDNbZaTAzq6kk7gFkStRI1/LCJhiySI3wlx/ootM
ZYQUcPxfDrINoZHeSADSB4sGwtvGlgoz4t/4wdnMbjlIlwvau99Mob5kao2m2PeQW9bjAhQQJnIc
Zg0PkffM53FlYTWHJE5Ok1goAbyNQV0whbW+lnycni3Wn0RB9y9HC3gng//vNDlHk5TRa2cb6DOA
5c3i8l0JLmjImeYZJocu2YgGrJx/AdPBRTiRq7YSBKxmzMYK1nAau2nG/v6cjYdu701oXddXcX9F
OR4BQd9yKEGdFC925lq77dNweX85EvXxTH3HvW9k1a/EeQaYZqz0TFTyfChWborINdM1oQUHFI0U
XxW6gppa8LgpTnwkct/oG1WS53vyI+KyVfPoMSCDcc9+as/m02menDQnsCFKJThY7lfmvPoxmm2J
QYHohf79ZuQfUlV1Fh9FMyx06VNWVyMB2ljFewp5EyfGoZyytTx0peYqQcLox+OAHGiLjtNASDdr
StoZaRq+U4ETrHUVVtJzzS/vuAEeBMYUWwpZRWNp/f8E3DgqyyIehyZXgKfnqHEJ2FNowwrz6u61
WNeAcFWidVr4s0NS2WZTFlvCM+uwSTy09THAZ5l1s/DzQMixoDimbH5DMXg5hKIaDYANu9jMrAIN
jYwbhStW0knJPGHv9gCVSl1u+AcCKbUjfhoRyFy6GtDYVkZR7XMVdoCFSLqbwAeuaFf4kDxdcYgj
R6yMlJMlEoUliCmjbijV9jL+pZbZeGFqSHv3uDSXjNK1F62PsfmcvtHSW2L2zSKQ69aCkul4/eQp
zkEr4HpV2zU0g6Ejt3Gs/+vrNJ4kVuhrrBej65YNkk4P9w9EXUdirvTtA5LhdY41jHd3FGZ7F9tb
d2Y2Ci3YZ0Q8227Tq6oYZNqVBFNYX20ENcDbIhWoJOXyXDWpEjr2jVmRG31Qk2EO9bicvf81dhmd
opQ+rs3IwbDp1yrm0mS1mad4OaOkBdzVJjgY7mkWF19lOlElWddo02Qjc9nmE5QEbiCcaYmrkNfP
KDcRkFdiKy5TV2Jwt9PcHmg3doKXv9liAOfs3hs3513D1p19FqmhcO25g6CX0Rt+Sg2fD6JBqlRB
sYHZ+ZtHpFFzxPAAyzWKPo8y4fY71ZuPAq2vpxw12VB3UVJ9Qv0ZZnnpiLyMKeetrfTirg45IvnB
MS0qsoRfJwUbZTOMZGofQkmcTsy+RsD2gOWVMMBONiJRtUzVznVq37GvdAf6HinFXs/htEG3KeD+
pLQZRiT4+GEyFOzJTvncqfwu2bOHkN2x4i38GOks0v+8AoSv3u/4fxxvlj47TQ6hIAOdlmZd+D6T
oCxWagnk+j7sl7oen5IxnEAPjYIi8NQddv+mW25w+OcXwdnJCD3CJwAL7oUntnoTQ6GGnlS8pBri
btwCgAsFGHC/CAkT1FjUeasHHN8sSL0bmQJgRUPrZTctxAEWGCZMmKxKHMtclMHoH0DbsX/cqdff
cdCztyG2Cj0v+btydWq3D+M4G1V9b2oIQZEdVhjyLSJTqpw8op5kRvQMw/On4AHKFsnZVtD3hrRl
Z6sTGtGPpKEyqG4uvAXBu0m9JFfkM/NdhnOj7PCNITU6la3SbduD1D9sOINTbmIV+ZywXsWBlkg5
+9p5AoeMDoAta3RFaZ3NTNnmH7RMR7ZKscJPSYEJSiQMQXYBlxEwZm89kkwd9w83qn/EZvcf42x5
JDsy1f78w64xc5VtQIutggA+eVQJEJcbg3DaoTrYdUi0kG45BpDmqle0eYDC9weiIYJNFIG4rzPc
yHQkSPksvtOubVCG6lp3OVo5CGPjWWKSA+jSVvHQaDp3tDxODUnq9z34u4Oqx7FfYuQqoZRLTDFF
SJMX+vnok5S9FTBoiy3bBPO1LzVd4FS3qWHrQV7kYPZiBQ/KB4YOQv3TLEmri/OMQRcSri1kEJVt
DskAij393d8Ob2y/akEgXDsuOdGd/j7x2VB7i3chmZIUUp+Y4EzgbdDkRUW2f5XZ9CCVSbKFjxb6
B0DWU3220sFmJOI7MrnDWDA0lcs7D0aYDXeBvhaCdZ6U8h4JDvvr2L43UZFmxp51x+OlHGl5VPiw
srIXTmw/4ubw5P8eEu7/Qk1XhWl5U0+955LyB36d8jPOjwEvQr6wxmJO1bR4JkX289saARhJpNC2
6hjsN1cV/qph/RKSDG1ecinGizwritsHGlCX9kE4AknpA4Y25U63D+x1OHwwhCejO6UNR765OlCh
SWyc0ChPMBtyhQ9dq1aJarVo6s7XntWbj6RdQtfCGI1ePVNDdIlQsd0rKVvJRH0Sj9TOtSZpRv8E
Jp4aKpotndIDxecC9uv6E7tZ/ZTd+XnYwigVRgLa4Hy6FU6XQLyoOJLYoa+taC/s2mKiSjJQ6Dd5
j6DBvV1rHWsIZyPPzclOJRELvAM41mDO1uLBQCyeavpg7x8Wkngm4MEo7sTpqzkYjgul3qaSQySB
Xetn5buiCH1QRRWYLXyOz8hZ3Kzc8ZgiqmePiGEhfY5fORmlonA6zAAuBb4kZ0Ss+NGtlFiGOiWG
6A3cQQFV3KmJdWB8ekxU5oMQg2t47c9Nw+hvrUwZjsL3bCtEf+hhd6ZrTewYkLmJndp67gBRFVl3
kJOatvE+DOk9i3NZFG6uDFO+BfQfTTwfaavzIIaOxZglIOjq6xhIURUCHYTKCyMXzcfK4k+oYnqh
zXZGkxOy78XtqdAR2Tz4NUeRfRnv9VpP/IdeY/5aYHHU9eWF0C5W9lgbGXGIa3O4qXCYY3gh1BBT
ybuUIS5PBTfN/ePAWYmU4ziaR/qfrfZAdyW1KjRQ1/HPb6bSMt0xwSdZKr1JjVmkI0J0rBEyfWBy
29xHINUHuFrpooiCXgGjSvwNKheMNnH5I7L84TZ/fomvkj4eGrfuGIFUo/K28tztigvDM6eigt9F
0tBf9Ec8qZ5JuUB9nU2dEpTLxvC9FxbycHF13dQof2ZNY1uLA9x0/2PiWpG3iMVz2SCQzmi3fVhb
2BzUDKpnsNPFAonfwgE/IwhkRa6QPNovYFSMvPW1ZVX4LaHwlukjqrrSf965n1+DdNnJB7mRRkK8
pXKXEuCxPSFOOUt1oHfCjLf15dp29RR+8to64QEAQz7p9IfxsWcSpwAksrTIMxhL1VYzYF+hU3G6
LJaVn400myes6ZqslnE9g2oyCYp2zi1P7UI3WITL8m2EI8HEeg6WF6FMUmtB5Qx4LtdlrQ5flwEn
r0FCIVwaV1MBfGHkCIz9UZxrlA2KYGlj8pUHQWnXNtlAbVHGmVKTXTHx6glQoN/3IpAayE3E4xmC
1ClzjXkA26x8ciVPBn3NmWc3hwbwNc5Jkb303al8/Up+nl132UiW8RZNCWSqpdm5C7pMJYDyJ8x8
iOdF3YVMSyKDl0f5uQZepnsZ5dIskXbUqHPKYDQIWvMs5V7SerkcSHUO6EOusyImZsfknUuCe1UR
GMeCt12auNaVrFxzrEfW95pS34gojE88K7ajoGwIto1It8vO7uPJYaLo8Ga959k2zZLBMo2f9Xo/
+DqxX7aTtsZ/+k3PiAjfImKiAIZAJ+g/VSIZZ3UTTt+bDXrw+hGlMmUikOwpiXx24ivjGHVCMwhS
YAasC3qNwgntMGExB+ATAYVGdOTVdH9SGGUyRYZ/RyORYTEjCG4K1b9qnzwJWux4fAHXb5mZeTj0
C20mjzFt64JPZNI70uJw78uXVaHzZSkPMDtVuHNPxhAcaHXNEVb3YSNcv+W3242B9BfyYz1qOrnj
vVwUS4m44K7OyJN4a9ln4k+914dX4vi6oq285rVH7z0wSpdeT0us4Yw9AdLxblkY2ZGiAk1gP0DH
09mGW4GFh63YBA8ZGUd+632XLtqss8MC9jnlNuiHSm4UXN/O7XZPktNSXzShwhshIQVr1wh2qD60
evyPoERb0wnXSVqQtTx5gtXDsnH4gFT+DgrwP+OgN3mROVjRKFUqXKCUoZabPmNUkQlN3Lbj4tQ1
OFAdw5zRWpVCtlsO1Z9qW+5LL94ykwjGjE8DegrqLUpiMu5iRpHBxO6QsbpRKXhn9zFt82oHWokQ
J9BF7xhu496w6ND7YYTFCde5SFsirnJo29jVzLTeJT9MYYNfYXj/S2T7SbOJvkRwLjEZ7WaBR3St
aJh8D5Pz9sFSHmG93lbNZqQ00Op5iE91vCRTraJDeUMHa9fae5AKJses7RpOMfhvWKaeBkdbHvtp
oK15gXFWf2Nak9aeoVGWH9Fq2Yf+PNA+3RLKFn4NsY0o47WQbudChMktLMkkRdVdq1ey9kUGKXuE
5/plNse7EsbLfb6cjNvMn1VoEfwzbirYczTR6T/B3Cej1oasrLOuZbV37mlcisvIXxJcAREoigmW
QNEGGyUFgK5hjBL7pNtTA+7869Y3f64iUf1B0k0S0mPnTEQtTGwFGQ07IXNR5bBCtW8Y9SP6bN0Y
Ctas5hme9tyrK2CQlYGS/m1JcF4lc2zVrwJ+eX/fzJQwwBuAVNImBfdlRoV9jXNJw899Ono8iO+j
X964SXT8E4011nMoexlKG1b5PaArPJZi+95EFgHGMm/4VIlDNk3QQt+eNcAEyYGZAsfTBANffCTo
Nf33780GRbOiMSL/h4iPRCvZg36dDF7zZCQmn/ckH1xtQrmFqncItmgIncQZPeQltNyBaVHNm+t+
1bxAUUFmaVEfzeBFwW0zjN+TsTM7mXZEzR5Ob94UaZtj4tlx3gVZfvPQ0nx55j5VRIhfzyDaCs2E
Vqp/Y/LZLDcPjudz+PGbe+Z1kh/K8AR4bfBUBek+mekClWWDVJqdz2RJwNZ72uDC7CgGpn3p1k6j
FPW2Q7v6a2J4g3Web1UbTMMN8DursHjN6nl+N2wPDPOZx07rWBmoejKR/FYs6QJPBVTSUSGPxjWg
HjjP6EWGpxoTNqd4wW2mbH975pUojd9ZLtCQ7QiXl/KXoqZYVBQ1UfqSy6GO4zvRi+c6qW/ZniNB
j7+/hkAoLCiY/WVfVJLVQFZ/MGOfyN1uuzRuAipEeH97koyrjjTbgIIsmDBQAjmlWNOXCCIGHxLj
Kbs+VKX0k1wlGONyHCqXi7C+8KidJ5CnpBri5SO8E2kavtdTe4uRjyleTZlrfqestDGm7aZ+RYU0
3SEpkvAdDLKjlUn01JUx30lEN7AyRwtOjoy5Y/o8QPzOAwn37deJI+zBWssDnZWv//DA8ldE2pDe
puDLu176ljmcBx+84coS2lZdeThFKw0JJQDY2X4U5hUKWmLiexcB5jYOURrwqJ7rbbD5+1edn/28
t5Scw5zHNorrnELBUO8K9WGuZWNHvSpgOMi3NGHY0uOuoyrLcPQLgtHltn6qeJRt9WjaIN0DO26c
rWHKBYjJ4BSLRdmNo+CVkvv/qJc19z2Hj34b2aJCClmyP0wspCCRLPpMOr0ZeNSnXEFrmbsyG79I
NHVtBXjz8JzZbtE4PX79b3k0EdsMX3dwPNnLsszIhQ+UUcran+4wBbAK04k1TEcDHaH1z6VN9F6X
us7734p5yvFhgIXkv41OVMkHz0uJAJ5IOrdhF5s1FDGUHQbHv847cfTEtphQdM8F/07Sgan/YT01
yuE8DZrfIJR6kjzVN2Ih9K9k98MQci611h867ugV3dM4wI1ANQxU6/9AiOqYx9x/VVytfQyrst1u
QbIqL6SX+tk4qqkgy60S3vksgXaObA4Uk3XTux3npHpc4r/5VuyajtbBfvzBt0LCRjUxeqja49wN
TX3WbrfX+X+OarJN2fMq42lO7n/840MqrMm8qCRC5Unl0ThvhjVDpSR3LF6faC0RFepbWTeOQlLc
AcCyl738HpVGt8X+a+0BAnKZrLq9wtCjOD0/VxfsnncIoTWbfU6i7qUgmniRzEozsOz6GmW0VTYA
HbwIzXMUWeL2tSdcZmiTWXNjNdBoYKrkjkdQZEHkGAvenSMlgWypR9l7NoJAmr5Ti+5KG4/xXCNi
cGcBvbMKOOkYXEekEhtTTgYs1JpXJs/KFqFpYJg9jdwW+QZvFOqWlFJyV4cRLKZzfzf2fxIA2uiK
gccJZUfPZjkB/VYdUo5NdLRD9fiVZOO2f1dZCj2el/KjHA3Gixu1gU+leNxR4n5W359mz5eaMOoL
fOc4RUpK2UnJkBNvHlgNBfm7eVVsjV3emR1iVzBbYv6zLtH+b/DNHotPRRwBx0RlBb+F+UHGr+uc
pCqO1DPMpKyNW4yTnO+gZ9HwDDyQ7RhfGR3n+V0vhq1fM9nU4QIScXsntY3gzqRaqBqe0/NSpTDX
Al96YGm/q9zLm4ZoVta9SgQbQtLAFTM1IS9Dljou8HiqbkdxGPFau5wsp8oA46K26wW8viWSbfs+
mErChoS6piMytyJG3bpW8C1YpcQXdLlWYW8HT7q5GOCJ3KTFFUE/LLxf03sVXG3hak/DUDEPGV5P
IGrrzkUi49QELlvytUvd493qSCuHNJnfgpJjDUSHjJT8wBPD23KpbPqqyRbeWF0EwdiaxEX5WEn8
Z3Q9AbNQrhjQzZSZR54P0HwFVnvqryGkNNbSu7I7G6+NPa2LJAPID0kDdY52OXs+7qLXzatlX3MH
0wuHd+ZwIldDM6HW93FC852Ea/88RsNRV6Bn3hNxIL0JxiqkYFnCvZNuZufLZQOkBY7tMiP56AH3
fgFiCGw/ScrwmFtOTMv+GpeYNFa6t+iwZxQgShLjGO2YKGs+FSk3hGq4TU06Cbgx5RwnB1T6KsZJ
eZoW9j3uML4zPYj/KeHg4PAVAzb4gESvbHFThSGbWxE1zBvTnHm9CPmlTBBmDoVhPDYH81kwSqjg
E75qZrN8j179IeMobDaLMCKStVYP3psVUxDF706MkWxBYNuAvdsargdnLpodknPE7DJl9zkSvJZQ
2H6jo9lRT8RaxqXdFSlV9Rc8p6IUlquLWx9oo6jYbUzU6EfrScdTlsPyIBft6ITWyyvohF+zFE2C
AoBIVmAqqyZsgT0EmNhYnzqlUeKEzPyDlOYtq3yYEJSDW9GBVq69geZgc7mjfW0bDdL5SProEHOp
DohgDSn2gjYJZJNueeMCAwyVSmm014Ec4dZtF6EhhQUQAFxBPH7sYJIlbjh9X7Zx9lGXg50UbnQs
7sYkZO+perdb+N12gyslp68KvbeamypASoDzjnyUcdzwkt9ygnfnhig5mBIw9YLMkJ7ghwA5TL3m
jnw2h3Mpa5uvGjKDFquM9qSC4RE/ruZQtyTk9yycGBTtGNptOZFiWNehkuBO/jAxNGl2TSKMOY4t
Sh2JpzCn1PLPzhAEwJNvOkK2M1Akk93MJcwkQ2I6ElNn0Ka07PG2LRrEMvHZnSMTBqKmxDPWbISA
Ti9RtP3PSMhcwy/anEl3wAMPkhyfLNEfELeqP/eM3/COWXHjwNaYvCAQQjcHj42gEsnSkb0BcOno
dCD+NhvNMqM0rfgY8LaMAvX38BD+PqEbVowlS4WX47fRZvGEeTq8m6xAI4GQcHLEpdZ9Er3Axddb
v9w7j5FuwyhomyfZ5/uAIHA6M8dkz9u48GP1zAIyPihrCxScTGsd2y16EsFeakoJbYfsn5iddmJB
NAxs+J3VYblycBWJzxPRyLUh/Xb3OnQxvK/CGRTJHttg2lbtIWPcYZ+44PyFIpreGe/1P2Rd8AzE
AecWDOPIbkZzt/VP9JJji1srsTACloATsF1BfHVWtLAaI9iFWVw3aqusTdHFYYifUXGKI2FSEb4X
64IqsR6cWWIYao4oUgPKYf9cd2ULrixrGuzNwB7KnVM/20xqsQ9BYsG6rmYh+qfkXZvHLf/cXZ59
4ayGpvXtYwTgbdN0unVIV6i6iSawU2a0+Ybj5gIEffEnAWzfO3FFfIogAyeUoqDEoDYd1k8qPGZC
i7Om5uq1zfXPyYbMpIyBcknqFrhpwaXDM08sJrLo5tKXFs8Gyukvr+KzL7wgto4ph4wPpms2Nfof
YRJ8/bQwY0+UD1gjnyL/+yIxXceC94coqOHAdHZ52BR+/C8AYFuZpL/Rmq7CkcidfiweNSfNNRlC
xxqvuW5OY7lvtXaq2aGxD4XAj4LTksTPQp8tGZl4lF0NzcXm2MXKw2bBXuhhTxrhfZWzu+SC9xnF
psWzhKYJj2qJCGC6cEhnym790CsqnwrYklnKuz6UkiZf6vI2yAl+UVcgKX2P+CgzFtgbxxAbsR++
ouaIc/qVgaPr8t71HQ0VVK2D+m7UJw/JXJsG5mjnyRXWlz52JR3F0yRy4PkB7lOoILLYiFfRK/GF
LJjK11bTnnHFRygDPh9mjg8orJLkn3+RykFuba/xoZ/KJHeqHGwQ4+kc3w4RGrnqm1/wtZyEf+3l
WmqPVoDA/DkJOWCxTWV4Y9Sghc71Z7/zVvUQlcDl+AH758ZHqcz7q9t3Td5S6NY+nrypxGnwUYah
OKdEXuN02RwZk8pmTRmaEHRTu/P3nwz6HyiKEvlC/WOtDU2PbcZJiXcFK0PL0dArmld4LrvWKsI6
y/o06aLHsIBtwE/1I+1ESuGe9gwwHBslejU8QiWQiFjDZaXqzbkSKeurZy6ustwWgqNIGDmPmiD6
uTAk5JQXom4Xv9WLH/qmY4uyqw+sj1nB9czEl3kHQSTDLuVONCRqTJpnpNotxOvvskd7VpXh4/Mz
gZgCc7hYwkucUkiCwOl3YRHtphiwqY8CTapheK8KtXBFjdWbsWt8JrDgG70UDJVz47LVhxCwyYCx
F11bev04kRDPTnB2e0PijNF2Wp9DbFKJaaIDcJUl8fN8PO9hnqUVMNBNGC1pFaJWXaurf/KNhLiB
mPCXh4x2DoIs+dpXHvuuA44/2Tz1v+rupjxUVeDyEDb0tuqb2W1DH8vUe5dNRpVJttsC3JuqjBul
LoSVkg80JLQ5B6mUB8od1Tu3thJnDPmEv+ukHDFqxbcIpOgm77x0uXNRHaKzc0hIt41SY/xt4JHu
sjk2PvNhXnUX1Y7MvN8yjhE66x1NLitI9+OqCCK1/oA1qVrwa1uM0XtaZbAfR0OnjQtvFFR9dbuF
uJyelks9woeOIGjrPBK7KjgUwl4CFfCF66mEVxCQX379cfPx9yiiWSnU0EjcXmec+9E8rZOlvHUT
5LrT0S0MqSldVQbgHPdIXMKiJ3pMcGJ+5xrOi1moQzc3TTPf0S+TUO7I56T+/nWt81VVGKvJO44n
Dh0wdFBf+kmFE4K6jM4zfgZ+RDzYsaHHIsatzsWiILm49HCMT5L/L2vZk3OMuAVuSDZNvyDySOMO
ThcphOBZDD69gHjYYXWlN6KXfmNm2R8cVn4AAgPhQTZ2j4op3yp8f99k6kxnxQI+AGmYmiItijX7
ELFkza+27lRwiQRzRJsg9o/bkJGOflauGPUWl3hVEW1Ayxod7frq8ajyYF6cDfM00aMl8hmhVj0O
SuXz6tvuqa96MrcS7OeoPpzRHlyZs/ZUm07YmVcqYM6INHA8xHroAvaun6BImZlTh04sPqNEF6oN
KjZdr3nO2AiAhDA21rEluXGTR9mOrTp+xCFovouGtbU48kRGdqNKVpXN8VySg6L/50K3M0TJncA4
BgatH59+jthCRv4ZdavL9fp7Znskz+Xv5scuzX7CF4ROOiJoQHK0AkPiOwgogyPJgYe+ClDz0b9i
CUkCTkQ4ns9GrQDcGzD6AgR6Wsi+ycErZnVZ9oavKpXejVDx+O5EXya3kA5EfsgCGRhD34GTmK3I
63zOXClH8ylBJX1GTybZV1OoxbHhtCauJG7Mm+1Algw8TEM3eihNi313UVfPQpVMJzEAkS3YA3m/
qTmLg37txDMquvnzyRXEtHPYqgjNscl37tsholRw239i8wpBV/qoM/2CMsj1oBgO7/IcEyoUFQRE
OFKiaNJmauNzt4E/n8OQOEhfxlhDYlnE5f+7WmyddofSBPRo9WrpCq85igkE+qr44DuY3iQOGGy2
h/TBiGBC11ySRdV2K/ys/evzbz8O5JqMwSPqkYmKux5cCm99834dPVBsWGR5rfaZZLBRY4dbcFMQ
H7RtquGUmNtoPy1IW8HNPhgN6b4/dxSuXEyAs3p4QxTR5wWS2LJyVdzjzYLbOrnyMcSX+GgJmG6N
reA51Vbn9ad4Ny9n/h4uouI23a4r2sB6cqPqD1/f0NzWSf9HsUGz+KjdBusX0Anf7ZR82MBXHTDI
lzKEwX+2D/TdXMm9ZYyAQJfkHeVFVrmBe1Vzki50cUS8+v9AJgqTFKjkRJ9Tz4oesLxwCdVgdHvC
bWsZKK6o3i3isfcbqfKWXg5T6Qed+bZk+YxL6cluakBjYaRzr1s+YR5jP5mkxNQld7KG3a7XwDlM
iBgeSTWsoxjYezUZut9skuoOXChdrnYepCVzOG0evnWCCDCRGRcf+LleRjFUVHmTuN00tavlcIXN
UlQPqR3UpOZSWiQAd5tJlmNkCyvkc7BKxhs60iypNYy1dzZpH/tvOU6TRMd9GgRm4IdXrKx2Y31f
heLV8dO4KcYNeh0K/JI//lrJZijQ650I9odZ8JteLDJHuWEB97AAIF2p1hR8JqmuAWYDYQMZrbzW
XhFvplIEME8J6KrmYrjDskf0sUUQ0HAr1Sz/Gmj22KHeNWGWLJ8cEMWzcj0+buKVn+i7mBoF/yCR
mbi/xsaqTAs4iBnTyIluoNbpGUyezLeIgyLLJxs871nNNraOCOS3kVrb/1Vdy3PR+irxpl4nNdTc
TzPK95W4B+ALqIEzq8oOK/lAnOMATyxT/XSVleC9c5dJc6rxFrL/RusUjLl8yd7mUrS3BCW/65Cu
PaXR2mBLP7fKLnkPk6wqQltTZlpZDeqRUPyGvAUdgNMLNMe2MIJS1ObpnJEzfUpoQtDX+OhxYWuz
VDodmdVo/AGAXQUeb4ydjLlG3lh6s1iDdzPiOV6Zk5pKAu2WWScG7xbbT3bCxevMs42iZx20zF4t
xMUhXOL7gYdc/BpIuEvpu0mvE81n7ieVUGzbmJcZBeCzGr2YIq5kR4tSG2xEprBXsrMbyduQtCLu
2Jl8ZksfK+jwbEnvlktvaYJWedNkqrLUvcGw4eE7TTCYcFAq1hjL6wNKhsnP5kJS/x3Aj5kou2WP
ijVhBgHeDbWL+wPXsHIit4FC8LGuigoahnW8AYwSUdmxhuDKgnApjJRz0bPpcbvE5fQ66XENwEzg
8aqkMh7sI3oJT+z57lph9Lv/7Sxo4+8SXD0tuANYVHqc6ZEb9FOW8Qv1Q5hJMPQR2QW+v43ELddt
mQqdVx3Ca6XCo9LvBe3h+y9kOqgz2dooFnHIPAoDhfYjPF/MXfFLQgq/iOfwXif8xyFShe8QDGZt
DJYNkGL5toAlDVqe1k6jMivOZdu8hBimPsb+LWcabUtKcmDMT9OCNEc1haMbIxFgHR/72j0zABkG
C2Y21PdO/oVc8av8GPoeuaLULx5CsdiH9+MWvl/A+SghnLhhIeruuwXqknqgn0JqU9SOxW6QlktU
Kbwsobd8gTdB/LVAb6kdJJ5t8yhtLE9SqimHs/bNCIexOBs0dkCThTU56QcHAliZBmZPAst+5xhv
hWWTpZYnopyUgX1maP4IY6ahVnzSC6mgUY6pAcKOwKrZH5ulY6NISyWDowkz2Pb4TVFOEne2nRV5
vlIUvJsSEN+l3VNY/F2N4OHGml1zOPRNUqyxdpwB8CpJsGpyettBAAgXtL6+YUAtSKIx/4hl9PgH
+KNVKpNm/yohIJkVTgxiVCtNBwN5rHZTHG/2Jn66/VWmeKFzxUXTWobO0vfwWEd7+fiw7B0pn/I4
qvGhPWUBVJAlO+Qq8tSEjIHNMNf41k/55FG4sG4EpSHuuuS0zzNSIlD4bpeMHJmyKeAQYJ2ahWmz
s0IFx3tZI/1Cl1DvdAfiVuKR1U9LluiFEApioZ7hVQxiTXNoCSpgjKzDItm2XB2XyKq1bDbayZGt
rBfxtaHQOlig3+mWmkBtFn6fVETueYpnDTSVA1THnt7C96ipolc0zU/EqfUfTyhpVSglx56kfxjs
7pj13ahkuUZQQXxG6+6B56wsycuTzAALWoI7tKD7Tr56yBpFi2JUO73yJjOvmr2yCqiB/kiJGyC9
yBGErr1rYKCvPF0ehv+xPEofMIF16a9IK4ofUjewoptl7VsMXb6sHcfWNFF5XrQopoX+OydoZGDm
VWpDkFy0d/D5XbkL0hLoNH/t0nuh0dXLgacAocdxI8fE+f9MeXwuv1voGkQuHyE5lUmAvxrJ5fAd
odsFdJhJFe3jBleatjw76vgGRQFMrpZnrZBhpqpwQEihfMGEsR6WEY19zSiIr1sLQQFJJzCWN3/W
si3+uqTbXff3pC2nWKKb2cKkzI9JewhCacU7ht1xdoAnZd86TV3tH0ZoXQwDlKcvHidy2hIn1iCF
yXhkG72IfQ2SAGxfCHwhq4vepZPt+xr9W608H0y+9W02MuVQeefD+orxBTXg/iaOvbnVWgq3R9Jy
ET01PeaY1dxnnYdYj9km8H75EAPVyH+uyGCzhu3rPrKPVdw2IXBMQsLNAAE9ZVccJ2RTVJhYOnkV
bAEhXsTScI7S7e4PulTIjcik1aThrr2AdxAsuxEUs0wmXvg4Wru5C7wLR5uzmdTEMkEGCBxX1Hj6
oqdFoVGLprpkRDjRDYzTUja8S+cHTE6zMbc16wom8hp4Ii7fVhfEbDwEI+Ook48H84Ggvu2kCLJS
KaoARNUOKh6H7vEQ8cDWeWFBo68enLOb7fW5Hsvt6BW88AMZeQr0C2Q5BCycYUi+xqE6cLun/nW2
elu81ailIyE8mgnE5ycxiOwBnpAWZNaXkVVOOYXDq2dIPiFl1OEi6yRfTlbkji70EE3qnTFlPNe/
ADlZy21n1RwcLy5s19pb1TcyrnSaDW/oGYEJ9Hqufh+uCtUf3ixdfv8Qqqd0uIZ8eG2huYlC8gRb
kckPRQM/ZJ9tzuY5KpRxUoJA9WfEEKM8HPILzBT+4yTeBV4WrbPXAQPCe2AFVBNU0DCYmv9BVtmI
7cSRonrJ+jk6tdeX1Dj+80s3g0ltxgBJfWVPaLw9NyA8fAKVfulAO0G+4ftHX0gVgrZJxf0kY6B+
lsn/GA0sZR2ZVp3dnsYym90/9bnCe6W7ZNYUuZSsxVEo5OBU66g9FAFsm+6p3QXxwgKCZwP+n1Q4
I38JmHRor1ao+e0Z7oWGYOeTZm8aOqOwQ+MTcUAtXIz1HIUcFEDDOdlLUGKTIAeWUZ+SfhN7pBAp
mxq2DBRqV2IAzJ3zK9fDoX3u7BzbnWPdzTmKhDXg8uulM/Gr779lPnbEZ5t8zoKJzZXIAOVrGp1v
hd8TILFbB6fiHIRqg6o5AoUENBi/uc7lvoR4kF7P5ekYHuGxQx/OfLjFXgG7RqrYtx/lSn0pVHHa
gRzUlcsGmMv4e9H8VcGcSWCGd3a/t0/z41Uo6y/w3FRRaDo677wv3JjASfMSrSewOkKVUSvhJEeB
dz9uMnPAJEgJvLDdYxmSF9jIGtJxAnMQqVIKXsKrd7OLrx+7uNcZ1YQxlEsOgVPPNNQ7h23VuNK/
CEnO6vXM53J5OFZUrLW5bZYIWi2eeqJ9YdXahK7+Rp1vFWug519rJMe87NeIah2IPdQqXTfOquLS
ZRQSAMa/ZpqvEugw+vInQjQ1nqPCZj9aD6vdag2txjqPefNguL5JDpFG39m1Z6jUdhMbeDAG+m4P
BOO/Z4rLYjYzDDvU8y5LGt63aucnQwWm9qljJLvKXkfdXIiDwov8R3WmYNHUuhdp5KBuxMs+MkaW
prb/zrZ0DMsXaY9AgvyE/6lvDnMyzK8tdfcXfKVB7JGQuFtoLndQOnQW/2HL4+WlZpB5wAaSf02v
yBBrqw1rOJOi46QSInVWO7y/SQsmva1A7IRrQLvVVb+aaM71V7dLnTSCa28h7JKVgXjca6ixqqf6
/8xSoVmsJp3FjEQEHKk+KcRc7DcRdsdA4z6bjBqqHEF/2G1U7Yk725ZJwWMgRaQE96Eu9oWbBJCj
rIPOIpwTZROgrMx7Pi0c9ZRIaL8Zd5nkG/5Mn3HA0A/G/O4UK+OI84L17XH1jsj09PEHKemuz6LN
osnsta9jrYFRk7LudOWy9UFqbquSZJrf84UCee83rifq9HKhS3kdxo1xCMWmhCCWd+Q4AJNhYNDD
sfbw6QPRsKQcJGFPE5uQk0sOQgTbsQ1cHB3d8g6dhUpLhwnYob620SyDfryOmt7OSlLaDx68EbOr
GqJa0mDw/UDx99/7/Bd92N86geAETFUrZ+JUgmY40I2WJRmRfj2iTYZGeGiDmZMIa7JBv1/GaloA
u3ucI1q3S4KIEO6XQalopuhlr3rZRQyT5KvpsrJ9EdO6ubvf/WCtGtiFPHD2HyRcS8L0oI3eE4Cm
y+2gzxWOCR1a14GQA/H6C6d7rUbD1axtvGYuimMOijpPX7h7T7L2wJEavmTGHV1RFIDothX3ketm
9T9EMd356sGJxb9lfQYEQVDzEcqT3zJnEMQ4D4Iu729k1S7JP8c+7ixc0gyK1Yj+dwgThRAqrOYu
S1I93YwO9LcAmGpMlFvwm/ikCNqkwd5gQtn2lqn8PbNvK5blDCEh+ZUjiSkwi2ZxoKib+8DrZNGt
h61Gd1axGdLCJ73AoVkRNAl500jkr948tIXtCkKicADPqDTLByksfowuUQC5bJnTOEfCpYfJxFu+
h5W2JavYN+lo2nzKWzdMDwQGPSvBJVD/Xv+bL5/4iotBBT1zrd1YVnEXUDksN5GlzTAsf6gm7Arl
nGXUGldd1iMG/124hrIFB4qCF/lOtB5+MJaxLw3n4MKgINN1vBkZbufS/cwDI+gRYHGa2Pek6e9I
xJfOajDVT206EOBlafW13yoWIA4HSmCnBKZAGNXJSh9esN1BAfY2qwgbH71Nh3FTD/aGK/PA7/Bk
a1yeWbwdBWPX9Fh/f28j5y5bS6qS/8q6quXYByqg1cXU8NpC0PHpEc8j7qQrffCnGHgRDvb1LC0G
nl6LsdNYk0LSjSY2karqMYfCNuP+tyTN+MHima1KyLmYkrzv+Umw6l06jARgzncXDYXNV6cACsRX
Fl0RHDthEQljB1aFqNMZK+JvovyeZ6bTYuLWJ2JkUok8Ga7HRgzIqYLwwndBLckRkr4EK2fBKVgj
9LUp9lH0zumxTitU6hRTkk+dUZQ7cVWFhYVbL9Im7Ow9ozeLqCfabsbpODAV7G00cbfVtJSgThG6
JIXA0YlymgyaG7uLfNFAQoftoemsCl5O2ipJxerod75FEGAang6CX0/rCu4rgmlRj6J6WNvouRs1
/qKG7Pfc+eT7fBYvn19Ff0qx+A3Rfb4GjW6hCiPOGpvTznmvOM+0C3Qz/6tul5tyC2phqf6TYCJ5
aUzogSgpn5gmRE9VE8+PoPZkCHzaGWP2Kvc4eTMx8oUVyLhAzxW22rz2m9ufDiO7ff1kZrtcivas
nFNITlPPwmdUyXt6XqtZQ6IaqLtGdRsLpamXTtAkeTKmpFs8QJxttJpkfz+UfUkyUeyDyqGXfhBw
U/0ml13hChJQ3TJIcmqeH8fpAvXHBwLrHknRKiVfGYp13nNuFyarF5oZGtSjgUloZ+9ccOIxkme2
hEevvxsTLspPo3PSaFkajnX1tzx48hGHLF/g0Evxl2uwinr5JR7gNbgeArDrGn4FC2SBNDXH0IvC
nPJ9Zvfgid+wIePp6HYec7J6C9y2Z0bcGE4ATCeid3TQ0cEXkZcUXzlSHgOB5yVSSD01BEOswmBr
30u6vm9OHMvJL8XZXmfYUp6W6j34VqQ9UXGkzdiYjPLsHVwnzn0aCEuUnLvBBFZ0ezn70ykhv1XU
oEgNqDsRYfb/ZKQl+WTVCa/XrBdTp7bef9W86Ab1rsYMdtTks7drvgQGNItrQn1u8YrbD1ur1h6j
f4lfGuro6gfAgpTlRZw5zSdOMuayr1LF3jOp5MmhXW43qw9PWwRzuVMGkKTPc9RnWM6Yj9YjBUvC
VSrb8xaVb8Ez1YznkiFb19yfHeo/8muYwZjqnJWHEGnJcye3z9Y+6tYQuplnhLr3mBPqLwXwb1xx
2giPxTKzDegTbiMS/NAwuTzmhhxWjxQQCAZ/GQEsKVQfNAa3ak18qKb0a7hgiRpoJ+XoYxfp98qc
0rDyH6JJnKRqkdedF1ov08KHW9/DacdkROfXPBtWTN98UDAtxbqA2gp7BJUGB2ODFTvdr6E8BiXh
b3ddlqCx1jemR3+XmvxReP+1Pp0gLGApWbmDHBHPTTJVBJOvHk5XU65ChLXPs5et0DynHQjFaf65
RXNaCYoX8wa3I3/09n9rFX6V1q2tk23xvgcC2S1fSLdpy7ZGrx7bDXWhOOrRKp25Zpm8UGf2TYfC
gLotaC6WNyLO2ZddB+R3VCiw60P3hVDRak2QeRRXt8p0lT3drxnN2wteNqMh7ddIBsmU6mFV2OIB
7AU9Uvj6ie317zMdEeplsY3cgnjae/BKJQUda48AX/LQ0Ky3PKkJ8RIsnac/l6TJ4NsDDKAYav8k
c/Mr6Z/RkWbeVMf1CSdWpkuBW8SxRUlbOQ8tK3/E9pjSrxAAhWuks9zCc3Qwbn2LMW4OkNG/qwFK
pDzSHsmjfkqAEhp4FN8OmLlgx3xqvXGJyNRhXBnovbSQ75WLM0pQMIqvLy2LpJgT96Vq94cvQUsr
GmUb+0CeS6viOh/vmcdUEwEMnVVcAudHWsVpnQbsQZhYwYbF6gHAEGtPiEq0nSAVbRtahjwQTc2r
ANRSidT7r24EBCVTSb2NyFm9O8mjxXwdOSegW3W6Z7ATkJpWP+Nn55wj/q8M5frJh4k8q0Z0dYyZ
cbSnlz+J7fn/Szg1tMz5F/lWI1CroEDaoqEwWgCOal0hwHhbnVlDpnSX/Hh1ePpZPG5bBrCgcSSz
1aGthlmAv/fGQnyoOZVoPNRa3DgBUAr0C3Rn0UvSHP6Ul2jMPnA1vu7NH/uzh2E1dmGzdXbzKUKk
ulB8p/JqcUyjTrW8KyMaWfSMIIazPKFf7DENhuPOa7+LVHTIIdIXxyrdKYYl1wPn9X++wtuvR+9D
pM7aa1KRIDUGuA+YSRJFxL3/L8GyndXGvT81E7gOytr/A1AKAIe6YjqARoOQVO+/3NG1b9xHsWmL
eliO08W4L1tRvdN8PmQx1wXli0oTNlqWBB9KFE0HK9vebGiB/L4sEocb4z9m65weTn5Wcrvp+59T
NMsh1py3QLDWRf2uRsVm1b1C14NHFgFcgFjYrcnTN5YIfDYOdLPcAEXAXLtqAONenMKKvWQOHHoC
Z/Efv0n3RQ/dHKlurTfWB1U2z04DD5i4guOVWaTGHCyQXC6w6XSPwgxgb+dvlvc25Du5Lr3SXX+X
WxlrTumkQQUuHV104JN/f2T9mikZH4++KKLfCN3JP0NTQUquikIiAO3qkXsxNyErc5JJR5IB1B9F
oydbAbs6cLqlO5Pcdl1/YuulfNWGG20z1jX5/YzjbJOsa1f2XYw+wKvlGSO6nAInoEj7vD9AXr6z
UO3uO/EPfkAG7Q1Z2SVC/NvSrVA2/QomFpmi3LaNWiCntDokU0XMb7sgX/RZH1wCYhpNojuHZ+Tt
7eFlislxLGdY1wkupS2l5Rbyay0EN740veQDRUPGKlUuOCMOhxJgicTkgUoQPDDTKz8Qkq4mZdoW
nqLh1yCRmOzQl0qgtM84ggx9yLOuvQUd/v2WDpV+4/Q0x4uF4HExCdq8HeCr4M4pQV8PHjf7KWL7
fLzKS05ve4OKPNt8/e795hqJEKy8ICwS/EDVDaC12uRO0vt4V/xbNolLyTwu+nMmNeBwohIGaUhG
41UaIVA1uvRbZEdB8rSvuW3abA+8KIjDzbPXYbs2LxcuFyLuMqJAgQCq+MTEt5fUnQztz6zWGr/P
VxEPdIaGZ/hUKPyIqCkC4KJNLyuMRZ63nkfFVMAH74POQhuVDlsNKcK/pFPYljYBV+aHmyl5p4IU
dZII5yeMioQ+wCxLkTROyXagXxCjVgIg8cS3J4S7iHJiGPJZwtX/rxqRu1dRucBqmUFj92cDkMxi
vq57XiwI/AX1OGT2ce3JoPD+HOd56ycU8Xv1p3RUco8+w52cAwRLWxF4DqJVAhZgWwVge/tVhKu8
h3HVoiBP+B6mgjGZmydp198gfPiQcfjDs2utaDLov+b8GkdWLoD5Tt1u65Tpdt/7U1MWVOul8zWU
mTs1HD4xuUidCvOxRRkk6+7GnUfm8HKAooZKBLclwEb/dzJ+rkKOqNGqIs4C8HK//SaAFEHdC9Jp
E+J+Vr3/7V0o74U/sm2q41CsfVaqcJzYxc8biqEISg82IRGS60YM/mwJLfcqdW+3l3Wd+PBfThtE
yheKPmoQhRmsdlCRzRD5wnL+qO6c0TNScuFUfCb5a+z3VVQlIH5/5e71fCTutN2luBSiLS86NYIT
xqxdhhRuQHttidzmPGbwPdY20c25UK9JbUifJo3hzgbH2JqV/X5kNQgpUNCbkdfxcUtZ61uBnjyN
dBEDk66dALTfx6+Oy5MlFk7f3kvadYlcKdGYv2oC03Uin6egPBDuhWyqqCnk7ZjtqeXmoKX8dXYy
90GLR3Vp1bXh2PHpx6ak3MxDRB1dOOfZjaljIWKdVBi2da4LiuuErnc66nqQeISXjwN31huExKYP
ViPtIurg4kVmYzaELNI3hUnRugArKOoOOeQrHmVJh67CGguz0TdxzB0jfrDlZbK5uSNqnk2k4rlL
GLy9Z3vcYQC7Vuh4t8jxsCjKNW3cU9Nfw+SoTOsNfHddLkiSXgcbCQwQmduqbXclX0gCLbbm+8q1
WvJl1xPL+ORbBrhehwfhv6E1+2QKPjGIYhsX0PI6IKr5S6siv/Rxdlo0CVZ7SBHgOlCviQlrqTC2
k633uff9gJkzrUR78uK/SKyo6rXbEfOWKuTUUM+YHa2LdxofWb6idn15MSPmUfp9p9o/eI9QJA0r
vOj3EIwbReFvasech+g1QFfnWisblV5ClpcmnmiKp+bR1HOueBmG1TQ3ONo/IMqaKhE/l5B5LCxS
CHSqrSWphHu+nRsaXXJqc+aeh/ZdehQhY1q1sp1q0e1h1hK3mYxCEwj8xvHnD2i6mj1eJbqkZVUJ
XV08g3V+uXfv+kwMIJpjJRrPBMBHNuCOhTDjf49fbkERHLLXzD1oSCm5/kkqXY4F56P3xf+MXvMM
akhijln1P9qsCJVHSFaVrlHiyfyo+56sZkAdh1BlxCPz2g0tgTkf08KHXm0OJwMX5Grrz1AdRG3k
imyPH5aZt5mSQOokazhzyfJptcXOBBptw5ShM30sfkpIPnIPpLPuRzesF/FKzWHn2fexV3jVXgQD
sphdBALIXYy8WTTKIDOG/fSZDlwZyUabS/vzXmqDWuwZarhZ+zLYu514aTZNWsxH5ETnfXhL274a
Am0bmjT7dW8Qqpn6zy7DO+dv0Tl7UPrnuC/uzENNxRACHvzabd9lJG/5U+RETxOAiIe+mwWEWxZx
JHt4OJk9/h42M+5T+CiCpnZalPhIUtNx/4XGfKorN6CMRpSm+iRGs5wyMe8fm3wKT7sXoyHEq208
UL9AZmvPIL44l+lQB4gbGWfSbTpzflAW2WE3Z2j/r0FOGRxzUoFIAJnRv0ciKtUTQXbDn4sEi6pK
c2b0qDnk7g7sH/BY58cm7Nlp+4jSqbzUANWXOQpwqbfYF2xQV4x2kypzuFSTkzYxcu3Fy5BB1x3S
J6pp3u4715U4zUZZv6Ey06PvP0FfLoZujM+DhBzF7x8bgRk2izdytw7VEkNYeInYMbOoT0xcnu3R
/cdANLxhP8TAsE56zvHtVIUY/4dl9Y4AE8ZLgH8t7MERjpr7EGyKc27WmEIHexUR1FcTKsvaiK83
1F3+l4p2y/vkXB1VEZjXT7sA7cmR1QnfHutjpP+7+v3ckZyer8bpxTD1YokW/v++ez3Ra/mex22K
i/x7veRHCLPBmZIXWZZ3cACvup8QEnc208UaZoxth/laTOkvjSs3W2g7msXr/0HHOWBOMsFbD5sq
hcIkiuOJJ04xzgLd4X9AX/zAXXZEmivDHi+gXTzzppY0Wa1LQUNinIcXlVd627lvyuU62MbEwWAr
MAjwD7MOJcIKFsNbPCyV3Z0ieNGqZnEaqi5LlHJT8ca5tCtk9QedPeuOsFhBRYFFPG8ZZjul33Fw
5FzcWGpEho1Ppv6YeebRYCw4QG14x9/bUOQ/DJPACOv0bxOP/WpBUpppiIdbG2AFgpoEYEqNIfe/
+AMaV7asiG2qTy7ou51EsrqwbWqSAFE3b41h0TXkjnOejBISIXsWw3qKX7MDULWhbx0TZ6+sKC6J
t1esPqa7/hnDIXaNcOzcfqakYDv0qIdmtCz0yhRkwP3Dikf+iwQrIcUN4u6IaIVxUWATe1CAurXP
qTlWXPmpzpAUc6K3amdZafre82L7rwXXtW2c4MCbTv2X0dXY8QYTrBwmoOV5O5oi6WPfJb9SEdBj
4trGHQ7vdP+3FOZnVrlanl+mlmno7SZ9xwyWM4WI5qbggf6w2FR4l38dJPJtEyGXHRTKmJ7Pu9tz
5uFFMLRoMuaosZ8cuM/bLX2BppxyrIwqtUBGcrdDqNRQ/mv8w0rn1riDgtcK3+hNSa4EnLJILnsQ
nNVebdMUV5OaVbbpirukJqGpkmVlUZsGxm9VRBHxCW9XSGB3p6sYj+5f8jG533+gHIrbuNEnap34
ZBJIcQjaiWSMBthLtJFvwb83tywAjdvRiAjwp6CXW+xkZ0MFTFj2pHJBLr+eLgYNMZ4ftZuEY2OK
tDnfvBKuxxUR3QKQK6x5T32tAli1NPCjPcjmpe8GSRrG+RwIx9tLeiE1yp8z9c1MB7ug3yzQE5Mc
i+Rnr11xfdTHcPu9XUyz0rYSeVtjFp567YvC0lC9S3DakakiAR+NVqdZ3U//BaeNCAiLYiGEYssE
hEPj2AqwqcL/37qlz0R6r+OC4r8IzxKaJiiGkpmO7hXB8PVeva3IzF2NyEU+WAKrxdPbcMR1WRpy
IlQICSrRsd19Y1nz7G12RrveZUcUMhE+zUw8Bu0CM5MxXbh/x35KvGX2TJ3A/RyzKQ90SU+dGpIA
1Qj+xRfvcUL4Eh42Z85VrMDnc5MLrbIh39ekm092yiQgQ7MEFjxzX5IkldxPiZeYl2mpTP4Vh0wn
BSF88/bXNxy0nldaDaqy7ysyGf1deytLE9W4Uno4YOEOROM1fh4HKP93KtDqJfVvbl/O7ArKA1VO
H3IaiASE7LR3B+AJ+FHAXt8WhiVOpHg5QLNmqgx5l+Tvl/OZj27O/3SCW11jYgT8gUKw5UdBh35M
FVPr5+eEslcdqSALqE5Pd4JlUsGviU0ZF3eYTSy+ANBjjfmrprAYwJG86u6YSRh0qvMx9Wy+d/X5
/d36KO/LM//nOcriSC/r4QeM9hkElRdRk6cnysTN5DdUHXIb2S6IrrqoZ2rO7z7/+t3jQsxjHTBw
/7N8ZRRlg3CNBiTGw7JPj5RX2q/a5RB9jW+7YPG1rIQs1FzM1X8J6EuX54cCRb91cHzKy5uMVBUP
9E1zUZj15HaoxM6faWe+lgz6ALmoNUfso/B/A6ZdJZxp1TDcFyDm1UcCOQ8rJTaTbrNMoruNVue3
BVBESyX+32IbLThiaaxM54SbtgubP7v+bUsBuT+boYGWYF15oYow75USLW2szP27WcZIa/vvymqF
FjsqC4CBc74w/Oh8ZZYQb+b2gyPXrVAWt5fhtGSLDgO9vhTcNFf2gfN3t/WIP6RrtsHVu2CeCYIB
VEViRg605Jy82BQMh2suk8Kt6ZOpRcTiCrs6SbJnXGyDTY+UW4jWHDmMDXdn7ZhMjHUdoYQji4K+
JmbkvFYmIef7/1g1ZyyMIvyJrH0U30tCF1mHGLhg8VTikHXYu4CCon92zyB26AqM4Eq1GwCuTtWF
qDU9kU2dGvT72pYy5sW2vP1Ng928HgzLkRmN6U1w3YJLMUokEXzJTTpQRryZcpSrlxTbRC3om3AX
ltca8jkt1+HIVDKg2LvLFNwx0aatutgH28HfQcfF1gqiBkTyp9kdjxHQyoSv6a9SCSd7CffBFmMY
I6hh+bM0qo2OZTvD8x7Ld+D+s3EhJFDCXOdM5hd2n41/yyKJWlj33yC+Ve1gzuiuBV+l7GM3DCos
cUyUTMcktyWvB6XtGb0kiyaFPaR9uJpPZXLfmv0z7+KQNUWm5mlQ90CA7qZzR2Yk/EGFPceekNHK
yJoiobF3tcBFEipH5sn6EzU2uhq6ELxf4d0cWfwm/JcXBiFp9AhOBZ3NCpcNDSdNYzcZk66QiPIN
lYpbXr45nEQ8O+HzYOT581vf+vPeLLdNSZE8lQOCMsbHrKcq7L/3uuyfPZm8L+ADnvxQEGizx2jW
N5ni+pRJ3OWrDR5+lWooo0eyqzhPhBOve3A8Xzp5lPsFSdRuU+LDfGRWLzty7xVaoKGE6JQHpuYj
JjFc0n7g426cqKCpl1K0pVY4dWmC5UIgiDRonTkw8Eg9w9NP3OPyKf+Tzlv8FOt7AABVZEfwpSu6
yiUYq2+t2cAEzUNcluRelizuJEvPmIl+5ME+myFWL8buVbiq1eCalZ5dp1ZdnssZj+Tra1tvTIIA
YCGVkcR8dWmHvtcsvLRT4CozVN3gZCszbQ8mLngMEQRDAn23D9PHzuKut4BJXkDhSDIt8s+G4eg8
Dl2SD9YTQ1yRDQeSua4rexD5WHEVjuOJnYub90D5ndamR8mWCb3XcGJ/K5xhy5CGFtreqlZjdz8y
ubkMowiKvODptGl1vvVH9tQFREg9rk+TkuBO5PxWPc1tX6oYot1qS1UwatmH7ZoHiGqftbgWqmj+
iOp27Biko+cWG3qFG/ZwZaTTiNapMQZ64xt8Oz4hPnkONS6lnsOlHbzOB/wxsky+XFZKPSrX/i05
T0Rd+Wnw4SkJkWgPX/L083hpsIgi6ExcyXB+ue2Ady7lmaO1yB1KSk7r0nHAhtgaahsKWoLOA2A1
QoliEvQnEh/GHM1ZyXfUmq3yESSKtK6qBmU3QgxOYI28iUpLpUiYtSbBHQ/Hh/V5X0ZI/2Au4fW+
p8L/d+sugYMI9L+TUXcN/LaaYbvZmax/ITL29Reqx8maYLLI+7C9atcmbj+na7Z5fKPF1Yph88bJ
c5p5bnQ7M/y7b23V4TYc4J+kZ/zYg9r8l1pnnmwQKejJG1z12HBIwTDa7YLkuwIdsMYl1zHAgnCC
A8b5GEOQX98ZPUdM/qgFx0bW7h3bm/6vCr1FSDpobwQodESsVnSLKb0EqGFQfAhquoCW5qkIqymA
6UdqBOPWaFCWY83nrLYgNhVwE/doJpEpsQQw4wp53rNnPqqVJrjvFEGv4T0rnl7pKFe7UfgmJE26
Rg35dLWJUJcwLLbpgTbzuKo3WBhcpY3SnMUkMlkRXESiTYjftyftZKiqA5HVs9bXVvqTW56BIQQH
E/QHGHy+dTMz7iwD1jbQSTIYqZ3Q70OLloEzkAkuAfatBlAlpU9TlQyg/UFSQurz8QaWEv+mxp4j
LSdRNdITunAiQ9u07R6hFghfiD9oQYWpb1J7N9ya1u2NWWsUjAEVKoskcopIgrU3tE/iEA3SoE5+
pTGMQTGDj2sX8i9DyRPjfP8p7R4LkjVhi/mNFf6np3HZ9LP+GWvXe7q5r4A8KVWcRh6W0ILlW8sN
IS14lhXhAHve0tH2cL+jbt2Xo9Y9PMUfle9rjUarPn40QMOh+ngvQ58EGUWUi3mcwSw2Z+tFA8Yd
v8Zhe8bLplhJ116PE1lNIb+Yin35aK6uY2Zu5jZmG1EK79v5HytfZB+LNKcxh/THHWcYJOgNbrjw
/zSU3YGhxGqfCuwn0f8TVf1JPSdQCt6OWvew1bsIS87WQL1iWRQyknagBPa0h1GokXU98oWIqrVp
/tVa+wxgfLpaTq8ktV7mqfTchbLEaCpcUzgZk3aelLioNeWWYFpiOvYPcStgPCLWbWi3jZDiCQ/M
l0lijNUWb7SNeF5OFlEh24f+TZyO02HzfBvYw9hL+eiaVeasQ6U+/KUN9cRqV+kEcT2zzZ7Hdq9f
ziEpY70pxOodEznHZDXE1BHGRiTbb00CZzhVgptrsqJa1AM0JIS8x2OLaOz69VfopWx/sMBX085y
k6RuBKTzdO7MrxdEKEOb+C88LVVMha6/OscuwEvEORBLpcSFDwSUmYjWZp71BjbApIUz+lJSFjjQ
uYqueGlbbPvsTg6n5sUphsevbtQGQBxXzO6K9GioC8sNONH7UVt6xuR7Xj0fRnJWMqMIlUKmLd+V
XeUGMQ5WUDEq18zh17n+hL09j6JT6Fz0VmOZGYOwZuoRIqeX3vIWgiPlyyNzRB3DcJFE9zfA+85H
AuXIOTfBxk+E7tOInSMlwXoEaJPGS2tEnTsom/3FrMIv8VSY+vxuTGrsOrNh1g8kaKLaHhVTpEnW
axDSlFX/e5Mv4/oS6FJs06si8izOdPhl3YY1n7pugeJb4PoUhThkcKJtNZ9uL093A3FpVZ1UL67D
3Nxf1+phi43kGL4KBnGhKd1v6+3WFopHW1fhSMRcttPZMjvsbcnWtHJO54I8q5QwvHBPfZXc1Fl+
qL5/1nh2KVv0ZvHrsTk1RQ2bLMh4AfGGuho9D5mJJgbjSFSxruAGpw4e2lXyaUtTaOudZNarEQqo
gIy7vNxIWVtzi/BKv90RF9RCR2Oq+UjT4UnOxTiupZWRnriX4xqUbGQMm1U0kKS9q2YXuQ/WvlMf
jXOgvGRqPNTUHXfceJuNFlGHoarAUvTxflSc9vpM06nP95xrT6QkgMjxBHr/C9MJ04GErtEG4sCM
VGSCiILaZL84Z5oT58Bk3wNZeu3cRQzs2DryXHXiZ6o0u50Rve8TLdQ3RAUoOL+dgxmg8SEk7Kwu
rm02j7zrYSVkdgaBeS+as9JKGNR9XXbPFkIcVfDsE+Q9G4ZJ/+7WXqfCXtijqHg3x6VIZ/alN1mf
4W9b12O2ZTPITY+jof9pAxNwwiwfKhA3G6Dmf/DYB7vjkhGfpeVvw+wFB+hUpEyijx+nz+6KgCT1
/Vth+xyjANfck9vndAcns2XrCFkWbg/9w067Nn/6ZDD5fk9fz55C8LA4pKOLk8DUohp/5B7et8Qq
z30xw1duagRioyY4h5WhbgQdXJArQpg8QwrL0NLoC5+DB5tNTQxCpkknzGYrezRwOSp6IvANonsP
Aa8n+BeoRO/VtDfkNXCe7xh06re5dvNrtGUeKX+Mfi6zeCM5GktepDhwpbyO8laZHA7Mhkr+61yy
+P28A+jZkQhpT/vvdIyKXqinKdGWdtLZxd4CbtpGE95L8kEk/CDgLpeicqkKOdpIqLsNdTkqQqQH
WbqH3y7cD4RW576HTukwRguvC44jo0najXXGHYLGQdg58i1BTffVgSl7L+XSRhcx3o8FPPNj4x/n
yvC/87MaEe1f5ZUbEme8gjA1RxjkrnEUgXcEBgXFaDhTO8q3L4Snu6bdenw6VPJwdbzDx60uojH5
q7zN81AqN9fE83P3Ym3apXez9O23KqDASSTM0cYJqYYLIp3qXMULyG6DKsd8PtcNdV/llzPJOm23
oDLOknmxl42uMnNSkZLl2MS6Qd1u9A2OCoMFmnm1TVXTADhKk/i/DR/r+ZDAVje5VhFecKodWTIb
45/i+EgTVoAZBgt+/CAnP0ngL5r8hTLBD0QsJmYsrBsNTd9kteXGL5timB9JATMDyxYAoHnkSojK
ZGym35aNf3LF24/zYT4oNPPO+fi2PUvOf6wn9TMMWH8zgCznoGcP0PMroZG3uSwaRVa5YyADEtp6
3+fnaHrhNDbKk6sXheKjIIZ7qV8yPygx8ZJbHPS1GaOkziSu+OhafgCIVEO8qdGHrLxZk/UB0562
r2ITggyRLjMHlcKTGTcoZD9CA/UdeuNvVAwG/VTBC1MnuWa9sXBiIpCGZc2TqPSe+86MkcStaM1x
Oa0y7sDdzQzTmDT/44n4LiM4AOK3EMLqtA73n+NT2X+tKi0tBrtN9nk499NUjNafj3aZbiEOCxCF
cdolQq9KJqLb3LkPeGRqF1M9ef+BR3rZS9mKMpgwEaPgHuMU5rPvI4l/PfhmkLS+22BER+lFGlhG
a50V9/2vH7pnesXGsY7c9KyyXfO1rdcBTY8mQkmwqEre/ST40z6Mqi8EhwAGq5AlWHLTUgcSxbcm
F4JXYbvEREV9U0GCKjkj5ikpxd/eN/wkvnF/Ig1483oZlpzNB+8BkuzpxUIj1KASur62l/19Nhcz
NOxcmZjoFEoxWLGmBbj0vLwR/6ZKyeeqEL2eC4ZaPikYkmviX64I1IuczDpMEK+bXeMJQT6Y0ahS
yxG1Qcw2xC42lFBPDLBialrCoiWEvCHpJs9FoYpz4X+W2IwG1k2TBymBHrfIwgp3lBoGIojhAoTR
c9J4vvxm6fSOBtVgms3Aicu7YQgCdtSd5+KsopMVTezEIvHAWVv+4puZKLeEmnnM89bBt/A0AnLg
V9csoNC5fLhn8yR6ARgfVaKcrqRWruorqpKXS5EOLQe7mum/2YHRvndx4N8yEXYq3Jq9bslUT9rr
CUSOFXQ+cIIUXL5NVUIdSBmeThxebrdo9lJ7dJZ1TH26XaBagWL4MmN4Ll3WNZME4lV7mfIKHW0n
mInP3xxTlGxY99INwSynY3NpH/WvSdP8dfruLJ6ibMvOyH8NQsH7WpM1PgyVersAOoWGjQv9LZdJ
2+0Pq7kg38zgGbgOhGfO7SQzfEGVN769GzXM7RqEZMCw9qy0jNS8NHIqA/JUiKMYbaGj4jFjt4Wo
XW6dMHSmBJDMOrdmoudm3oX9064vVHqEUp9kb0Q3YzJTGnoAGDdK8EjT3alKxynro+ZroRYU7FW9
YV901/e7tahFEvn/0VR3b0VOndaX4ghf/BAaUYSsULt35KC6SfQd1fFt0h+bSf3WG64VTLTTBSOt
7SVwfd/OEQwgwq5UdD7eoMtUOh+abv3ZGVOrSmyYCg3e5vge7dM1xna9Lvt0iI9pfMrqTxWTCqqR
Iv2pijB/2evg1cl6VxBpBmxdoUdvm8cxUUcsgOPAJ0xe+qZ7I/kfjfdKd71IZKhxIP64e8gHKLGS
X9BiIMd7+9FKVrtXVD5yn9+63zkpSFzhqCB8tQfOMZ9MH0PVtlzfC40GEAzOzwttj160DVnYbhbf
Qq6wZqVOTqWgifEtHIrTYwREGh7cmvlWfxUvYPCMw5JVJFHNBg/FY27DhT8kutVE6KTVcoxXPRVn
sZJpHLE9uOSJlBXOwgJ/ryZOOZreLoqBFj54CX0Lru0ysZ0OR+fIRZ85H54d+epKLnZiNXNohGpb
gkN11H0eX/PbQUMf4ZjJqmUpSEmu7pZ7tvn6IEF3U4hiyKrz60SDpE3E8eWeT++IB6VGJwF69arq
artGLoILoHgSSgdmi/9B0xgH4T/imN4RX8pXlx15C34uvwl9U/NvEsG4UMvilnYdPSkycpfKQiiq
b6itZO+vxKdIuBdkQjTqMIgMoxTRXDtHGRgnD+p3cjrfP/SloU3UvNCC2/eKTgz/yXCu1tdKIM6e
XJOgvBxe83f1Q5zVciS4upxBwE/g6db3kiEB6HHZCUR1TVYU2jMitOVuD6/7c8/OkcqjCSqBSLXQ
4BAZOo65+KLJHrVJ6lI1Wq8N0Zg8FZATNUJBesWqHqiCtf7MoBfh764FBb3fMOA1mcY9CdPMley0
7m4IM44jbG0dMcitpOPW6enJAF5ijyCYwWWga272msjb+6P6wV06lXDpq/4JLexQP5ipigcEjO4b
svp/tD+7cbfPcNYr9jSVZE6vNdrcwgvG1HrdCrxgrt2MotG1ILcHIr2ofYggBjTEXbSyBTop+OuN
1dTHFgqEMDRMJD3y1RVSorGpoyiJkDWA3J4DrFAmPBPr02bWPKLXzfp4KTcu6VKq3Pmyqbg/c/87
918KJktozuTGMjDZHUsxRFpus7WfQvED3zyKx9CqI5zxt88QgGI+LUwN2Q2JyoX3VYeV7qgsQlW2
CE62nKjt/Ng4yMs55WFPoI/MEpJ4fBil/zrBYvlxeNgB2Z/SLfBLfZkT5Jq5sg4eX/gXv/l7SMqc
Ix/TjCsryHFALzawQe0g+fVfVB5Y5Pacz1WirnGz6Aq4qMlObF0vkNWi1TdgwrK9psU5A529vFaR
peh2ve34aohiYFeGquo9wWTXCehfaeNUBpzEarwd6OOMyDUeBwUOPpw/SuzBzPw2SuY77gAS02Me
SWarZM5FMgUkwQE34JTVdu6LMyqo34OdPluiO+JmiKAcojKAkbymEKTfX8WIP/0hNcr1YOhSFkA0
0IdbSmfO/9uUUjkc29RaGbo/9Wds7PVnAw3vR9SBiIBAWOvb0bJqFuOSbgVJRUFj65C9X8cTel+F
ZTqPCStujwD5Nf8Twkw9Bti/PdShktuYPBHA2ej3sKkupthSzZybyGJmzyZuCeMERYtGJJiPeEFe
Xpd0e9xwAd9kt+/5sjrhJAJCHCgD9nfLIBbJZpB9T9H707gMLxD8TuJeWOAX1A3a7HCYR+esFfKm
q4YILlHotXZHu7Ix6vhQmtBdLyBHkZo/JzCjbx0bAItW38swbn2Ts3eeNX4aw5QJKOjaYS00osxk
NhXfq+XqCXAhm622bZjQ91aMqhFEaJZvvSnkKrYG71xhubn3jtoScKqylnasZ8w8dY4X4Hth2y/8
GrEYjcGeMq2fg2daK68UhYHbtsiCM3+PlishVH19FaF3o0MneFj5iQ3lYEkYIcwOXnKGq8x9smW0
rfhXOucPDf/BIQoHg2C4DEisIoVVbrmHGoLyxekvXBDVtkzWZX6XXp4KrnQFwG9QzqiFtYajz5ll
Pd5hDKhI3jopCitWx2W5JrKnocSP7uOrPOIhEhN3uyGlw6jB26XOabduVEL/E1kbJ2n3ObfZ3A+w
9axpa6C9Q1nH54cLvxCQhNYmQBxlUL9e8IRPDxdVb1R/NAZn0qLr8uPKbpASi4ZxaJEfFLXqZHUw
HKA9I8OJGM8VOGDguxho7CSTsX64+cBpHsu1NmQyIu7cVW1SVGE0AT0saxGG8Rb3sUsAb4sehyVA
jRQiMUm9+E5kKffSCLR+Upwp9RoNfRxkPM4OeKWeCC0X5mXhyEJtESHf+FbnwqC0W5s6k5v5Puej
hs9QIwzfJxghM7/mlPjqIsZ5Tep3+cq111e95viDpU9FJb5NTME3JJvu86zRRvq3AELdi1OPIjyy
+48m0ulfc6YCA+rlBQuZYCMVUvXV1bTwdN3NEPkFeZLdHr40yfmSm1FQxtlGnC6zjQULhtzbBey1
v3mSs7mBGAR1Ut4SPne7X4Sm1cfw/0W7uYR+XygW7b/2/L2WV+8zquSXIdb0OY+MKPIKwF6P6BKk
kIbYfBSgQF99PslhNDoD3Uo5u6Q+fQnt6WsNW/f+ntRdAa1EfFQeNGwW71lCJr3H/Y7y3sQUZ/sf
2ccBaqkvOFIVpzj83aMoMp35urAKf0FHOyePqLefuPPSbYfReW3xuyDA8BrWqQ0jpE8MkPUSeoTL
llIKGyMxO2fsfIHHY+bkusFQJfx7qBZo8EOKX+MK4NWo/+B8axu9N9PZQP3uJIh/iT6eIwCwlrK5
R4KiqXuCS/ry5geaC9nFcQcntrRMQ7ImQkLk3BUA309EdHKtOaG23sU802FwwbffrVhV3Shq8xKj
fsIuEoCb9yf0+FDYqUWg/Em54RfksEFfkP/D7aJAQpFDanCGE0nwWHeCSlKt0u49o6N94xO8cITP
vkPkpXteE4HjHiSk/GcryrYk2AiAuKQlzHsuxROX01hxJ7R/Zw/23YKoAWKgAlLDXQNYoez+M6D3
s0qPQvVyLvQYMCQvR6mwUXZJ6nblwykjjX9TUwe+lxPzDwmfPb/DVLMAjhPVXzxUSpnOZB0l/fSE
iiuLNj+aw357nEd8PcOBXdOwKYW5KkQR16bm+Jvy2iuvAG8520qfHpZPWviKm1Oxryr41LgTFzVI
YsLTfb51uZdypyfQT2r2uC8UhRBA6dQUD3mfr6TGkkUWrYevfig6YZ1aevSZ52O3jcmcXU1yfLtM
K8Erch+Boxn1W1Z/eh711Wdc9/PfVEceCGtm+a9RqNn2P/LBMd5Hbxo7kHmof4EwKkhx26HjdCY0
QPHzMajj/ARXZimoBEVZ/UOSFvgniz6Rr6LAEQzlTcK9nJtGzzTDMO8TLKeiM+pLpC4niEg8kABG
V2SeVFsLnuSJN7xTNUpMM/Vmohqe2dJgm+JwQ/dPfpFeVwjeY+ogs56cGnz/s0VZXfAicoYc4XR5
FJC6NA3CGW1fXgCFXcynxf6xWscWv95z6+NTaJnw/hqIDcNPSnBl8ZFXnjLaSzmsn39f2eTBY+PX
fd5nwQmdEh8ZYPYXAYB0XOuYq0bmbRzKQkFShtFwe2ymfno1TysnMAqPp/yEveVCa5/qgrU9OJZl
0mQfjt9db5Z7u+hVrGZABofQGker1wje2lS6ZojUx29/7UkA2d98fY/3G+vm4IgSewuYo0ffUbsn
dONhNU3QmS7BsheQ51iurm4+LCNms8aLI1XCLDpgAyNxWgELh+gNtXRSdvicK+oAjQA8dlsV5ppf
WCR4vvdbEqJCDy8HFeU/nsanBzltOPWRamxbd8GKKcWOIrg0q7k2kpW+4j6CvUU36/D+0PAxdBWP
nGTJl0ugnm2cwyeGO2YfuGJaDtZj3GRmQhwwpMIgPcDz5tb7LQUDGNaCaErppVp8RXTG3z1ye9UN
MVfjZhFtyBs4wVd4u7LI3o0q9pJJARfYLLN9dCO8w1Zd30xrywHor6S15+utX4h/6N8GKIXo8SNK
ufJHX+8Ld5BSn3ow6U4EEDu3yv9Crtw++Sc0JyRrrNUfnrmZly/DQ1Q3DyYIOW9z+/PScYXNxhUF
j+T4uDkU/YVAh+TRp1c9kTCXtncw7Rqc9cVPY92L3lyQCEN79zlD363LEF1m5K8VEidMRv9HxLam
AwUmNqBQVuMS9deWtXZ5orEQKovrOhxYfXyB33ZKEjHCdh8J4PQ/E7cSdSmiO1V09x2ZshNt9Nfo
mzxmKHXvuoQjxfogTlRjM90pbATR5v1+M6yXt+2CXnLLOTWBoqQQ95ZZkXmplFI06ylU1QNKUx9F
54mkBV227DPiN0+LPPAmOAY5UGueaB/CZAXNW9yO3WQObequfjubvTs8gzw5qPuwjmjW5OMoIwdd
/Eh0xM2UR7Zo4WREbYOVmvDdwvPKUl7zxw/CkSY3bxkOE7tRQ89nsjcNzKKv1TS+xY7MkNif23++
+izG5ylCZsg0/1Eq3DqRaeiUYqE+Ue9JrC0Z9VF3ddqdK6321nrCHPiFrfLdAKeLgsKw+YupxbWr
T75dYo2T2HblzcVn97fOx32ob0skasZsfBq9wH8iI86DkwEBWW09T+2vXbNyOQ7jgoRpE3DcXsSS
hylp2YzLbJ4teVY0zBPLAyicbYbB21CzRF4Y8hmS3bbZUUjHSAkBIYRRx4zxVr/6Btrz7F/hoNZU
NQ5Xi64E1CTzwvR2/vPk1s6rPPmEGfMPnw8fJcgayyiX6VhuGBkosM9pXbziBA7XgG07eAVoLPnH
CRrk3hqPbjIEw4HZaTK5EhLVX8EghX2vyGyXLGtGVQ5V98qz1zz9nA0QyDe8MI35rPEtMA4I4j4K
6m7NG/NoCO9XGSmXBVeNU1u3YDVYI6u6Dsocvt1YVtO8qTuNS4lxJEirsphhpNqV1OXvVlCifXxg
W3DYQ/MMkNqgf0LTPoMDPKWqD1VkPN5uBIK1bCm5Dq/HPFMqR4o59UUlI9D3YoGJgHxXXkxlD5sw
WbhOvLuLZddS63fzUyxVGp4asD+ubsqvJY4XM1V6+KfnmFmwQd/JksdsyU5fQSCcJnxZksrMBJDh
a4Te+rT7SI9vj8jlAOj6UQq6KODk31oyE5rlFd4k3uF0UofW+oFNI05qrQiaHuP/bwI2sZhBju23
dyrDI0weVWL8oGWiSZLYfyz5LTHxhBFL5LWRjsG2A+YEKaB5CO7ymBR6d2NqMZhS8EHkyhTY8HDb
xVT30jm4bUK9nhvDABA3P2GKYLwc4IeY5ErNCNRbTto2BhWuHsCf+UT8ORz7BbgiezUxU5LwkI30
9vYTvoVxoEq2WNVJRuwKObBXZMNfL5/I6O+9sjrsTTpCmRG9olF2hAJQAABgTpUzNXyS9OYpne2K
YqLlLRYpWkMoKekCmhPi4xz3p5f9LY6qZSIFSUaNh9aYS2LwvoRECjRIx1yzIqAHSvlhZUrmY8Oy
0Pwe52ilGfqPd6vxnxUVljKDyH4ExMEFhS4WrJg2Mj7wNwPF/0VCopRM0gOWhLf36yiioZMmhsv2
B/FrsqIioKRfHcebT9ouazeW7YyDP9TIOxFPGyGfiH5rEfuXXXm7kC0PqYQ+x2oDf5VKflWS21IN
7m5M5NnVXDn25Zl556SXME62hT0gci5zVytwE+o07M0G/qEUjKctb6Kqb4IfuNi9JYpndNOkumxo
/3rRG6oZAiIXFOzNToGxr8ShoEBtuYkXMWEAGHKlrYcJV0sKeKOYvn7hgAeygZQx9OGitxARXZps
zQW5pyzkE+yrnjnZOPN17g3EQXsMBO36YWCVcE3u0q59QLZbYPuapl5lqi7TP+z8g4rG8mhGA52x
VOtvr2dNIjxQ1ygQd0vRF+TXPVikQ8BFiIzvC5MlDxjyU7riIDwLN9lefa6MhBk9oM8z55SLh9d/
TX2FSr4zCxQ/BHFagdqV45OLKSIC3yvgF9d3hOgYOi/b2yLr6MnmaXcd+MdNxIRu7t7wdFSrK4NL
IQSqWGei8p5G3X93RjmEq3PbowxwBkuo/jKrBmvFkd2mtDz5UOqaurbhRC/T4jn4GRAQ7V0kH933
FmeNqAL2UsCDOFOYr5Bwy25JJyLYKizkp0OG8ugt8VUX8MpGDsDzarrIbABM147W4zAGqeSFjHGE
uo3Xwa5AEHo3msERJiRH7NdgHeXjfD2KOOEuNgq8nqIOdwkFpfgJKNLVVmyVg7GHY6DW0BOHlPA0
CzwlA75daC3Vd05WGVPHdJdUH2O0zX5BgdCCrvBB5K+p0N76lrZ+58QUe4hXsh1CbV90Fz4k2cYY
+jbqXvygAJ1E4mb3xYt94RyNB7GsCTSJFvyDKEBDb/Wrdb1wNzCzDtqWbEN8KpKBiYPQKivHBBcr
EYnW55hEn1V6wh9iJ09zKz4pre9NEeZwqbTNMUQPNysm9JtygGptFDzpXUPjrXUuGq6jg8UU2vZt
HErKxPxUooc1q9SSnIBi0BnYGk7LkFau/vGYfIXXqaxOwllMZqlK93xp7osj1PTc7nMTpouwHfIY
vnZ/2wPr0zcuR1/Wah4Evu28v1G/GjsQFtPDKz0DROtHIcqhj0KPuOB/Nxlb0on0z1b4MEXl6N2a
s48BbsMl/ZaisoEnXAx5kshpssEnxVGPMkUyGjmdwwcsmujPdJEq+KhqjdlLuC/KrjM561Awv/uy
XTpBZZSx2F04bALDPgiWgp/DFA2XnxURQwX/0mBpDlunKYu1VpwYJrdQyGBVaZCg8K31Idr2NCKJ
73STolzBR94Q5TV8TD+cTNrgrwHjvEL5N73a0E2T0fYUNP5FKuYvzj7lj8n1gyNWESFJKgu9jtAw
sIFCo/Z/y1Vz8XSZeLclWQlpCyUn50vZvIUDMeViSdBvLNmp4NhFhcks/sgJdl1cm5C+1j64+rBq
VAeGdrx8aDqSltqATFAdbrnf0+i586PBNi26P2eInGqnWeiD9mqGL+2Rbpu2s9ptdcjF1NyJA6Q3
jSZRwW7L+5EDB1Dx1vqsys2h8upk0F2GHlH0Y/BpqnRQ28Yv2KzqxIs8MNBBN4MPbFXwNS794zeD
UI0M7DKZQSVR4X+x2s313G9BicIY3HNyV3krMjZnUCzCA1M5Giq7lquY7hzuGM4KCOECW5VWe0wj
19hvHJtIyFqpY9db8giKIX8LH0e2zBitsNCYdqZSNahCZvb40jlzgk2zzXey1jaIF8UX7SoHYvP2
RHuo38kqLyKjh8RN2MB5QrYb6uWfi1bZlDRn0aEM6Jskq43Y5VbFLgEMy5fxd+W/m+5ForY944gf
j1eRce6kAdXVYt865n9RpkuU24MGddzkDfgRNj/CPKVrftFIwZH6S1jRIMxs0b3fpCXGXHC8yEQc
XNSxH5n/nSf74n90KkSymA2tEG28ZY9niDU/D0TiHLyPBTwa8GmG0cOxCICMaRZ6c5HIMUoQot6t
qEMOz6+wK2zq9gWzPMvvCkEjuDSGp5XNA35sP64/lRByG+CmI8TRjtJnPe/EApz72lC9dfb5DmwZ
jTtePrX+zYjjjMdEx+QRQp1l60+COvgLmJE0G+ZP+BkPORLaMoT5/M+fDyCctYEdnebqJIgO4xQa
Ev0iy9av0hDVWh6NGigTHti2UKrTWXxBWVoKauf7OATl0cfPj6di5wDP0RR1qrYFIN9uIvIySIig
hG9Zi4XiRpJGdRVdcId2wCX6NZoj9MGO+5DpdhP7VInZ9eDcuZueolmMJbSvz/JBAmoM6OtpnHKT
/A90nVOTR3Enb40ztUgkRDAcuAQ0J43zjP2qTtjReSt3629ISVP7dVhikukfqJ1o5NfDD1a/7BED
IGrqma8fiJsZdS9zci8E1KYzq0RFGwzsFcsqRDZ/4mwkkVUd3RKzkyEypdO8c0sG59BsGGOEIEej
6sRd9H8xNtlLdN9FsnqNpZeRnSiIRKuE2agmAOgSxRSRHE3O8gbrbgSzvr4iUNGbp903xFT68mKL
dZEoNZQ3BVYTEP8hielJ1q7WIPRA71Ui+AMFzmI2OyenXw92CXVdZ+qEgSwIcuchBYdlRUa0+f0w
yAAlHpKVf4rPYu12C0x8ITKQ7sdDxyghlC71SqfS9j52hcsyJIGe2IKwnC3vBILHfy69FJcZwm4E
kkcx9VlsQN/cRjOUAAu8j+bzrMkFm1W1N97+geYDT4UYnaJswkJsLIiRi+y2qGJsSWkXPgCqqDe+
8dLBGE0mUkHcJ0OrpppXVaHprddZEBeLbgkRVb79RbQFs4bS+sSCxDOi7IuMC5uXIy8n4jL92OXA
guQAcowuqJLmKaAL8tFEOfwePTBErFOXr14CxP+xL9qa1NkrCsX1lxzBIiflODp+V3B3A0NtwQ0F
XndYboIH7TufpR11uMhYeeDKYEDOBtvwHb7hDs6/D3vt0c4+dt0wd38JvC4bM6AZ++gORriWPfoY
qxmhdKaNU6RoAUFz4ipNb6zi4StP1lQMuDk+YJx1GSbmcrvdvYSmrmh/SQsgFI/9L3VxERqU0hbY
6U4FGUQyULKx1yu39iH8w3cBTMuFJO4VxQ0BS1T6+nj8QL5MuV4i2O0E4oZGv6P3eL1MU6kyixuk
VuyNlNgN2oC9rjx2Ae8QlIrSKgKVrKZQfPcndM0N3hJTkzEkqLaALWpz3kB8PHHoY7+d7FCnASGb
/QPvhP4YTZig4gq0dmlY9o2sVrYPSUVh53unhn9rIZcJgYbDlFO/+OiVMnU/tSj0w+38VXST0COv
V/ctscVcbM/sx5oV9/Kv8FkJ4nByidxaeKuv1z0Z2KjnlshtdHQ6uDqOrdxLW0RZL2hki+34svIF
ehnk1hzRbPdOwknOv7VbvT5KNmP4N699q16+EsKLOwQK1KUWjSW3IvMvySFcCfKy5Yv8WEfxX6NH
HXUZ3hvwmWudBNtxOouLfvyNWiM5bm09u7n1TVwOnZdN1wuMQ/uRws5L+wdPyAEH3DLiILtRukC6
sDCNgt7gSi5lWzk205n6w/mDR8m5juDJZQWXfVl9iTlGzaxpyCbFaKZuxnNFQdVESzuQmF+MUMIt
rXH/SABF6/MuXWwjFRdvjGrMMRyvsTZKleFOqRug/gHL27Gw9k0NROFoasGZmEFrgrZcaRXk4KEa
GUm2CLtTzBD3j9/mCKQBF+5fHeKyvuZRfySDCTFQQWt++iUCT54K1LuQHan9EDHQTuDnHCdOIu/+
yFj3A3btCsbxTY5ZND35AoWX6eVvTsCZ8r353hW18g147O1ux4C5fTKw+7ptuQQDfXGA4bH+f6QV
604ZUuPfq3UE9YSe2jFUM7U8yqCYXIT+G84Ad6g5t5kW9fqHYl/XWnGYLvx7X0tOttCfBxYFo7np
pS1nCsCTXdVkTTZbkF++V2NzxqnCkzoxLEFjX5o/uopHnsrIKx7wKc1IVstOr2QGv6tOmIO7N/nH
6xUUfKZGhgrpt1FGDsVhA/rvJ+WKDGmf9Pkv5KdpA1y2mjMkghnL5caye5vlewmNvzFecdqi1O02
Mk/MMTSRdG14mG81NuZNcmgLao9O9KqLQsENoSIRTghqM/aoFyQPNwSwewJpXDaze218FSjfGE4Z
KbeCUOOCtvLz2hIQKozXRUlaBVbkQMuIBN2bbD98DS85G1rTZQuMltOJJjAuKcEwI0eVJT9ED/6d
A/yjEP4qYxfQwyM+VHr0XqzmsKta211JnYjkkKYitcVe7B6QD7x7/wDWHU1tDpAulWlk0vIHf3pF
8u247IBCXT9jKhxruMPmQ1yJ4uvkWTpQvP0HtqvD3yaRFbSQYFqOtOqu7wZK5B2HPNzKeVNZn0xh
PlpK1oW74Pa/u6hNzzkeV1zpwKu/eHDFd6dWYyJU6WvZ+E56TCf3qzVBZbSqIFJHQpY0MU3AzeiY
Tq6UPyldX2KO/o90sXblHWSN4p8a2mv3yHcrYpt1pJkDMdnk30FwP7KvPa4UksS6lGrQBkdoifvL
NDA9fIfqaRlhuYDpWyuypI4YGUIGWuDH9rEGFTFX/adYZR7ILFKbRYQFbcv3bj+sNyogsyUIhxAL
AILa7dpF9KeguRbi4L2x3gnF/YAUy7xRr2aooE9irGXc3OrA2pV91bOhk/srivdKsxeSR61pNUH1
CBjg2RnvikhuH9ahbdsopyApnSDIKuiz6SH+6c1N+LrhhBH6y1k4/H0mk+mTzMz6kSpZolhe3Uhj
ofrj6ULPQcSvRW9Aq5LnCtmig7AXIByhypXyBxA5aCJ95g2IofNldtSc++99K8CCe6ROjs70lCBA
eB0cOpMI82gdHX8JHB6t64sTuEIIjs549gDJ639TkWYXKLvVuOrzGyanX3efuZnwtS2dMX+Xg5J9
Dk2oSgRAluVTupPO8ta8KIsHgD2tG5zDhyDKH8oAskktz8AORlKioCUNfuOpzecA1qHxFlYjJzh6
NLFjC+yvSqr52HA+PUmno3kdZHdkE4+ahYReE55e0AWlR+aDsv03D5HbQNIhc3TfVwpKoTvEq1Go
1HWLqq9iHLG/Jg4TTVypyI0p65abMTH5GqUeIwak+PAXRxEX63vmuP+Zfl5ZX/xMBo8De4Tb6/7S
1AOyCnHSjSKDUuuHTFTnHbMESAUn3zIJ4OMhPkQh3ByphOH2gz/zfPz/STDFFcSwjfWb3yO16qUQ
IIMLNfPrDkBPzpNcP2AFsvqZrwXrrkd6tqDnbbmn3oErpHIbJAAvbiOlcLadtysUW24FcLGVUOOp
jU4MJ1XpaUsSCPyjQXU8cLtae2ZOpId4MP4o6opJETASLiZ/6xYDqOd25UkAXD4iJDnURbk29o6X
A2Ge1sBkpboagmMRb0QmTLnmtUVd7cC2LOsyi3phbjS+TQwwkvljYMLTUVn3cYbeWqlYdpks8XOk
hH/e+d2+wjX1TUxUz9T1EIE4hsj+kvNkVXnkfEnFFyn7/o6Dvhp1LE+5GEvkE4yjHohaEA51k713
LVPFcTIuPu283z3cXAwQ162P4XiArQHmzWmj92orWvjclIi6NzoScplnninI1z3/if3WSl6mudBk
c/+s0ZrvBoY1rNWUzIgEqgCPWNmgOclXG5EWc1h5PgA7qaUibm30IEjA1g/3ge6WubxoPzhRCfUO
YXwoXiH/2L65iI8bfa/L+WgUjWSQmvCdO9YT8KZ+5J35O51jOffrrLyWSSVNG6yUT+qdT7Xt1Mre
nw7Qm90O/DzR1p1MhZL06oWyYFS/vY6w5VXJb6nQ4ZuLc3rZNUlnWHRj1MBGjql8PobwCyUZNk8W
WTfuj+5KJCKj/HXhBnJwv1A5rrMSFQqEZ6DEp/wN+sX2Z7n+rVAWKJNbOzjCnlaPQrwvwtGVtPP2
tN/XdEoVOa5T/nAEsTm+FOo0E1o7VDHF41qwpbtu+dYkDR5jclI0GhmnCIphD8qCwAtqvQwcfOJz
wcijTELTlkWZYnBShD45v4WI71PSzW1ueBzXsOOmiLDCP/LSMEDi5KIjsDbEgaAECnZa4aCpJ+gc
QL6pn3UKfslLP1rfYlxd46frFlo/eWQLk/6QSgMSV1hJLfSyKQvoWvxFCEzsN6ukX9WshKV3kM4V
xEi0pPTSuH5mnfRzFXqvOIdN7SvRDKOYgtNAstnioR/CNtXCTIqDQyf0ng4RS/BlEWPIEQP6pq6x
ji4hfj8i08e+fLwTM6EEHp71ImJPweaXVInhzJtVusYk0FumBlbdWrnhlqLaOqGUg9PN+RwUtmNc
L1JA2tVGT3m/pkSske9B8K9to4xu6p9h/QksQqTAMp0ZaBU0BWfBlqpQFprpcKlOl0tEuIEmTNcP
OcR6zggn/rEWHFvSoJFVsW+AJ7dDzAmEa9dHkWAhlj2Py2yE2WtwHZP7XzdVQdOp7lMUNl2JeMJj
Uz6i8d2sX+Dz8kbm5JdcIe5Sk+brg8upOOIAHQLOiN0zsVe7sadnlr11GXvrfJ5I6XXLoA37Hyuy
l0eDT0RbeuRvkHj4TqdTo8miCVnK3QtrQw0tte9Q4P0xxcMbsuVN5mfZXZ7sbLtuibkgyNDA5NiQ
dLAi+4OdxvX+7fggMo+X83q7VTF6hEfpA82QsqAJ1JJg4lcoqdhfwQBQhaaGpqSzcERdZedJw5qQ
cn9lj6wK+c9IkkBqstITGWM7RTEqMUp0b7HGqeQhb3yjjy1Krpl6MJkpbITmS7ekElx1pYCAJT+0
dryRNMmII5rjk1DxBNNCPsgZeNJ8I/xFkpntmEaXBa6YA49st38mUMbWTz2L7ykB8CNIc0RRH3Jm
jarLd8uHpMEl4dshKvAOVGyHcQEuCTgr0aqtsSBSAucPWCDayBpT4OYcpLfnUTBzOof4w9JwMxWp
82PAu8r0bdWnVMNz61XCPRyV2ccKPdEBgcdPvzlTv7hIqOJhv8qtMH3erjVc9s9uzsI1vBVM6pbd
OUAME4LjKR3nqoLcZhPtcNPhn8YthNJrbrm/7M3ZH7uM4yMUcie/z2kDyNOTt9WrmySA8m/QgnJL
3xJfSevG4bwi+OudE0hMrpHjO6uyob6qkZSJARjDCTDTRCtgdBxMkrx5ZGfY9fniXbMyY7vLzWr3
sTuicjJ35Wlh8XEOH8qQaTJmErt85GymUStVEyOz4kyUIXv7WVkTLihdLYsxb68Q+6QCXALQ4O7d
FxgFamEAa7/chfEME/rYx6h5TdAKUJnjqKSkwQENLmGqBuv4Uf4nv2CrgUMJM4SaUVoTidqdPcVV
pOvUB/YyiB4zu7tbYd3BK2sMs0M9fsgVxi//g49I/XyGqDA50UX9IhB9hzzowPS2z0UbRlImeXCF
77RBeRHpKymG6yxEYrdYYIBc1LIbfsQl3qX9kENy0lMhqQOnm6BCLnVpHCMFPK7UEjCYW+OfJ9Jn
J+BZBOhWE2EqE+x7aMy1g5gYzZt9JuiMilf2n+nAJ7isUEVRPhwGRuVKAFBNugwXCGNlGSIldiog
iw7sa5DQi3q+1NbDZcAoywnVrQBNjdWxaW6T5GhAIbrJz0/pUSROnEeqXOZsNZ2o4Eds/yKcfwFG
m/LwwyxYNzsAJjZ8xRprRNVlLlVjJcC7qyOspSGgqAiAZmVoAE7LmTFAQng4qLq0QSjsrYp+TADM
faZpw44aNvZWxwEclXHy396rAqY8+WtifJCqOMigeag9SZV0Mqcs+Wl9JjC3lVkQDHHL43eG4xu1
VtrXLlUD/0xthT26eUCQx/z0J+UScPqzE9vFa+AjOJRJeBNRy57GVSHRjU2RR3cKy4uNeI0UyXt/
VC6gUrec6VbtK2ut6vfEbq6YwBmmA17IhPH/LNo23y1m7NyPYtnRFoRy6kJqjMZtTrpnkji+6NoO
5f2DhY0uwQeKdpUnBpm6gZD+sbtCY2apAkQcjDpNW4H8ARagEzw1DwfzvovsRONzKq4mzFnMZ0OL
zJ3CfWAUSvdBiKko5Ow7D6EHwrW3PXH+rfiXnezkmKbPDNwFOE/WqTauXRnR5d+n7bqRVujFOuMM
e1TLQ55KmWSUZptznUgx7CMTJc7mVSx2cU9Fl4/p3DWbgKHsrAbooGLPUj+/MgjPLlk/A2AQ/dRX
59NaYqpwwzs7IZo25viyqvuzNOEoGpB6gpaTAu+yQkHJApwpcqbkoKFEWZlbI4ljzoJ+yfqSFJhc
n+1sZGSo+V9AhCvBnhAz4lX3V11V51ttz4ryNblUjVeV+zxU8zVzghBQ0dIUMpELfqhZoJc4GDvD
KEDTJKFSLyWzjfh4T/BeIVCUeJD5VlFitP+RXdTYzCMdQI6sRQCOpPogWMQbPKVB88MzUQZA+VA8
0VBVd9XaqD0VQu07d2CtmDxhyDcpesxIHXlP+MLVAv8OqO/WcqXrmS59fS2oROIWdoePn4X5fbLz
c4r6FmP2AUcqWPqnW3OHFsr7czCRCyIQbEXdv84PlvZduSyi1WzW+z+4LMPU1IiyTClAz/HV89uO
EqpbdVUULYbWVTBfZWXaS2jRvYl7pUZXIN4p+3q7pOZUeb+2J8Lqa2mGx/IlcsUn2TdVsKQIsVTb
wBkLZmrYNDmSFge2AvWTQGTLIs18EFb/l7AGMfLwl6xz46NWwEyhPZxqaB8OGeyv52pT6hgmgDOc
7FjqTYSE0xbaO+XCCRK4amCkKs3gq6RIijPZ2IC61lFppkiIHaAV0d7RoacI28dMXSXo8H96SdB+
TtsRfiMfXjS4VfD0xh4N6f/QbqeNpcbkLBxhCkz2IIK38fgKqlBkSEr0+akYuMXWcrfhx8QsMe9z
eudloqe4Mtd355aHPg2ERBk1/Gxl7zgHB0MnV1YVI8QwlaW0nE08HAvniPMsrez2FMmEoAncHvMw
tiSoxnKJ53A93nUdG1Alln5NQlpNT8MkbJCbuNWkT+CnN9shEnbEr/f6BiYF7VwfYIN2SYwSdPhb
4C732KtW0RDNd55a3PcDQkNvHQdCpjfAoqSIbHypPxUKShFLPgNGpBSye/avAiCAFUCW+BXy/ic0
RAsL61Pm9V9HAlHHhW8nELV1M1DVKRqtRhUvjcTyGsRq7VV6JbtpyuLk6kY1qdrfStLl/nw2sJ6q
7JcCeGW7+bANhesUGB98DFLNwXLO3IxYuB/gLw1Glr2TwN0OlFqYRN+phOd7UwsLewSAvjYzjCWq
GMoLd9Bh7cCkpzTBmOabkXheJUeUSYILwV7Q8kfxRLGN2k54rvXZlRT/ONYryxQnjFZSUY2kez5S
6TH7xCO3r5/3lxzGe9OybXEgHc2ZLnbgwwOmbLRC4uvW+OfDQGIFGZP4w9623++UXCo991Uw9+2T
eyknRRvDu4q/69yGAv9jTGYBjm/1b7pKS27AkfzQTg7MRvoUREFgbwFFw8QPbk435mv5d+DtcCgm
wKRvyRFUD/Sv3mRovFbkG5Pov8YTWlCjL45Aug6CGQ8tPB85v712K57CbwK3/4KngPPGawcY1m7j
LeCdeYFS4i9n6rCHSRwns1W8HLgVRiC7O9WOsEVuowfmR3h8NMooK0Pc3JRS9WQsokrHquJBgI1P
lgOG9fATJTxV57d6Lj8Ns0J9mYcD1Z63Dgm6XxEjk3QHahU+8ZAjbmWtzclIP5XcU0E8vCZOStXb
ZpmDXr+HYXHuronrfzA1tN9glWHXczKJF6wu6uaZpVRb6/kbKnJxSxLLyV0anNaUE/N+YuREd/9j
UzDr9dJzq0LkmKt/Ztjjd5PJMY6DTRtOFMVXZpei6He6uAdlFY+1OxSxW18UKQc1Gp8iM3/ulIee
4APOdoMdnupRr3ZPNNB+skzXgZglKfZImJzcLm4vxF7cr0JK6CsHJ7xh9R7uvkTtmG4meiVQ92Ud
X0y8FKFdoQeIK7dZiZilvta1tXSpCkfAPNXtF/B50iMUVPkv3uBgh2fU9MCdABwHTn7P/gNnoG4E
3KiG+opYF5QrmqbkXbe43QGGCQ/78tMAZar7puX50fgB/8qybsuoNhwuAfffmuKs7GG1/gJwA7aY
5Qep1tbcFwQINj0UN0Xxp/Ug4BH2zVdPqSFPkRXgYt7hMtvLfhnLzrcKL861UlIfqvx/mcBX4iod
h/GywpsMUpau4HfGE6KUZvK6fg7lDebOiBGzCdb5F8ZaX9tf5VKEq2CMvL8rc62BQO4DIflJKKQY
cccyev65tctFCwCwmUjOQ8Ntq8efdwugdozMTeW2W3r3Kz9zQdskKrMCKeJZniVhszFIWJVzrYB3
CQ06Dw5xX2zE5QU1c5LHTROaB6Tpc2kQaNW3SuXTefagkS8yfysoVKrBqCTPIJ9p2UtSj+SpD8gU
elu91V+wOPTj0EOqJ6g0pYnVz4mFh58vz4GuNAR2TXKbrGpchldXm5bYO/edu6Xk8TD8J+KPHkni
VgSX1dvggaRIjxNw8brtP18k3K3Ib6RFiamVByUHO5fVIxBEmRRIp8J0wG0owJmaq54cM26T4Qup
YTlOgHpjYwA5J+/gjq7tgx0WVuD4NJh65Qxcq7gOP7miTTXHMvhcfdnQesfiVblvHs9WhHVEXwZR
Jd7RnxJaBe8Qyu0jKybQ4qkJNl1K5jcWV+EzggQz/PUb10YPUzKFuZUG9jqPjOdpBFuCrK5w5bvz
05lVBWWvYPBKBGp9W2uYPocwKBraYTddGwXlEqIywWXpB4/bs/K0hl+I+cow5XRf/Vf/ns04Y6Z6
NUpw2LYB3S9j4H6RkiLcjdvOhBvZdrF8FdjlgYYIaEh/58MgBgyrTa6lN7nIdcLAvY3ETcT00XBP
IarBQGKNLvlhg083EaEeMUH9V0CZRLRwllKGMHTplBgvGeZuUUGm/dO25eWy00LCOKjiPNDvcamP
OnS/3OuB4v4M3TuxPjMEu0RH3CM0CRms3zFsJAZImuvNk2KTTwkS3SKd3JxHq4XHjuWfJemygkZU
I7KqiuKftwb8ORQ6l+pk1IQLRo0y8tt+yUyslXsDEM3qsc7856PwvB2BrtTPOs3rlIrPeLunMDMK
SWbPpiYf2lrJuUw5SpwH6X1JRmSlqLJzeH09KRSq/FupHpT5v51Tp1ALedtaGrHUnRsONyLU2q2H
BOsbajuC08UE3tt2pAEAc9XwfsTgoOt3Mn+L4JpoIjUIuSyLfKUcouMRabCRQpizuAEx0xjItrLK
tlJ6KlQLIw7Zp7gsBAk6bZ/rmZuDxJUJGzlLLc2+n4LEEZEDcOHC7ae+qwY825iwJDCn+egfBbJl
fvmqIdL1rTHeaPTtWPAWdl+97m2z5uCxSP6VIBl+StDBkEwqVj9496Gb+5JoCoUkWhXYm56HpWxa
KoueryWuDewL1gnardrNn1tcCHq+mmDfO15FME/YcXmPlncKn8lwcktFNL42ZIBMlM548z2fm4bC
657W3EOFn+xVLtbqfuDdaq8Q32mt+hMISuLdZNnbJUQVYEFelzukFQ1cQNpQ9v2EfDIkgB3plIHY
TCoH4nMTF4CsPsawzWturwTPDBNAJPd63gzX9NkTI/fpWj4a36A5efLgQf0UEhevMTIrUDCiapuk
lKWUl4YuUTaEVd9QFwAmJnakFjm5+Vy+CP72yNcbzNatzqRKKPInhQh4RakQGH2Hv6HSqXxItXY+
S99oC8MnOP9vA67MeKFBBlv00BlSKpY4htyExi77sNg/z1pmwimpJ8NNm7wcLYJGPNNimg9kKmPV
JUPkBnFF4UwJzTrszewr55zRgMutMiaCkzZo652uaXD+8m0IccBshqG/Ed1e8ZqAknBe9KdzQGHA
xgYukLNLvlq30tH2N8Y6FHn5mAYAWEu2uEocYBephM3wF1O8ySJmbVGX2KvYx4A3nhJDQM/W3RZE
m8uJ4sWbSl9XvU+l6Z5w+o75P+98PlyRaj4XtocKet5fH7uVuCireg1nE0abicPIefpFlrf3ZOn2
nmG+ni6xynaoAyCB+tz/Zq333W3mnVLYy0obXJ+IOVVQQRiZyHqhJyX8z34jQUt7IiQpNS1fiHbs
lDTpp/0PFvpPS8hM5ngr8qRTceKYeL6jxSlv99CiaQyWbIKcYl0i2cbewsNE04oHA0msvS/rtlU4
EPv2c0rWyLhzYjh7PJeqaUDGpgRP5S66b+u/mdw/FJXApY/ijoi/U6iGOS6PUlH+Xgwt2tYWkobK
WXNzbza8ErivfEYY3BDEvK94WWOZMhsE+XijGxArAdXSDrzbW5C4OmLci1VvdE1pSzITKgKG1WY9
+aMuOOvcTcX+rXnaQ7uA2b0RsrEK+ZdAFB4TxCqFMAUAvVovfhyHlUj+6g1hGffMgsaUyaMs81bj
DKlM1q4NAUBGobmhrdBmJF870I5bx0GT/gHcVymRRoFpihTvacDIkhBni7BfXYjwRDoO0Txeg9OW
KGHu+gqae509otJ4HeWLIlj1x1XksZT/3H7F0YrYyebVw1XvUWJm7Nhvnl6vBhQLeOI0O/zdBoc1
BnNd0nil8gEF3BluKdUI4FfY0ojlobS0JrehUONfQ7SFVgC7SxyDS8Y/dhjaouo1fx0Zu4SDPeZy
CnFE+oZ+kdGM/hEiRGJMs6SIGIGY3dpqQFWgZjEBEfcIFC9tqZVGtkg2CPDSCci7X4lXfJOqEZlM
3XHY0KCV/W7ChDR4C4K1TvuPxlVSjxuXcmhNTB1VEn0wtuQrDpa4uQc3fGx5y5uiLSr54GExWWJN
sY4HXRQfrjSkSYodm8BtB3WY7OM4lZmQxzYPcus7gjSW4DHogVApn2LfGIXHWcz+J54encNb3nsn
xJwWtmsURaLFtC53/WRxO5JypDmIj7sJLoBluIeLdJyMV+dYWwVv+69uEQd2vZZTvw52n/KoV9nE
l16gKGE9J9S/0RbjCl4Lee2yYOCNNDJK9JZCtKzW9rETlJFWKKrtf43LUQg6TR9u6ktvs81dwyLX
WQoQzx1cMxxx4fIIUlrcQjKMTxA86w1g3fJcvYAmJAX+8EsbS5+TJkRjFHk0gOAPixJ+zWnpGdnU
8nfhQWpfJL787BofRA6B2dDA7+KAzwcmTlnpHX46jHaFrZpk2obtADVWcoEE2gz3sDmyjJ1jDMzC
N5ctc242UObqrnV6+Ylbf6Ayt5sM+vzqQiXjkbhJpV8MvAAp52ExVzA21L9SP+Hq/53Zc7YyChbY
BhPLXFExE3oI+Egnbl8bIWBZ+u1YmOkMZ1Wa+FFdgJX2VREABQ0jtp5MW2xMGvlkSCyujj0Rbm+X
KFY10+0rsPCoFFYwnOyhFB4SGJ++1kjlzVO+6+NaBmMONzd9RmWY72mpDFwzsf4YaU4YND9VcZFo
DwaNO3ANa6I+uewDdMKYlH+UyamauOdcKAL61u1QCySzqwloZj7ggKkqWCboAFmBOGdzLBTpGhUv
9DiEKZ6QzSkahLsPzAFB/WCkeZkWTixj5XCFAdz2/pWUjVtMp2DAo1S/CZPiT6HfPdEuqmravH7E
vGFzmXI2Eu9tylgGKs913eFlijtPrxGyze/DJDxWibRaTMw+9P8ay4RzyrYHXn876yKHodLUPl5d
l+GIxNECoC9H3YAb2AN6UZh1OsQSVlWAxJz+3xKVfp+ke9Di8s8b1qlIscEX/okCJmM63ZgTjwyI
WIm+SuI0E52I4J3Mq8qA8HfZtMN6yXCn5F5E0qWQdj7kD2uCl6ngnXbx0YoORZKEOmWoDtk6ufbh
aDJ7eLfxJLkkNHl7Cq+PNsA8cO53SH/qIDQ++sBAsaWv/qaO12MbfmQ4DLT9JKglVzUClMD689jk
AsI7yWrFayJ2UZK5zGCZNamg0XbifJ7MwDgOHl8DDrmSEENT2Ycx8BIRVt/Mnmn1/Fth+3+j7Z2+
VLWb22gyH75fdt7ugwunBAW6gRU6NfTUY1kmY9dgY9jOkUPIjRYhZfKh4ULvV/ImQGNyxOYy5SHS
HuxdQUutpjoArCj201f2W6zmTqhxPSVSs+wTrD72vOmkZgNnwQwZRNndeet5mde0cC4K9IxYa2rH
pkhNZpGylr1GMGM8qyQftuajo76QoXrmygP3Aasa8JEm7TdinudRuhyoNbCgJAQeFafbwTVnw0Lx
2Bg23sXnbsPZQmQT8/sqmQLO3YMGoPK9JrAml2Vw2KWTmctfoUJ6TTy7aSJXJS9HgqAFTSKoLts6
580m/Y4YxAfIWfepbHyUDzvuD20MidsRoo9u+KmA2BJpQVw/Frp/ayt7LZcDBPE+dJ+G6zNzE7f/
cufInWCopY1Shf8+uj1acWILAiBdNEZETbkesf851WwqW7fwZ5t1Rvdl3mAtkPt++C/Lcc2JMgoC
+YBonvy/CZotPz7If0baS3deE25GPLFbH5wuyQe8yckSI71Pv7NJGPPoWG1yb+W8oMbZPNpKwQFz
pP1ziQqDtJ6kBlGbLzqdYCRS4C3Qra1WQq2iMubZtShTTKZ9gBiNKWcn6IlVmZ/+bQQ79OOyNG1n
T5cGqz4AFkih1bn0Xp1dYzVD2HFYRTvQj9TmEu08KXxMq/xpc8+pq2rVv+1C589ighbt7Ynfvrck
oZOtM/ppTCAXlypcBYGUk8+g1JyPdYrpxzXQIwFk5hk3cfyRjIilx1IwasoDtEfna65BkbXntyTX
/pfngQ7rUwX1UO06my5/TgcomZrQRhG62jNDm6qZEKhkSpROEdQWFHnEd5pLlE2tVcjZ11OjlwK8
RG55IbWTgoAfGmii8UBtNa70qvWq8hH6jHuDB2JIr0XFeRtzITKNF05IyShSG3hwf7W6BdQhwFkf
Q+KPnrcd+/5Q3XWakrHAu9kvds/pHYAiaGr13oomQWCnJA6eOvgoQLXTlLpjvlnZqYsc4uf8pvNU
EBruriu5AjPPgT60NtdjdOJJfuSL1EvJ4+mhdNhWz5bXGGTcGqlsVi+DMNClAZTg7xGg7SUtwKYm
gV30Dla6IvXqfzofDyPPM9fwiHVxJzaoDvM3NdVCfc/ESncbfLorNoTChsoICMMeU2awK0TVWBJP
VTd1YA//LWKlvwZzGcD18bZI0/u2QqShGMv2xWwxXyPibz5Z5MvcYuSp2k7/Xwz1au+IIROzyL2t
zCLeedtHQr5GDPegXgDFDweczgsXs0cgzVIb3LJPqYTOLfVRs1FhiFgV3KLABzgZ7sbKAcv1cwIZ
2ir5ZPZgViukyiJy0rBRbuNTNLmTk+xOznawur5zOh9On7wbXavVDf5SBuzIev+NBlxmP13vGC0F
27ASzSNJNl2XwgoaHhkODcP2SgDRJca71qpIkxsFAXbm4TYEnoA5x5Z4MFksULixNhys41KytdX/
Wr48/Vg7Df9WgL8vRXbuyTS+fdYriC9qD3iDmuJlmB7N687U8tI91cAO6wbu//q/v76Olp9BKpQ5
IgAWwQAhtvFTWr3lXWFC+Eag5Xl8sgDEaVwKFuMUg7nZ5Ipj8SrHN9xU/c+OixkYFG9iwWyIjzKh
5WPtiW3iyZTSoz8Qd0goOgdForOJY8ruRwwnGiQB046dIlDSxr5nm/zrRUlva/8bwCu9ihaG6CoB
mHotFEyGB3oamAN4zeNIqdVMhDD+KK0NFwQNdDtl3oAjxroa9PfLRw796ftZrw9Ozs07jaABCboA
l9eKBe7k/uhXHBzqMk6BmFnHV5HTqxockAlQNVsJsnif/BBrFhvUpyo+0uw7HJArl7k3B4/alq5P
rkJRExr8SoDkbysR2hrrFmxTXqM9i3JDqnZKX+4b515IArRdb3I+5gRamfjJXoJN77pxI5y6c9Tn
O/JP9r1zr0JTHBZFchzp5Z+UvCv3y5rhrw7of9FZKKb3u23jfmSaQlUCBe4TpFoJr6H4vPstDnJj
2rGghgLP++jKuuIUI2QeNMgkKBRZrzrDus+NMs9+Kn4i3l7fl96+YwlcDPc+ZoaX1GzgUZ1PQbin
C0dUqnXPKmD4FhWsa9qXPecYEhJ3EqAy4IL/cZduu6Tx28Vf9e359Ane1Vavt7aouCrFfQULjUiK
uequEmK5xyexcqd7Iz7a9fvu6x2hyBMi603d3NaOa1wIc5Vdt4fIxDil5djc3KCqdxS0tUpzrCsA
iSSN0anI5XLP4ZJXlX0MZd86MKMwjn10DqOqPR3DYKsypMSP6t00PsdpOOX4VjuRSPflir60cUhT
YI4teo/sNgE6ocg3MJc7QC2GHXIVawCUV14vR2lHDEMdPia1PzPb4nCF+gj8tnfb8M8TfkzAHfys
R+KiXz5QMwB/fRlQeuBnFD6NDRgcF4hGtGn+92bCr7ZFHC6iaEYNoSdLpKJhYDhizKAMoSnMYdLR
8tpw+UGJV7wc8OPh5bi8Ez0JNZGkSx85zGpjcSO/bADsLnJqm2arZPviv/uOra1UbPghgIUkYZYw
3veoI7qom2zPOsd5YYL6dS9CJwfQ7V0uDjIfvSLqrzq4WF6gtHLZSPZq4MNnVcZd+jJaiMxGzdRt
tQNv2fZZiIowcnFT3uFArihCWOIkFIARIFxSge3WU38dB8LDtshBrstYcSOoqYQdGNhbJuubY8fZ
U0hH+jpvI1YKaB4OrnuDmAIF+ib7aVhUT7i+Cb+C/dmHTF2007u9KCUt97xK/COQ1wrWx6YDJlOJ
n6y9A1FrUPlGO0hfL9ctjKx+wPkCMDrMyo1AB2uGdhewHJvZxJmM6A1MfCMImBaV0Vu81drc52v7
NDLjWrmJ+Lq3KfABTx+L+OPZVfmyfaVqYZGiKkhNs8OmXta4aKdZvhK5T55BHCtQogjhdImmRQ0/
1mvJExqwv3oQhmlFsHcDDBRMowniTQBTbgvfb9DavG54KkVvDU1pZ2XsHGaobq0oupodVMVIe1Ch
r4lXBbSMAMXeaQTuO7QyBR4suxQ1q4vVTmIT9h6BWMo/VSKPVQ51+zJ2FCOiqG/M7n5NPX2Zvb1A
8pR9GCmKM5eKE26BK7ti2aoqNL9udnHTchYPTazk8kJrGHkR7u3P+InOjXp6xfYqd/JFgXBa/hb6
8F/NtyGWJBoiyQAZnPVgQnXxbV3BkWW5LuX99l+tgRanSJ27aflYnbmz9Kmuv26CddYzHYspDGIJ
PFt1NXWkt4eLcMw3XwdK4cShGyuQ5HFknbcMiklDGn845CvxJdiiBDqQL9Z1f/WplTkRUNtFzsBF
U+VVc/fUbs5PzloVn/kTYPHycpfAqnu71XVyzRjJyRgwUdZZTlvh65g+J5ogNP4ODJyE2ACmj0fi
1ocp1K4jS9plbyOl/hn8HwjvErk3il5YAaOnJgIrpgbUV7fu4hQg38jzsYhOr5XuZnCGIuzAxxiR
7q8clic99K8zm6Pl/gdIAHALzO+DIvCHrAeOehICHKwer5vqgc0m0hDV7EUFNbUVuuIulJwqSQZx
lNdaw2my+BgzS+t6/b5edtIjx9VKYdnlwC1Hqj4msFy9RIsX97FMSWtf+ZfhI2j6xKZn/biipRTN
YmVCjbPwQcGuhyHZg0tflWb6sedaaqLhUQSJcVDfRn7sbI5A/anhRBFaORmbUg+fV7OY4l0xafZh
GRcQk/KuneLKyG+SVStX2/riIxHfMHAlzw2wHlFtlttLB6a4rglo3Ed0ZsEuwRQZThXHU7Xxl+ip
FZ0Uy5SPwoP8guEaGgAI6gNElGF5u8NHFeWzsDiKB15q9KHDzKLEsM1m5Twnojybv/dSVvrpkT8v
pn8EgrJ0MVie7TkEsn2V2GYxadXgIV/DUaeOcU/Nh4dUvqq73mRjUwIUqUVpMEperHR4NiyQefFL
ppBOeN80r0cd7EpgEVDNCWUCn1WwWsPKMWc/dDrNmveL6Dc0c7Cy9srOWOsHqE1RjCprSVuiz4V1
zrA4S1eSomSDmTSY6OQLiUeYxiA1RodxZfyY4O0LUh4lr+o2oMX/2YRK38+BmxF82MsE6uTe1lNS
CHXHGwMCzDxtcvx6BnP6LES79mSgmOPNpEXxIi5DM7AAozIIVakS9dwDoycEO9zJ0F7qoL0MkVGc
GuiVeP2OBzxIhPoK6tQga321H1UVPQ7lXeVS/V0g+Vw2tQ6o9V2ffBKgQ5ghRTKx9UxjTGX0bujq
rQilCsznq9uPbwsU6n3luYypmj7MHiN80S+o06DD6QFZ1oiyJemRzdaeyTZOs45SIazkaUQDfPR5
FyscvLCOE1h5q8ff4nqieu3xfIFTj3J6+OMfMygOMxVfeUq2RCQyrZ0KwLTfzL5BBsD2zlrVcVQa
Cvb8E/l25Dc8Ic0Hlf/K/K3hw8ply5jirYQKq3xa94LVqukaQNfTLlIcgyaQsSH9KmiRQLaKxLnk
tlIijX8RnPtNhIlmUd2LEEkEJtXkbQF3MxO78e7/j1dQF8Vdr+ij7dwUEgJ+KeeaabLOXUet0yLK
13ydRXE9tSezvQYONzY6x2nHb+OTftGmPhPiv0XxjXqWpz2OIIUI2kbAste46U6jOfHJv/ij9R2I
q9TI3KVPhDamAYpFzzfhS1LphUa0E09nutg/Rrm3auw1RUubx1TJck82APSrSjGaGvoi8z98Fait
w6ZLTh2PEf2Z8zMlnxhjR5cDMsGQKJ0SbqotMjanXt7IjaEzIonpkK+LHXz+NrGQuEEGs9ADQ7CS
s5uwpOdiD3v3KLRXVXOi76RCc2e9PdmSJzpLYQz4N9vWaFOoRoC7EvjOGZl95rVY9z650dMox+dy
PM5oOFffQkBzVJlHJlAa8qZZxjyqD2rSCyXApT79xT4bnA1AxMtEsYBhgASZXs8dQYTrspfPPOXW
SiFNGBp6amsGNGWYldLtOtgdaxnEt7ErEntnBaJTj3LNpni/exrYq3XxvxSLvngpkU1OUAlW4cJk
3p1xWVQgucE2yc4CajhXOuy1Dk2pMRQAhVB0ATxn+dAT7DXWWGpSmu4eMByNqpXF672/crdC2nQz
f1E1u83Lt/P0mCkD33KSXM0lmQ+rZRsDcfx9RJCYfiwuA9ck2xNx76ruBO5SQAf7XXa+v6YotFqs
v1JpLaCGXCZN9juXwHHyY4K2EXMu55a6aUhYG9GVBU68JVYE0IofJgBWXYddioedtrpbVdgtpetJ
xuCGumhQkcnobLXD00/YkLnEpGs9Dhg/HQ3aXCzmkbZgFjD/PCeRbV4LvdYeh2Md5hHErzm8HoSD
/e8/eB3gz3MMIfs4PMwMUYJSo5HK2tbwG72jCRiueotes+3++eek9qGfUfHVccUbjkCK1wZVAHp0
DHnWOYVZC/sPhLhKqtOOeSMaKGO0J4lIYou2vppy1u2yDoxQmK97u56G1dy+UkySKHpxKXTy/KTF
IkUk6xj7yfMZEbFqz0dn+Q3O83LrGnHzrRapNrqwWz/ndrU80GIURuCzeOOoHrjvlNI3n3dUElZh
ajJVR2ujsxEKpMFpRqfhKgSBcFJ11DCOuKKw4UWUbop8XyF9h3EPR+UAwbUwphOgfynIfJ2sbAo7
+Kk4XHQp4uKaAj9I10bXvyggiuwec6onYtMIfbCWvg3IlL6gMBjiidrYyLDTAlGR0yY8w9yq1NFH
5tvkqaNp1iLTvYxegr1J9P3Ho5i5WlF+xBTYiMfX4x07i3P4CibDTqslw3Gf37bqUamvI7CVuDth
vjtbCMqaktBjT8ycIf0GIHcUFHuyK9/WYEAo2FOKRGKLCqbQdtmXzfjg+q57d36xSRBOKxtVqYz1
qTOgLM9Db841u5dr0aOzbvDlzIqdKUp/bI4lTqNpWzN7JQuecRTEHLvB4QRlCgrx4NKWUowb7g59
uwSlCEMuNlHq7L6IcuSbGMVp54zr/athD2tKs+p8DyAVdAQbFcx0VemUoF9pwMsyU9dqn7MUZdCj
s2HZ6u2bumus201JOMxSw1TUKp22xKXyliM+AxTw9EeBmkud6TumLa+f91ghfSpOQwpSXqgKVeCJ
ToMNmGVkfpy/N26DNL+pIG6leKdpn9Uk0w5a//l8Ii1e6//rg4QkVxgFhCPr+BLOtf+r4YIttyY5
ygGdIv53vhrvKKerh+0DKR8BLZtn95FlawsftRsgMVJIQm+1WQsxxHGshKHATWylftyywJzDPeWk
OOhFlpqLzJTixv+XU5ZKwTGOtZdWr2qHxB2S7evfHz8XuZALxUFCGsKP+F39gWYgi6JUnf4+Jm/y
QMGdLYdwtKQAqd+ufkBXr5ykxJn4rI+AouYkk7Pzg0ZY7Wz/cQUb+dt0xIR13k6+zapWuGo1AkOK
B6xAnXX3leuYHxVmJbrg6oQralW6cxqzFMutf+dH1cH5Q4Sp45DyandcdYuD2ogbXow0eHtNu/zL
/Dt31BpTL1VkaLyhYwM5TPCt8n5yeQn7/YCJZbRCEQegzzUXSk/QZmR583QTp8rnResU/mjN6xMb
eaqHgnqfXML3Z4AIZ/ruZ1F9rF4pQVVn/okL3AsxXkJjwjCRW3PwzI82dmien4IdxzNsgFvZrGGM
+wOJY8j8nd2Gkd55SK2mrSVgwa+1sf+sqweD0A5pm6dBqQGfqsLcEWhc5ymZZ4UGPbs/XW1wuW7G
vjm1fj2goSPILkXO28fcZzq64StV2UYNeziuzibRWBzCczhYu3WiAsbh7+/xQbQ2zbzWUzya1ohU
bt7uTGdwue7pMmlrlaELR//G/n/zXeaXbUAXX5dI5EGseziaBlcpiHt9cMF3vGtFspRoaFu5iga5
NCkvOohpQ1VCwzxDJEmr65XgNKgLTXPblhg4jAqgE7n90ZtsFIPKBBy4y+5UUWIodBNRoF1oUNNW
BN1OOGmcxrO2VU40sHzCiWiX9HP8RPvOlm2Nb4Pq5HSoxYU9F6qmHBU5iBVC9lYcKcQl13hcA9kd
Ys4GBUtHC6mSYDnh+j5PsEWBBxEd8dEezUwq4sF+j6Einpy4YYwTrCtv7JEiXUwPu7N/QYtXsRa3
h+Lv2kN9DNS7+rXGSC3M15td6wLfWGSn0kd75SPa2swojJveAQu0O4U1W/f3XJmGsKICqpIRcLFi
XGAZ47jbzlhUuHgNQb/4E4ah3sMP4A7XVYpVcVtGBI19kvuM1+9RcYx632M+Wuecqo2jDcmeumlG
ObrlO0qUmvmpWN+p/b7ZKWrGhxAMhOMo7V8YyK+btPG+Qkbh4BInLxixbXFASiAIr0196wukz01N
GAev0BzjMZViN3sBP41+I3rH9sg6TsIpU/UBcYsrVbQgImJ5D0Y7p1VujVWT+2DVEz0G5XjnaE/X
KOl3zuzsD+uk1RQ4++LG/L6jeFS4pSdQBTHmkOAWz7zrLFOx0tQIOr10sFkco46d7EP2102Y/xlK
hv4aLzCwu7JaQZdV+Nhbn8krKkp9pqtYR/y+/zx1NRfeNoSnUmOignIUxuRNgh6mMTxvg0xtLK2X
Uyji+Gne2mXdyvlnDEAwxaDHT37/EgDDfLHljg+d0V3pySRI3g8fsTaztBNg3T3yqL4dIdy5m48e
b0VOVSmDoS1LiQ+5q6dcvePCL2JyP5xLFsE7AGtqFERr+uOocwKapPxlBW/imkSdZcOyeZN17pzg
SksiSCZK4PwfklkkgrPHNfmE+4BAehdTfPDaHnVha1r4gkfsPawp/qzaYqtY5EM5cEy3yp8++4Es
afoneUnIEVxhpSPHwnyLatIR7ysyoOTyGL9B3D/3JuwIOR4rXeGl8sJDyMDLsa7En8fF++Ich+nh
68XqOzsyCBpk/ZGoyMx0pijH0flbC7BKnIL5zgR8hc4jtuaxaX+yLwwfwP+7EJLOyH+0IL+NFnbg
t8YCQ35pOddn6Ws8FhYrONhO4qSTDUda2E78MwuONDJXTltvWohhoSZA6Sfi34a9Sn5nlgkP00HN
vWZyJz/g3XkZpFBtJkVvsd040u9NE4NA22idQScZzlUulvdjh47FMWv4uJbB63+i+ZzTDibRP5ZO
3e3gnvx9d71DIYPEAg9chGnTWY8MplzNS0eibvSEjzglc0hdxVJDKIM8s8e3IjXDKEi1ooJA1lo2
6cdUZ0QI/xmh4FJJ62sTWdqOhm3oB/ZPG29IhHL93PFy8wcnHZFLp8MWVEuOeDCM67apdtpLgY0X
425/he7VwOcpIrycJCLdRACpSBJk8+NgOACUB8O4LVmGbSacDLzIy2SEQxLK18WbzW33pw2rnVou
ctqD/pcK/JOLv10gN2QjKwGskIjL5WmrqC7RWnnu9+bqVRANCS6RiRUd0XKdZh3XDdBOBP2ba69c
U3jt1m1X+i/qEI7vhI0I6OqlvUMgbH8hzdC/AAeKu3zmci051mUm9AxV0zTWHOjf9Uy6M/PNQTqT
JXTskQTMe6AIPRFF5/t2Nc3NMws5siUDCWUmDeg2WZd8fRmYxfgJL+A8oiKuVE24eK4Mo/Mxweaf
BIxUgtBku/9JgAapRYbKGXvbh8buK/aEilibFVyN2mvz2pqUBKt4RetB3JhlJlr+i9A0BOYpXiwl
F8XSkUOfv7JukHlFuPRpGq4hl57dGDTAVUaU/zL1sxujdxHDqAl3C1ymMoUjI2ZF8DDCd0SXUz9X
RgvRJyZaQ58Y/s2tyjjiPNCouCi+64QCfv9e8I8ezFfpFyxc5Yi4fjbAqK2ECgdPH4l/XFxgmj4u
WzC+XYQ/NnUtDnwsAZFVs60pl1XnJe2QRJTKcm9oCdJdyZ5p1EW94Eh66d4i5vvLudP5buas6GPd
2Vkx+qC34jv32YMLYzHN23wAThDgfMrgKrS+s8sS2PTNedSLwnXRFgC+gA/8tXXXMWxGyEdFdvpq
nbF0EpfXBU6Qe3tFBm69glQ0bDNGEtG6Gu804PvgbLAkCnpRgWApjjZzPuozey50iF5hbhRT8DG7
hbaE2pyxTHFB6YTBrzhs89b2ncnBLR0jsRu3bNlOLgNI/VTic6UxuOLb1ZMY+qauEQgbObsbOTm5
j2avnbl43pR91vXXUf0qsGoTIYVNlnuh6+djgfIr2aqK7p+ZhaSyLFQC6vSwXkeLbAZMpeUKFimu
LDRPa9M6t6lg10SC7YQMG3giQswKk5ual/Pv28Z6MCLqoMcselNfuS2K78Hb8wbX4rO2XD8GuCFR
R5T5edOkOMZV5VnB7CzF2LYYKBfxnWsiVY554wK15ipBkryaA+3dbC0tvCFH9DlTkv9VqGAFU77z
HtbKu0ZRoNwBLliZgK370JpjX0S6TqaPPjOAHh6LaBHIvjezU8W49C+hywSSPxS6ljidApZQr63B
nQv6J+PZ6UQvC7rjxi8cb754IW5v8/ZOdeiWuOqEISjROPNbLqOERSwGQIHDREGt/XbjPbSah7V0
yrTl7JbFVZ9AItOMag0+oS9fT9KgaElGZ0vkmR1pNqTm2HfU6zOtynSFxWEZ45cjbXzpOm35uFR+
hz8w/JX5G9kiXkVxUdbz78EdLopoevABIva32fdaibztB1CMqmj6CtXPwv7nJ4vnjeLNWSR6WRP/
YZuXCRKjTQf4QUCNHqa8Wg3KQseEdBrbZgeTmhF1L/ZuVzGsgVrBTMIkDmIDOTa0FRHhFPe8WqEI
wnT5IUg4HmmTHB/Zgrz38qGnhlCKepEM0Ziwgr1YgG4Nq0vbEqCNgckJHwjc+14JSBu5/e/taXbV
z/ZdFlY645He81pGbUc9PWJbHI7CCSB0bgmu/YjTkM4rZ/Z19X0Qj3SJikks09pbK4cfXdVYBzq/
JvN6f8ZRuwdQhcivKk+TvZ2iA3WBMQRE2fT+N++iSdAW3VgSIhwGzQQPZERqOougkUaVTX/TZ4Le
Cboln0jC0PpRYf3s8R0+anVTlHA6/ws3hSb7yIP04Fw7skYjgMMMvvVv+mGSOfRs9kLvrLZyKT/f
dAQAD/O/tOhH+6tOYOKWSXDiTorkw7IvqWNyj0FkZrMLx68w+uMjgjYcx/gksY68YTwi3RBOwp81
xn9SZuWJ0v89b8b50CsZGqw1glVSV6aOSJiNyQL++awLFuy5vAgxvvb550WNDpYbU+rohWICQlLV
KPMbGQ+BIx2r7E2+X1bIaFyIrJl4WC8IDt0gL0y2kSPEb3mQ7R1L6OCpFleeN5rJIw7Ws6laqT9d
ofJ89A2QbxOV3ZvlqpqZJQ0F+7RXMX4TXBhqkPSE+dmw0IOTDxjuedXGkvODNA6szDKXuH/k8JlN
AKgEsFGGFA0a/AxEgE8aVyzWAZSCByXlfTqy3DXXzKQdbcYZyIaOERB6Fz/CQkszIXxtmkwkRVLw
nECb0MnYWA65K+fWHumkyft7xSvTtRd9KbjlErXQnYiutdrSzrdPcigFm9Opa+V7l75/XaT+A4EK
ab7dCgfe95UQM9B1FaLhUkjt23nUJtLaY+CiqFQOATPO2puwSFVrRCRE3OhXfa2Jp4QTnWVqmBDf
A7SfIYM+O++mhBxJJyAprJPUedBrcqY4O47jh1NPYu5R3aIEhwwZ21AcUwm61gwWE46wlr404XXo
AznSVRZo9wSCcrFYA+j70zzmwxATlxmfeKsNS9WZcrzZoAMXi1NZ/qGKgDWqb+yHn/CHdha6m9SP
Yg1iDxOaTRw5YBOo0fRwE3Am1Qj3wg+dRkOD7cp1GO/0e5gp4kDSmF4R7qiHdrOER+fF1rzOHLx3
0AGZ+L9RieaDXBu1FGzDsZfhyYMjgBtwOG+/K2+3U6XZca9Kwm612X9GNyZFD8gJUFBJ1RaYd677
OquNDVbQXZacjxw0pAkQhECY1PSj1tcrTrhNqcVDcBL4H3Aw+deY9qG5O0iWXj0WjMVNI72kqG4t
MfaHFhJitbBT9Rb5LXaImkQP90pPTxqFXgS6csDaoGv3oUs+ThuhSAoqmLpB1yBAbKJkh8YzAzI1
gLKZkjQlShxx1FoDvRVqsFS3vLwCHXEYDBnBQh2Zh9dIW9znvVYLBwNdFHWt+i99ShdNTtxgzQRI
ORc0T1elvhnh/V1TCcX1unbbp5vEPkHDL/8NuHvxXanp4fxtBdxL6XEF/5xRR1UDk3SqcupV+SHS
eVrppigUM2zdkFn/EXhZJ2u13/7FM3QjM6Hb+S3BIAzHCI6VIgr1SKRp+QC6hBTm5M1SBqdZGrfm
qInSgm0dHAfD9/Duj6QXA1l+CGT0b/C9FVCb4Q/RTr/t12q5AjOXLsEmTXNVKZC1s0+dlxjmJN8F
GT2rmJkM6sT9s6epifUdQgjmeu1OlZ+nlaU4ZB+8HXeDu2iGqZLVm61yWW2zecwKEm+PT/h058g5
cpxL7/0a8gIlPPqrstV+Lfc9qw7hcM62r9WhNEMzq+C36uUQgYLU1ftfbzMErXPoxA2DpYRk8TnK
qU75GFFpajepfh8RUfA9+FCpEjYe8SQJjz9UYbpXv1BmDDMgu008jtjn57z4dpfJSObOGCDkPiEM
eFaQe44ihr3bQeH5jKVwXz9jIep15PT7Aflc41t5/e8dy0Xj8IgK3UB5AdkmveTpEF83WEN0W0u1
ZfGk8oFx9kjm1i1ltU5+zuwiFJja6dSW/kgc+qoT6n6MpBWdPFVWBvJNoXFhGPK6kUXFtpz7coJr
wEHOevb8ar+V6UX89S2GahhntclZsW33LBfBW1Ng9875SEq8iMYKIFEO+fK2VtLeHdGuWcwaHuF1
FoJnXzbu0Eg4neWwDvDuEZyoxQmoTY/tJb8BnCuND+ra/cFaqnU5HSA0LRYyg//xpCqA3YVyVFzN
moCNS+2A/kitleaQm1yCVZ9Xge8nh98fWCn++M/6IBhJkMT6szfsD45gukOAJyCS+CKbq+q9lCaQ
ngxoTsWiDG1xgtK+S4WX/mHpWudpo5jlppe+ZMqEJze+9mMtYbxxZ6AgRKf9/vuy2HxGVW4i4Ya5
XsmqVetJ9IuEPbaSd5tRfXrFxmh2areU809z5IB5XSymj8xDOo9RWWIOXVetAc2yp0jknmQCkafg
mCV6Dtd0fk/4o6jqdd8MwHWi/0qG5JKIN3nu6rysQiQ5XYLH9x5YhRFQTdaiOQaUaEZNoEyQFCIa
bERSk6DmGMVvwk/DZNcjRXsdFNiBp3GQHCxhuOUvrtO0j3x6UvVh1tiG7QCDXPNV4TfRxj5GWXTK
S7O0GAPe6+TqUR18NY8/CCURZ5/lBcdANzt5fIziQQhAFxwyl/PfbK0If9W+rM27ep1uBaMPR6eL
EWUwUikTxnkZcpVdC5APvCrEWa6ABvmCt3umYNWX8d1l+/cEwe8xPo5wIMyn0LweEuh2RQpueD1x
GCP48Pi7RTWx3w2edz+p7bs5LIxgZ9Vv95Kz1ME3k6QNU9y6ueHU1QTJz+qKRPpPrcAgqyXnmtVj
wr3HqGn325YhZVRwDSOokEfYlhgoOPtE6Cm3u3Afk/xi2aT4w0zz8HiuMaoqa3WXPj9IK56r27KM
2fBX96f3C8YRWM456SnbKPW+LBQuQmJMY6D5dxyHUIzkIWtvuf3AWkNIJTa8kE9Zy3PYkoOXrEO+
+nGT8mJ0ksdSBdGb8tTMMDu5knc0juckYs6ZE/k5amJPpiMyl+raW3+fR3MHF7fBc5ssJZShhUzi
4RErhZ161En8nozJhuxu33mD6B7GOAh3u7y3JLYmqOoqYznBtVVxBb/gS0GtQrkN8UHgqojawBds
YqmmpawIEBBrM0Hy4U+qUds9Jvrhu+rMig2ZOFS9vvQ9iCSt/3MYjQtH/lOwgu663Hu1+B+kQz8h
+0PWuM8f+iyv6jTFUMx96joVUSVG6il8+cvA1NZd9T7Eh2iVoQ+AyrrbF6LZdV9TSD2B7Lb3tdgK
A62ZtDRWGcYJX0aUYGYHMijQ/iqiEtEl6eyzkWqAxOkK8iKNgNZkVTv8X8BYh2SHSoruiq0COWkZ
SwIOHcoM9uTjnFLB28t9MgitWoWPIPt/v5DI7/uRefUqENq6dEVHR++3gVRq31e3ymSaPRFXOtr9
fMO5M+LQD2DDJPAmFbcCAkCOg+fz7DwSvh7wQ8F1sRfwWskhSWWl7PS4FYifUNINwdtaNDHxoFkf
0a6jSGgPBIoeh1s+7I9sBPGEGbOogp09CakwXhrD4X/wqK9xwqR+QhxuUoPmU2JRsWatF0EuWKmX
F/cKXBGZ1oQedZE7VlT0amZqo1yJPdcVG8L8Uw//YUpAGOdEnwHC+BooAma2btNh7fOXKn78/Rt+
9zfvUOaf9qX3CiBZsiM2hTX64u3yv74DUdTdFxutu4iBtMHoWG8dOB87FZUa5n0zzJiZRTMUbA/b
Ju9Cwjku3ixIuq6DgZyH74VW6lijEHzrsDqsba+/+oPs76HocbBGJwluW+nqvXP26Y/7b2mQ2OZ1
f5qeIqUawZTuEeOb0EFaBbQkQpGBpzan+pq7MLDEPPenuiJsrJDTo6mtwd5baXXXDOb5nAnVfIAo
JXKTQZ4u6pnbHKTM0RurJzyFZGVAGfYRP651L4HaLX+zZiJdcsBv6MmFXsMPuRvhz6/2ACmMma1w
5zaFsXwf/73AKXU8QdL/QPj+4c8NvGxGbnpyPUySj9izVsG2Zg2Hn2LeEqIYie/uHigO7GaK29Ny
BF915uIP6GYIggjj4/Gt5e9KUcZLwuQ2zi/w3UjsCu9smGleAYUEN5z/OwB7gdgZaW9sdneMU0Ya
rAtKH8qKUMV7A7xNOhOakiWfknlLErxXLPHTTdjLb7HB0M20QB56EhCqzRYOzbvq62GCcnyHN3wW
uDkdXHUxBCGKcFyXN3whRlS8XMh73OvL0LYqJewypnesTdcn/4s/DOGxAMvug6BNbAJOYhttrOWs
5fxgZBITTG58/hT6Yr0SragHfjtszT8bCRJzr1JQFLGUazRlCj4rVWTSdF34gIUfg0/htjBiGNKb
CWPFihad2PGezQPK0MnuC4LdhhYyMCn5FFRl1ulafPI10Ixm9xPNjSno5QIKh6lroJEjv+pZOg8W
ohOxehVT+WmZY6NMWv5KUBvUplxMXQyUUjSOgedJ/MRBV42J/s/PMfZWR8Oum6o9RGezzElYkaRg
oEimk6QBLkuEM/A2f5UGsb/b97QT87f75rKtaaL0fQ6KUIDn9C0YjnpDLUASMHE8Zw/7MnRKpNHx
ddXHM4+MSug0ytK1Qo6lUVQ9DTtatllsNkZqF8DFeKiz7Jl32RdBzV1V/gtii6p8G4LmbfqISwLx
uuGZZR07i5q3CIHTbdlmLJICOx8YXfBVPuJ3YxDgtyo34N37aRdARK2oyPwXJ0t04U5joNhsQ9hu
2WUCuBsHjWK+xuISm76AI77n0UvgPm8X4NzDOHfViKn3OBQY8HtRPFIuMsor4lnoRG8sLBzl3hA1
GqZvi5CLZXUabkGhRfZXkfvwJXfVYtcgQsILL+pCn+cTCRHd+Cer+pJ44IqPei6w5Kq30GUkpYO/
goeOCVcp8jknt6KNw5R5zjA72Z3KBMfW2Os27js2CkaHY1ag8NWMO65R0QpDvoM6vIt2O6yuDvsl
iWhAMDxTA/R8KviCb2pdm3629b9G8OQX4qPZn1lwRHdchJgSyh7DWhNeYfZjDsJE1Gll435XpPrW
m0mVfbu5imNvbGO8eQzGuIqIA3ddJAXowHW75XtbMjsihjdOvKOaTYtZKq+AJyORHHB4VsSiun5h
6G/iMTMEXrFrlVjaRr85WlJ0+J+5CFkPsXgGuXq7UpOQkSE4bZ3WfxgGVtf1rXkxXBYgYgxSpqKs
vVGVUq4WPUHsFS92f6wAisd5DEdrIYK/xi/n9oxdjiqnuJak9sts1UGYdfmU8K7YYNTUqXcUUQvR
UOYSsIqjScQoohUW3rtOFtd/mzf9QKUnfs/JGJYY2ueHu13mTMaznardBVENsD6UlygJdf+5eVWF
KQOmZt3bxMqbMt6aHPwuBzNmFjzKbe6kzkgXGv8iDUQm2dDXJ/e+rO3cVQLwKBO5TEjYi19dPB6G
J8eYktUjPz8fvyPIJsVSDPfzt61NllqboxIO+vlqyaa64awpupAY6E/StSkMijI+HK2Ib92yhfk6
9X2GD/8Wl05uPVSgr2WI5QgZY+hqgHPO0eLDEnlZ9rvzSdH/qJ1SA2t1krC3DZtnKxbhA1IRaXM5
QrATPTLnDP0HcETHLQdlgFeAyRlCkd/b0ZqC26hizhcDgf1fuD8aWaVYgM16U8aW2XsTECud/5zC
WdD1fZnELwFaeZ9MNcb05D7XqW5uQD/KAhiY7ovXWwihEPMzLkWFGXp+L4doXc9wHTXyEwgvS19D
O8RCYViH7dNa4/ECoioh0LDkcXqvoZW1ClSBrwF5QPwoOwR6sDtHWEDY0yv8eFXpucnlV7PhFMuY
3gCWfCCEMxt1oWRL1rCY5a3q1is8ownnV2N38aWcXQBTeDOGXd31YoLgVwxua2JE527LGc+yGz5l
WIWSiTbUuwd/L131j1wpepRfyeah6eVggv7ZuDdCMgKmloMXRwWb+qshu7Xgn0xWxA3LWzVjdpBa
AwnDxCwQNQ2+bEDkORwGM+ENlmgOGaj2FyYJdiDyd3qS1ouvJpbxe5asnfykbnz07gpI9WqC//EP
o0T/wOGe4qWK/9jty2kYyOc6LWfAUwXoF8JqWIB+Er0xBFZhVIBXEGRxK+bv0ZHP99+8xjUm206J
+XXIEA5IurXUfWngJHVHfrJ6uIbMVft6TgtOKgbmZHnjgJ14Neq/eJfVxXFG0j2Yi71iadWi6sef
hqDNzQeC4zdQkLD0veRX6EOOFc0MQHLIW4SBWSe97l0Hj16c/OzghotR7S2Wqi16ikhemiyJCgrL
P64jfPn6x/v4ue6ERlH1XtEJKswcxdGlCBTvygSAVdujN71BseFYHC1YqvWOOhhF/cBXZeDwyjk7
3963nIFMze482pa8SH/J7jt1k5YCgc82ggGPdcBPCzkL2QX+E756e7GdtOUy+xXGxILCh3nOkkxk
9hwOCucMvHzX3C5UkKDYd7KQ1vLhUF07Alp3STGQ3/XXPiPVlMQJzQ5zrcVA4MGQN1Kn5/TSb2fF
o2AnQfVxNbM8/NiHn3zDYgRkPgb6wZHFg2FtaTvd+hOaA9pRda+NwAZejngt1r+URtAAQZlGneVL
9CG69SUSm/CGQIXlquLx0duR7ol+qe3l8FZdGhzSSnkjT4l8kB40rjgCCasGJyBH7G6wjNPIxTzD
3CUQlP2n1E1rJ97QXkcQzTYJX2FebAxECwVF/U0y6Q8oX5PpmtzerA8pmcSfNFGir8vu33Grrev2
eEOigHQhmrS2Rhs+/GBokOMa8cN6J++CINraRq4/asD67UOPBFWddADHjwYEGeHhFVVw/SSMzN20
U2hrqhssMCHcabqWVahIe6+ciE4hKRcowVIoWwpVUIbI2yZvJGeKmV6jT/cVKGOaLoylVsf2u2GI
2kqmyQb1GyBfkPg7H9bKxMRgZDx9/B5DSNx3B7LIdKBw0MY3GnFqzqOMJmQWmfVF6raf6+QJPH6J
0tGUM8T4Yx+GILCc4pRDovO0vh9tdNpisYc4hHksLOIP1GmcKozl1UVG0bR4hPgws/1WARcYkR71
bQVqeMwb3rOx3JXykeilQYLCVCQn4FEWqUy9B/V5q5wHR6QzrZ60ijjhgtGJ3oc/VdCFSswGLRZu
2EpjTUIGhGQalhxXC3s3AQu9IBJ4yvbUvwBZXZnmRcTHIXa6ozK4qvUX7UJjNsQ+llN6JeFnPB7Y
r1QZT/GCpBociaOjc6r4bJWswtvqaEuRlLAKwhmTjUEM55fVk4p80wWQYZ0X4Zk+7I1DuTs7dDvW
VBETXQUPl6oTfQenTYIaa+2q27JlopYqU++wUyQ4RePeAjVo26n8Gl59Hp8H+fS7zrzemCXu2o3D
vi4cxXiRjp2cv5PSZWD6jQ7AI2d2d9F/2fW0z+SE53SqV0Wj9gqMvFXbrevajQZSDa04lDOBIMkK
/m8VN+AOszf6e+4TxE2zGAwwJIfy6ECokuLNi9WqRUuK3xm4h+Bo1tdYK0mahixlVS+nKp6AT178
7YWt8h1Nd/KdlhN5s2LDNRWIBQn5XDDIoCDig6ERPVjZ95igFsPjozhEJeyoLanNA/0JK47uHwHL
LOyHVNmEjbLwc3Ec36MyNq2jR/eD6bokvAQqhm9rKLSTuFNp+8RziTEqpSmnsej20HKkoKcmZ6JT
XiSQu8PkHU9WQTgv9TNlGBrsDucRzAJgO8prtQlQxsz5W/+JSCMdQ0OMo2ql7GX0Jb29ol5MpXRl
+ewrvPKnHCpXfTJ0LiUEDkgYypGnxS/PO8cUoHnYf79L4yaMmOsY7vunUMkGroEzkRdkwrZS/hmx
Bm5P0lyZmjjvuNOoavX1pj0z1rdLnQs9ncKTQx+O/IAwppsGeROJDPg1wu4fRuJexmONsx16PR0o
nWisw+PFGpveV+WZZkyPS0pxJyqSOXn2roCrGbsyyh2f2m9Ee29IgH36ruTWkYFoY294S+vb10Bl
f1U+rV/kyRqaRW4tonermsleJEtsyS3c14h+j1p4JRASpQckIWf/rVDWaWA3+CG3QHrqmtSIOEYA
dLQ/UAS7hCpaoQKTYzS6QN0TRpWwfUNijXwCfxjfHwqIgdJ3fAKentzJrp4OwUCDlzLvg1YTxOWZ
ocgjI02erU10zevfaOh2qDoAvPZFgN3fVBNB2eLBUQXqyQGZMBYW6pchOAevy+BBqOTuO8EhQQVy
Nut6JnPsWPcXMMQyZCjdCRs0Oy5/juTzpa3yA8/NP0EtDiO/B5rbHCqaT4kv7tZ5p9AGn+swtS0P
Gl/QLSBhRAsh5SUnCAVYucpEKMSY0gyBJ/eceuAWg9y2tfdVVXYVqMvCmcD4uAfAdUNULg068nxx
RiTTTmUsZu9CLksNHSW9nhPs9yhhft4/7TF3MypEtXJQJ69x6s3Vc4NbbG/M41fzzGWbYE8OvbED
7G/S2UwbwLm6Y4uo1WKfGviniHJiLSma5GtPKLGiiv7JuNTKWw1aY+SwX6rODmbD3a0OxGj10IrA
1TbldHpL0AXPKUIhGmje8uua8jDj0BdXBijx0oLKN4BhGRx1iG9glMFmuYTCYttY2FQJgbrjB+cn
XHIWqE49IoR0tanGws+hE42tXh1BGToWEklV2IpnqhQnLuiQsABLUcR/IYx2Rj+imcNTMkgkAndA
ZIRyFBPF/F0jNcXwBeiibRJMm3RNbfXYqC2XxbVpKjsI/YtUt04Bu1RnG3Keth/Ek3PAjB1e5Vmf
BTl736JcSQx5noe4kx5QAxiOA/YFGTAuJYmCyo70TGIRdToam1BkQzhbIY6hHxqcZJQV/RyLz7oe
iBdlX47GEOhymS/dWJpGXUx2ZctU+TGe4bSLdhYuHy8Iucv7N5qvfMe5JDtj8woEFrciTOUbsLyU
QGQpYIoRM1N/kIx4gte1Ydm1Op9zeYLiLz93oOVqYMGykzFDBLNL1Q979XPAjuzZ2t/GX+QoeWJi
XAhTki22K7sPR4p341+7ZoKUDBX2oyWPXyyH5S1EvHXn6JuljiYmzS7EM7egOlLp6S8XRnm2pSzG
/v9Fue+lAQlXThxax0leadtXxS9kikyp+DJqm+0n78ked/COjX6DiDtkW6unuLx2vCSfDIheBKr7
jbDZfewC2/G473PbzRUb7yVSWFQSEc9UssDwGdE1uZ/woFmZKviRjm5nkhij8BdsAC4qo3JmJfjW
9K8BgISXAPT76HuyNoDEKRXhwufkOANAKngW+HjQcwQsz0r0Vn6y6Coh+FBYdWp5RAHSx+nb94G8
QYuMwkufuFh6bCvjZTcniNcxMpZxb/YzuwYrDP363y+cANkH1/GAE4U7CiVF8L69aopwdh18FqMY
Edn47g1ietPtR0Ehzl2E2B2gho5thI80gHjxsrRPf0weN9/My3eYccLMhN/au7S3E0HDn2jjbrgQ
6GGZgfr5AdEdc/f5BhNSRu9ghhrlKVmyy8cMWYaEXinEjyvacNfDHzEVQECduYorv9H1uYAQkwTM
HWCjRalr/sbu9dSvLL66ChOB7Esy8F0OqYQbRwg88+nT37yyZK+0dNa2rHiO1EnaACR1j5nQUxAK
71nvT4zIgqO6UmC6SwpPwykJxI0OvCbpkwpXeC8Nmz7LJX9k5A9MFg3rDbq7cVaM72HjsG3w9kXy
iRd42kQiwbb0/Gfg9E/k9Mj8gfQo77fRczpYGTdHx5GYxvd0k2ezt7P1zEhzFLkZkFvILfS768PU
G/Rj2dW5vgNCAaBvOrwE99F3TN/vK+rca/Xj/N6wbK0y1SgDSeiStnqz8snVv+P1nX5GO9ZK+inC
B8wU+ERWp/zoQ4W86qjF3FUS6y8kcTsbIKShnERuKeNbyP2J3e9VcahvNdTI8gXXgurkBj3I8P+P
B+u/X5ezfw1+YyDq4lmqfVoJzAG6RFtKFQ3duRpWlJY+iHY6S37NWXBzoKVfKTQO2EFy6tMfq7Bu
rCTSJqMVTlIgPb7DaBK3ggxvoYiXB97DU+rWOg1BT3dolwuSDGcB0PCqaVdzGyu+4gxRw28BO+Hg
raBh/CM6QV+2+p2KfCgzKC5jNTZs0iWX/KLbt4MDTb2C2L+mXg1BNZxN8KlPZR9Ek8sGT/CzIxbO
5PbcT9Z8/ktLG0fuMcXZjrgRjJGx+gjUFj8/S4QtEbyxnaQDo9viGznodPbB45Y/QAJr/xQ9F0QR
e8rYUNdZbYaRD/BM97BwFUkJRLehgwcHQDGXvBg12AhLfo7QcoD+dtqL5Wir1IrK2wXXU5GG1vSg
pGXuxx+1pLiZEGyHbXlUgvodmQaESi2An1CcJz11Qo6wQrI0KTlBt0W/c94rAL5eJTlaAnk+lWbQ
rFKnVWWvUfZyHnkYVb4attJZZrn6VOowU63QdgpYFmmY6SP/JHPHjvObeTJslK2lGyeDS4+qYpZz
IdSIDq5MEUpM6Wtw+4u4YCTPfUNlqbTH4ouamJxnG9ZxO9PFS5Zf3T9NBK/xRXKM5om7GXUpU3vi
WOMPXT8UZB0JvEfiAytYIP+wBcjuXArg+KpHQpHpsWFSeiWLgN2eeFtOCDXPHdCSRgsiQkIM0j/W
aDXXJmxAZmR6J0qgnu5Q+ZrmBKJUoBnlDe/FtNHfpTm7WOEShs8dTJEdx5Uoxhe1Izdti6dhn0CW
79RRXZzEpaAqn6CrkUyLR9kvV/gZPdWsuDspmdrK4jrcq6Ae+ZiQseMTxNfXfocqwHbOtroJFw+X
UukVPd6tmHiiq7dIeJfFMvFDXS/f2JH9ABa9e1KbcyGHtS/yot2bnxvfI9nAETHdGR+K9uCUMGcw
egwVEd4ifumZtp0AC3DDEVV3Dirhj3Z0gjDiPuXOF6t2wytF7T9yhn0KnyzNuxWMuUH8FoATjM8a
IKggHus+4YGSAp4ofwC12iqchdt8nAKyr+G58/xa8FsqQt2KaHIUvzXMQIqWYpst7CTo1hQ+jqWa
QaTcmAM65PsT1mqcSC0UDuv3qJR21PZbFVkGVfd/eK4JjBlWpxQGEo59FnDadCKhJQZmh5iZ/jH1
VKjgWqdZZxRrMbWv6bHcsZp9vvNA24IRJJDDHlN6x7Pz59+TD8+mbU7H/WPnOvNbemlp6ZkutdyT
FMOChUREnWp+7rq/5R28AO0+GUnONQQBBZokSjTtTD0E+BmjTWW6VcdywDm/8PbasMJIfIW/tTao
gKVCn9umpf568BQrLLKtTYk0/CyM0ePMqbtEGdDp1ePMPAxJlHXv9KSzb56nCJoicbIQjYmDNMfA
JO5c0auvDpUR+MZsE7twrN69+1mMluLStk/nx+IDm/T6a/4bG+ndqo8yh8TApkB39KIPCGMpb/be
F7dCMdt3+nBtY8WTciBOMKZuZwVaIqqwVlPv+PElDau5woX1rlbCfuVfPoXqjPgTsD8xJzRTV90J
0pE/d3H5oJMV+ZMUpJ5UDS+iGxwj2AuRXz5UgMrsay6u+qd5orgvcaStg/QW6fACjPVzTNlQe7x8
smtViLNHRxDvH/HudbGD8b91QWQuOvhUgz0jO6J2g2bkynPPbELOJO4RiTR4x7yDBCSNjKumf+Uy
QO29SD56Lo+LGKjxSCmBR6Hi9MQ/oUm17kram6PC0MNre2XhNGvz4k4PvNdtH3vGLTDziYhQiE0T
jZ/b2oXjm9N9Wi/d/zDdBB7cFNUObjJaPplM18Eyu7t3aSUkCJ6ZOaGCZs05GMI1nqgjMZTjqIpQ
Bsk3O+GwVa3CO2cMvsXryZqcYHTrM44EVXrDI3aQuxn6X/ZE8vkOFbHoZ7ByjIP3BT2X9+1P72h8
lZ1YZSYxJqoqg67EHgro237D40BTUfdx7ct6dJBsPgFQQ8Bst9uWZBXXmBvX3fFhDbFkV63wzlat
iTkaTXzCzvqeRf5axo3qH7de+dRTx4XfnQxrzD8CJs4/WBZHWegmjRPbl99rQVF6/HKbsucVJXTu
mUU1HqVSfgjomASY2rOVErSkrE+kydQhF1GBUxKUTUjmV3nhZJM2K5j/Osk8KyPtW6q52pBwMeao
TdGlt9P9GV+dk+9YsVUq5aC8llFd1o3VyhkpihGMPOTiElaxatmf2YKVbDxtWSx4qrZjhQiOA9xe
DYLx7BkTT5VaFaMWUQ4dN0Ap/OlMc03fkBc/R1BmaK3uLIQJvKG/xYO4PrqYi+HOj3mvT85Te3aK
f62S3ZhCx5ZNbXbbg7FBaZPeZw9UuUx1xvL7wVfKzRNfBG32SAimqNa+xN4L6K7Z1K8r0VYxMBSV
WNlaaFRyA2VfWVbL+LrpxQiJL7f5UPcpoaA9M93Wi7u7fL+NSxS+5LzvL54Lox59x8EeMBOlAOQI
zRCY8dINxS9aBj6uuvtEfJR8M8gvZ1Qm/aKoPkabqZ31910gnqhiipegEyMOOC53fUSwGJLGr/m4
Nlp3eM0LrVboBPQmN7Mwjx1akmIl8s8uJprtGH/sPOKgVntrFdNQP99zWRFjC3OmLQm46JAPo5Ny
l3c21q1RocNyTvh7SzOfMl/pejDdqY5EvBwnd1J0d+BocM6djr9sB0ptDmSpKtoCvy/nYAI4GO+u
ANWBptZ0d9Zu6quuQIM5PDJ9WfRBvH4zIu01dqX11d6eEOAv/NBvWZcC6IbwLhhlBauKJtDLFOXA
Il+Xl4UoyOpJE9b8eEjGgwdv7ELQAiGhdY/gV3vH5nTbx3MZ3Hr1ycgb8/V048adSYoQLhEItPaC
LhRctz8+ij/gSbt22V4pI5GdYXwlbLuhzNzUyN8DE0hNzyTFEcuGtugOqUQEUjkX5NXrJemeirlf
T/9OGH8FxygECTunCQw58+tnNpesiO9Xm8sH/49/XleLKk48AcHtzeSfpH9Qi+s0SyKDf/jDz0Bh
Y2MKKUsg4s7Wlvz++vsTKkc66lf6ISHKPs3tcQskskXxDkl4PtG16NEKjxsdix5HY0nMyBOuuVcf
Cwhwpe2egoNJtwsQWc9J64nMvpcq5bmmt3Lgcw3s4BjzNXMPoC2QOhjkl8FX7rlqdos0zmBIYOM9
pQOcmulbKdiS8CvulSVA4AcHPJ8lOkymmqazE+f8AQR4XRyb+9yagzPlCFn/Nduk02uIJigAm6SQ
L1mP2vdJfmto9ES56NFRfjhmqXjmZxDNttVOOdZpLnlcTtrNqlb3H1S1uaE9puPz9mxZEu6RI++X
ygzZBpTMiGbaWab4PPTfmbchJRQwxANBy2OXpxzXkEn55e/PeAOuu++5GRrG0b8dIJxfEORNHu9C
f4JrjCdRiIXnBGzGghXoH6VBfuIF/9cEusnkMj1EagqE4XSDdNl6wZVanyhxz2BcSJQjCIPpl24A
Nhpp0QfVS7kmDzVqOzLf7guVoiqTy9cvMjz1MlZmeAxUmEiMv7QG9cAtaLbPOGjeRPwDZbJDVI0N
jeibyXccwm4EBg7Hwl1Je1BlagGFlTi+C/VLgEbe75+FpG06qVojZMWQzTZgMPhxS6S/uYxcSmZ/
nSpDgi3GNvMpa5GEZbodEw8L4jWjGQZyodQYdcs2kLcqcsuFivlOzJMpc52oUIDtJ7IWJ/HZUtkk
U9Z4YDB+XVu7yrIhzXaISH43hEBWHlFim+hK2kEpQ1hNPpMgIYfECBJ91NXkxdnRYQ7imPkpc8FR
KzQQug+sOlUcmK1JOMDUl7OWo18ALyQGd2Ilg1xNqSxhPNm3H3wM+kjZxugHWUz2/H9+UZvRL4T4
gQP+JdeYW+NHjs8UykVM+BpRWFteKGj8KUwTleTOu2iFFTZInFNj1sHJII//xG2FKW0SS0t3jjcw
wyI4emmujAuO/OkEtLnf6lb7xNG/eorRjeYANAuhSUJR93nu8HYUpPVKz+93Sqad1DSN3xAZE+Uz
qxbh0f9GZaVhgq6x6A2JpF4tmPsUVR9Fy0T6u7+h2Zd4yzPHN3oZOO8iNyRnNF0olrI167nRFcVj
hz3Kehws+OzXJTIAV9nXGKN+VFwvrpCZgAk5fBC3BL5q4RyUt8NqYcn3ubAEo2PP4A24VmwTY0b4
nrM/JoFNh3f5jerFJrz2SR036iFE3qDQs01GOVIrcKHJlruqdoL2pZA95KDhjmJ/u1iLC/dsgcpU
rs+8qrYgaLJaTag9aOMqw35xmN1eap/1YbMfuAKdibj3r5iAyYXCuMjvadWRk3LVdbUv7S1r7TSq
Mty4bCIb5e2qHfHnCSV7NcrtrgrJ5VMJNh6ICqvPO+ybxcdHN5uTkcRd2zWmh+H4WEtKuY5oS9Oa
b1Kug+vVy8u3wWKKMXmRUWoqS+w5Y/lDTX1TK/ELZsbhw5d2kNKY6LAiI8jOP6CXMhvXQ2NE3CNh
KmtxCxaGMqpIjWNj/1ZnDiWlk54ftXsFhpM4hA9A/oJeLSmGWft3pLIiLNimFeWohTG+A4UredLj
tML53pEPaJHrMBvZrRyq/D4kWOD9TEzxisXhMIigA510UJAbjDFtlIuokYAFdnhJQD+C6wFRL0LG
aHrG+7RLzX2O7jBlH38xM0T6Qxq5pg2L9GLMgcPyjPACssmP6P6sjeo3VQOKT/aSaHn6Z88S+uYf
R1il4pqRcKrRSi0ZDNHmOGxXu3VCh3bv97guTSJLBjABdOkvlQlidiNGBq3XvpwX4NrwRQFY4AU2
M1KLH50CJlYCdVIbo1mzKxN9bag6HsMA02rjgjSoGw4Q+EkD0BrnwN7VUR25C7N91YmwOF9b5ORA
y6gvAp/bDxjklSbjrFPa+H9qtaDBS452Zzi8UN0g/gQ/eJJRsAfD9MguFSJNcP9W0FzmEKz78+xc
vpfZkQmN51tBVt5X+7oHU0r1T5Six++6WqNHLnynvvisRUK7xfa72uoA4bUTzDXFXiaunP74I+Ml
Pd5gMPFZQcL0O4fw1XZTMgHSUjDqooAPYp70eRDEM6g5BXIvKYdRkxhgUYiPwOvP5f3hD4b9fiOS
tl4npijg0w5N4sCJsGjnND/b/6ObD/Hz1AlFI2DWPSmEja+X6/I3LdGplH82f8QDOiBFmxPKR4wW
WZP9VL7mg3RiFUq7E7fmFD0IalkouPqPqh1PvjrmLJKNYI2vIbf2DoaXp/ff3Q7MGAnMGxGD4+bG
fFHxCiLmqaH1mefEEWSiX1MErrrp+25g90NNRnZjjHAGeKCQ6BBX6COiOnfw573kH8U9r2j/iPLu
/LlmVxt3SMZ/fVRkg9HwdARQy9Ujx81hdW7gVZ/+7IShZJFd/FENg/gbKzfIak3qyEyutzm2jWQL
bvw7PubBiCyzSBoVtLMj0rxlsYOziOK/K5fUXb4FzgRtWHdl68lYAWOFJhTdANboNUKbzxWLLyFm
SyhsFemvGkmN6byAlUzAywGU3G+F6SYv0u/RVkmq6/SeA43oETjlsQw+o652C/oJMmKRvDLw5L2h
SurlTSam0aCZAaQlrrhDP//L8x4tCONdiFLAnItaTYAWq9gNsUyPgFl9yu4D2bpjOqz/2d+LhaED
3Lt3ecNe4QUt0lv0OLUX/a4wZS/dZfXEQyNBvpReMqc23HDS6H/LlGPd5qRpJBx1eIsy4toh/xJY
Av6RijmTHX/km6SPKj+1ajhdlTUCz4sXInX+syrG2iY9yU5HMe1snpJgOyq83RsmPpeaoD3Jn4gJ
qWtJDjW7cnXTfGoetGLluIS3BWjFQvplyroM6eB8bxfc0jIFd31uGfToYD88PXm+5rE0XtDoT9hP
Zka1Ai6HHVeAt80VtmSuqC7pNlBzh3rf7hHXCUUOhEovoH3rVUYhgAfwj76f2x54qijRSSTG8QOJ
FggTfWNqQXoPc07n+BvA1d58zLUZGUEuILBYP8e5fMr+gf5lcxtADmLl4HKnWyTcxOM3Zlke+09F
+BLmQxbeOczIcPym1IN/tFN2+adtMRhDFrjbHnc/WttZRKwtUz6cD3D3WvEZawTITdRpS8AgmLPc
UEDkCwctH3h0Dcxl2OcaGzeXRcY+bcUJGbT4hl/IRjE0ZSwX1QFbLAUu0YWyXtAgkOY6gEQZ/jJH
ZKPo6e4+dYgmFYt9eAioDRGi5tgp5D5NhGUchs3l7v9Sw1uIPWVFbm2nr5ZxNqzz7x+tG30NDa2i
AoCYvTzoNCidbWQpLzHWqxA0xSYsAyK+zFNvip94U/KpD+yoQnDyJX7LMbJPAK2xQOQb8KuRePZx
HstX40ifHIiNI5yAanz7CYCYseYdeXSdrfz5B3FjsaB1DETCX7z9K/479Ox3ufsiq8zE5WKu2T+M
xwOhUKwnJZgEd0J4CEU0xzAxfhV/tFKK3DhBwBdqiyy02X9qsrTuMGJaMKfCqLSlUZtqdosjapzs
UFiWTrkJIyZjhCqZyPw4as7BY9ap/47T2ZMk4BZmuSIkNYaE1ZMnviEygPDXUwRmEvl7HDKfDOvZ
3o8M9LGYBmXSPkUh2g1HgTixyjdXqASkgdUL6eyPdKl5ib5TPIV91BLtIiL3fIqu1ozDfBfg7nk7
Cnle+5tF74JeZ4RzAjIGPdCpfe1+iTCLcP34Mr3i3QkuV5O5tX7ugXrhGEA6ZJ8qborJsD6DtcJi
mKnqg44PZic1fKH7B0bqlne1r3dB2yHJ2Ge5xZqjRmOk5Lx7O/F0PYzGPzIsb0kUDZ36CYcG/YfX
2hj1+wy8Nyo1wZB5KXAHUOf+85cIC1A4/AbxgSw3Zcc0qcDUbW445guKWZxEKheoTABTBmMGWuLx
0OcLsKMWY9QD0B0Qus6Vs8B4NRdOI1KKUylR+uv05pMx/5v2S6X03KnfOrxxrfNx45veSDbOOpLy
lk1h6gwCfqdDBxFZ6RT7fRWJ7QWCR7EtUPQap2f7YLjoWssbVlf01npckB+rwVbO9agEwLdBq/0q
QfQ4ohxssC1r/itCb/f4F+RLsaopxopgri1FIxahQye6/0Vf2i62TOz2kj6ufmhCrxUN5TbmRTya
fSkgc3zKMg+zM5OOSG+cMZ9u5CzRs+38Sh0oDBTvUJJ2+50C4lCW5tXztP7hi+rLL/6oBikTl0bk
RHo4siz+usEMbdw0ShfCFHXuUZ4XYPH493Oe72/wHEVQOP1JB+tr8/h7Pz0ACxS2ix9bs227UzEC
ZcUd3Lrme0Fdr+FDQOggAkNPwoJzc5TvB+po8hRiK/ovSakeabJSa/8d6cKZH1FlhqtZPZ5uAN9h
0MmBnpQI5hLs9VuwUW20KZpvii0gmr6Jv61nv46c0mKmOpo4t/JcIgvkvbMyCyprmrOL/IhElgzo
0VrwJgWHNGVwchE+PS02GVpV8+efDIVzqP4vc0RCG50CNYVgDqeEJhat0RqwgIqkaSBTSaSXTDkM
EA5sSxxj5sXHxsZNWtlBUokfJdNJM970LQAY9PkFK38G5nzdMDQXtMbPxEeY1wXJxuNPjYWW+CTQ
6s8WU9BIwLzLbjTBqR7dMzVvey6OU39qGT4zimVABTbtEUSp9XfxCIWyDD0U9isnHvB1C6EM9a4l
AjkMyFMZHyW12KpO0z0e/DFpU9Vvp680gDIzDv8UqOnLQeqr9IJ2zfMlkTiSwCj+qTw2D5j7hJ1a
SAFgdhS9CRKPw5xg1+QIKy+9eS2H3/L0fi1nzmN5bX3HamZP1ptfaP2hK8Xojl/ZkuMUrEjIT5yA
I8JB0On+ph6vicZWon8cVDKt+qURFeYdvLHKL23wlguhrQdftiP1jWUtb7Dp36bY3alLyZ5k5VNL
OI2TXvsogRvNgQjJUiObiN5bRDd4XvkmUhKCxCHKnTCSVsqcXkrwlLKNdM5OQCdkQftuHnueqqMu
xGSe9xPzl9Xk60zeRi2XtHxJfS09Tcq32IHI1T4asrXBbfpRWzkwQtRBBggghaU+AS2imLqLatc/
l62Yi977h7pUzikupHVJpNhJBvFcpGpX+nd/oC3GyzgqViX4euFKxPheRT4vwBxAzXot7SDJVO2L
8G/ymSUPh2rpUOWi+FnO+q7BYqdu1TkjlykphysTq2xfvoCiaoGfpfDKihAIl14epdq0fQPZOlRX
wbk/rM6u74PWE3j2pqwsB3XpwZHdemYTgz7oRDA/eGVjrOdzZa9he576fKdbnxeTxtgaxL3rEXp9
XuuAz7AAWa0jvOpkVurUx1GOAX6z8YyoRqCp5dCKYpVG+0KI2uLOTGFFl5vRsfMLzlgzTpyx7f+G
W3lpoTaPiW/Tf1k17J8v92wJdHHZIh1ADQVbsdM1jsOL04s0xVAIv7A5TAN4AlJPw2jJ0pM9nfRk
X5Hm6CPbf1HVbJhz7wSzXE8UGTcyGaeAwk/pQQyaeQ84dQKjAhlJgw83k2Gg7PDhcOdU19S2Q2WD
aNwApq1k7EE5grLyJyTrhoSBWHuwAqm/FmnGnC1fUXtTdLdxsUcTcwkvOv/F/xG/4Rq45b/5SdDM
vNY1ttxwwZswATik0iubQUmzakpmRxxM8DusPisUV+iFsgODPgE3tSrEp5atWvvGFFeLTwgMUGDN
frKAoRQNyLEJwrJD02SV93ff7RLgoQQ40NeUTf81s3XL4sm/cPe0HxC6FKUNrZjQcQb/lvtPK93N
u3iBAwrrzpdTw+ulEPJTEKKp8Kcoywc0atQh6ag7nnYqs4Ffbv2ye7K+fbM8htDA8K5RjewTI5ja
1MBD+hZRLmf8+Zo+RBr1GslgnjCHAuWmFRJYYSkGCVQnD3oVM5FHu1Tn4+ubEwz5TP8T20TfiHbs
a8mJiBIUq35rChAixVMLnNAATyQCjbLEFglG0qz1vE5EFOdLsa0WJSMlsXPVlR1/vccunqc3tJCT
qq94p5FhhSj0d7QstOH9BPbVlzKrQUr4rVWn2RKSCCewuAMON1oVF9BgxQWpeTQvd7wGzgFPl/4z
+Q+g8itgYXOyi0ifrOZm4V45tkzZOzWkXXFARdAab8p+Jh3qdigROPZY9u50IodAHTgBkbmbwH8i
oHiCeomWs0yGT0oEYQa5WpX+o2kU0G+5ja+KtLIK5w25v74mwEcK63r4kKHq6FuCpSN9Y61VaXPF
eyNbX+Kx3HxUjnzQKEKtmrOsMTnwDn9GFSvkaHxB9XMuMmnCLXJxI+Xomgi8AVWNz460PjDm/s/E
G3htNlS/+TYAXAx4qSYDIM+/iFfgNYAsoHapHf/vvnPupSkBvwZNLt53kzJW/7TxKb7rsJt7wYlY
9D/5Zb3ujvNOWKnUzavoP5TSKDE8E6NTLgtOsCXr1JNgIQ7toCAHx/frpzbugKmIYReFn4r2IUpQ
Iudij8EmHs/gRkllhUmTM2aoih7p6EJSvjxtwujYBLwBI3mznPnDgxpKprQC5/xurWaxT/9n8nCm
M7PQczax9H1BrP2DXe3GSd9OGHE9MFEBoJ6Tg7fW0dNm7mjymNVh5RBbfxrDVYDHXNzKPrByGud0
yiL7I+LeGHf1EbVLQEVuFMGuttGFgR2/fcQiUjp0R7FaUILSzG8YFrLVnc8+FOsymI1FdCZ/jUbq
Pykxv4albWa2zQKNw1Fdk5NtYQWi2ezHNpkxNRB0EWS6AnnAEsmPTOJto0NBKOwrJDqNC7/wL1GJ
I6lQ1lOpjBnWINtHUfUDfheqt3cujAApw3ffgfqMoYyggk0RficoCYnwc+H/50N/E6LoyOKDddDq
6Mh5D2D/R/OHV3By8UgjbHbaAvf+47BygQhasKqRZYd8JdZqqdT8BR2QAlBd7UynB7+ssZoqWR6L
KqFVqe4AH2NbGObvoNDOYz0YZ0bj5t1hC6vAdoT3MpwVEuquC3RKZ6ZKJ+vuBF1XDE5MRn4T778J
V8QU9NluSySzBjM7Hqa1aX7UN0tbHCDKs+bKNJHgt5X+0txP9UJmpTVQeSHL3IoHbDHt/Dr7zNgU
wAit/tmr8C2Vt++3BWcJejrjN1w1shzRP2OHALcLKJiOWPF1nG/45cnkZHu1JChkFr732RTLXtKH
Kw6XHf6ekb8Fic9tGdOKbVYwx7uJAFUjhS1Nw+YQBg2qgX0TaANI8yiBa8p2kYadHnjeg8JD4aOB
qqbsnmXUaLXT6NoA7105k9+ficFpTEYPFjVqIR+1EIVdXOQN+e7LYOIh+9pO3lEdvfTYnX1WSDkS
YNa+V4y26K1um9vAgmQCrnV9vuKCxQ46pmde7JO8ZsdBuXNHcq6tBLj3Zx0sAMFW6OQ8ogJKclBQ
/RppkTTJFvdfxTKYIphPPbrH6z389nLXYnL5GRDEmRHMfD/uMQ6x30ZLFvPlzS+ZWHaQu6HY5orc
H/JYysP5GDjD1sqbBaDEsSlsRm0SdEJMIqyzLyLJqgafw5F8T9lK3KOMTssv+k0ylDNgnLdOBDrG
CWB/Vw/FQCG9jbAc7DkQRRReb/Vt0OfPIhURe7xHbyLejuQtADCPjNOuFKGalwcq8ZhB8yiEHrI6
jlygT4iYBYOQh0xN4fJfuDFYzb477aMTGYLfWpW8ElkjFS5JXRDkFAfsWHhOXb/c2wzST4a7OQ6E
hoepbpmKkdZMXxtrQmFcRanJZrjmOSo+Iq073R6kZW8OeBMtxHVR85O/KxjW6kOW9mzlFG93zRyK
66jDJ4hPwHeXwoYIwJ3r+szZMiRAOBQ/lYFCsyH9ImHCUJq35v2kkfZ94/Tpl8J1dcIFnmFYlQA9
nmvKf4LfH492O0mIJBner/eqQZErLvn4aHRAq4ETRm/EhfGM1lU8WM62OSF68M2N0Y6w1d9FYKfj
Y3sQ9jG0TE/6IS/nYiiEXoeDdNiIg9g7ilEW0yQQpPoGdzeRTm3wZhzL2EMnsTtWEVjheLtnfyLo
qHwUXwWpJmp4HGJfd1tlbjXGLmc+KNb01iwN0r8bRfRUKdp98ojq0semQL8JeTVF30f5k8EUPQlv
URPZbyAdHUX7zcxNbFaRcbnE1P/OIFnWCjxBzISTrmBLz4VDGIGv70wY5dF6ZtioodCYTh/Vu9eC
oO2E4hpMjDb4gHiU+aTl5iuCnULlr7rIEg13H+PnJRoFBKN3jn9P7VFJZJfybUJ6vRwJRkgtRSP0
tN1525mZfSP9Bq3GhQR8wuedONsXYxB5WNfFoyj/BeWW8vmkjncJGm0RDf2xLYoPy3lgStNd7ZLH
Qzm6DclgVx+LZivyxyy/DgkIGDuAQybpTf1ox0Pr9fa6YSjf6xG8ZYJGH2XBrhiNaBY61YLFpWZi
3/21cz4bGeKGAeBOcpZIAFwXcDKe0sE7WUVlzdUQTH79Vc9U0nMxUbsCBxaBmftYaJXGKrVVFeFV
LEc1ayFRRK+5MFp8XF0Bjx6FzZFQaioHPEHw3HgLhteMH5AMk+Y5CnM+W5XBDPJZcCQL5eYrwIMl
89ZS9dKE1TePPFeHBWNzQR6/WI45Qh3BtVgGnR41Y5Pjc/nE2ux8pBoxPGFZGiP4agRTFZjAMZcq
02gnv++OuAVbUl7mHKSN1kLeY2C0KQWOoLI9Iz3AeJo5IKmDWnE3/2/v5izERzga6/ee4Nx2VESe
0Jw1FvDVtP/jDYzCfAGZghoPk2k0ERHSDIdYUFhSb+cX5kyFdLua49CV397sJuPRLrrznEXcEl7H
LPxzfT0zC8zpqBVYSep4ucVACDY8pAWnEvg54rrA5862PLkqqxyYIecaYd6NH/7SI67eyvoUJaoQ
qdCv0G9lq7kG75+gahjRac3qPYOgBoM51X09Ay8E0HyQ9G06pBqle7YUminFMadiUDwyPhVQMxqt
LdwyoIX9SW1+CmAz4UFo+jY/4fUfvyFXl0j7KmS67lnNid4ohaAsBDWbxBnruKywgjxsXIpZIfsh
PjgidLnpD2wgeVblrIPPnIQbmkKDEZ7T9CLTBzPzvwNjDix8HimSD8hEEwMXu/FJGJtkYkp53dWv
kGTP6SYz6S9kXwOKWiLE6QeO2RSbaZxyribJy82NgTNWgmcmcdD6z6h9GzE5MFhuAQoKwZiszNT3
/NvoD+2Mo5lPmY9RF7VgUGFbn4afB7Ca6bcg+QZHxn7MdzzKt1s17rXzhnvKooe7ipSUoR8TCD4A
KFU45XGDMMTascIqidpPXuIzfrI2fMSr5de8UqH0tnbsJI/LHrCgJbvQFBurUOgEZqOu9MA5Ieah
Kup4YCP5pIE+2A1ggfX1LAW+qp8FKDHYT7t99/SM5US7Egzb41UphPqT+WCfsmjTCJXj/61NJfkS
CaDTK7CJpVAv9BeLWUJGwjtYmUMmJqrOhdww87L9gckla/6DIybiPftlYWkhifn5D4vNYM5c7yw6
MehbkihpVHUqw9yxKWUrUuKa6KpSxlt/chOB+fhwZkq07LHDlEn+SxeUTqsNmYP+2pSnQ5Vlq+ig
+Q25s6Rasn4L1BDlYq7yUReihVsKm5ijM857FtKR0wWJPISEZnECr9omFZjbR7NyVO2zMuvaUrqh
u7v97E60xJafQpjHfbww3kgH7X/X42Aa/i0bJxujSPWQ6+skU1LXhKpzty0I4K3V1N/L0O45BM5g
TKjaGepgYdp4fAuypWUdTsJc7g/bdIPUskEQWFgd1BsxWW95Kv9QRRTdR3M+2/rB1M/p2o2IBsU1
b+td/jKosThec0gYb+z0na8FlcJB/Vl1v2k13SqQLFzS1NInk43yl1UpLq7b1KBUgqLYUyZ4oQud
SwDK1zJphth2O7HK5KykqxdMPzIFNjUTRL9tpy/gGihlAFnA8N+zo1UvFvT7wRk/rGR2aHvcDuwM
VE4hWsptYzE8ov0PLVYArzZ9TEx4lcZ4JS8ji188leYnCMi1R88ciEZ1Bneqm4G7fUwfGP6lcSrv
d3cJQJgQcthZXxmDVEX/fndgzDxKC2aj+X3VHC7TPJxND3vVA1E5WDjCpybs+iXdIPBDwXnCkkhQ
70baVt2orBfcpuhV+k2xdrJn0pcVTq8/0YjMfuH4SrOv0cmmQYwL0NuJvpf2PYOWU3tuT3sKJl/5
Ft4IAbmfpDCygTP984uWEKaKWPgYM4svlcBVgKFeJfEPitFHS1DljIin4ow1YhnW5e3sic5DpviZ
EjDcYS3pndS3dw06n9Yt4l993R5+RGbYXdxA8Hp3vyKPr/rKlvBkbM7572CjLAUFd1FBOVrVvBlc
ozgkrXIguXum32ON5HJMPpfUeD0sJ3kATYnW1s08zNIp9Fx0hqp7D/HEOj3P8UGVvAgVCqJdbk9e
bBKPltx3JRIX6IHjSyvzwcSlCnKT2VjX7QILzJU0SXmdtVcMHqphrDgv5YTKYWpEUIcdPaqypRa4
pDccyNVsbMEOJKKmbiWgLWTe2QLE2l8eqIhBed6//vIKj7FhGQsZrTnqitBH7dneZsa5SeWpIa2Z
LUw4RCadmbYJpvAlJSLQBMkXHjq7Mo91/ebi1ciabj2UgfeKZZUfSjQ0Xfl2BlDoB/gc2Qpd4bcs
Akc9RSqCCc6+6pJYAAGdbLRnVoCV9dvtFWjbJ8ZpUOBh/Obe7tuikejaquQ7IkpRcYtXwze03vMR
IpY+N9vJsIVZcKHCsr+C1h4YRvQzPGbUsuHENfBcdOgvKVtNMkXIH3cABbDoc2rUY4RKKO6tlkPY
C1u2CtkpT1333OY9STAvjA8cR+DJlt/q5xhgGjMzYsYejvKJtV5ac4QjCYzI5YsXq2uC8pADY9J2
380JQq/5sh35fNgkP7zsgk5K/mtC51rslHqAQb5MPcA8IeMi2KMBYi3xEukHsbSgeCyEE9IjGceR
XPJhuOSrrLQk0nl6WMhoH7nYYTu58NC1dtic8hD9kPdKTsKHWsL86LIB6qpIyDz+dARUNRTJuWNW
ZK1l9t/lIVaYCffjAmDIjqB4YzXBsQbMK1+cvpPYmT2MVXRIH4Eb04KvUZoa1YuWv6iwsYVoGMTU
w0lEjbuNi7F8QOOBgtka2eYzqxb/XtwFSwTb0Yb/RSL9Lb4ADMJ/4DtQRSYvKfQpFMMkTtOc+vjH
QLNW3uM8Ni9OMN4DFm7QwYQi8VB5fMz6Zq54jLZGPbQ0n8svPcQSpxIYBWN+PSPSPMZtrdP9cmAQ
EnhFLvC5Q17Cp09Dv+bd1NYk+QBt8/np/yyGVhXlGfYbEi4bkW9Q/ktbQ5TRh8gJT4LktAZ0Yp1S
dHQBwjhy7ufHNiM0fhsvveIxCowyTslZeYIp+8sVbEea6OL5s5CNzh8YTnap1EXDhPA4hSL8R6aJ
Hp+A4hRIV9qz0NuAEW4+nAxFvSrRoLMc9a8PlmHIqMSdCKVTAUhFLtJEVPuNQXxTeJ7QksnAwdj9
NYloMueb9juXAJR7/kookSPezc+B4klqLfuiAfCMAqg4hPjY+RiGZCPC88co91Z9s9MsKV5GZQvf
KEGQCFyyAfEBIx9jaHw8YXsF7bn5EKZJOaPdROd+r6wBC7eH2cGIn/yz1NNO8zEknBJWm5Z6folM
fZ31yQtS5u/YL6c87/bbwsMih/jtDj4mcH7fCCNt4I1+ykVrOLY/CwdUCHaZaFblINJNto/adXTR
pg3hssSOelJCHxkgaxci+JAce51pyzki6in+aapSxS92m37KBYW/FdYF1yJq/nenExj0yH6HEkF2
CUFZ8KGX6Z9KvZ2Dcn7P1eDZbylPK1tB0b3qT6YX/p7zjS5muNzOZv2hLPWjnrjTVLv8O1Ogu839
OPKs+LYaPnpU8GTwtWrufspD/KDeZg2ABWSkb9O5QmTB/giJgl5R9mFkNYQ4VeXdo/sQREatwDW2
46yCnW9f7xk+b9KbgCvwXsXykJmqEeL3T2ALXCHppLJwuZUZ5i/rWw3SKJTnAsGVk3ofinslnsf3
9H5sB5oQxH3tvW5H+lF4zbciWMFhB4hoYy6287UhU/c6pBJmtwOJXNjCrAKyhbMfibSy5THeVQ6u
XKdLBNhi2CGpmRulzfPM4+f0k5EyUJ25q3RuRQ85wjzCR6zlGCKSD2TpsEN2g5KAeS20TtVPDsAL
ij+ylJucvo8cPh7XNNtFjNBZpEoosG+A1iyTymNPtbdniJ4NSoBK7mOra23wzApUp/lqpXjosvPm
TKQnEFxJ/eNc74VF3qPtCNpjzt6eTaiyH/9py7PXhgpo7Z10i1sews1C2WimAcVZjZaSNCFYOFy9
xu0o+7JDc9W/w1zsjGGzhBP6RpfvmPoTQGoM33CDkpKynV6C2c15FAaB3lg2L8jCn26f+pZGjyBj
wJ8RQ2K5poqmfdpZjgPfG7JbOh9Fr26hmWysID5eNJ+gMv5uaH6yo2TtT3Fi5GCbw7ebbfAjQyT+
kho/BQ2FCS1jBp7RhWXO//SIfngw0gZat5vIaDmzwQ4cABqfP9KjQ0zCyAweBwSR+B8f31amjGqK
KmF2pejjnyeJNzCHl8vtm7tHXAStbcUJd6sylmw0Ii/GQej8OzgtDlSkohnhBKu0JfqJg61MYzwE
xkZ9MnDU7GgArI3zEy30WxUD5OYdQHyWfKRtx+vVgpVS2MiQlqzuAcWMIZI+c3rPZl+xu/H5SHc0
Ke9Q+GVZ6vUfelp15As/Vc6uvc3SuN9VcEDweDNaTzXNqD/BBqiMCXToer7NePEp4dp7KzU30Lk0
LPdqzxoB+vAZkO6iZx4rAuymRPaOM09kZUWPueVEZOaqrIB55S9Dnue0VdDNC8OYvE2h7gBn3W1Y
rrV9OPRWjYBTZEyoBA87WZ2q3wfQXe0j6I9Ba322yBfgq6oU0CUJZ8ON0MAC/qvtdEI+my4YOPp+
Gqee94Z7p36mrDRe5F9dPH9lwjMnaFn3Gi2TEzI1ICe0lQmXnektKEOkD5RDxqK5IsIzVewum572
duKot5cI6coU5TtjPwOvtwiKWd1TFy8fa43j9CPCHbiTEi+p0klrsbA2i+GZcbE+WeMjgMzTOmgN
OYWjzlR/hL1x/1EwQ2BysqpH94xZvuTWBQ4C0Hdjzej3ifD37KqvYeghma9yRa6xvZEREuCAptq6
EnPTfhkUD429YQn1tsvS6rKtLxqeuvHL2CHSBa8oKYHfT5/9VF7yGxFeLu/8X8fDCeVUAzY3TFvh
wOBeUATKPnzejCOPcmlfcOPdKHH9Y7cNLaRQQUIIxmQBr9+wBbzlx2pG8AdcDbuXpAPku+LmWeGx
HHLHEmSNLnMxZ6Ek7x+K6kbH1RVclVQksG1oTu5Ayv6lGyqNOR06uvIe7WZIIyD9v5bZjFHTogog
MjClgKEJvp9yld9c5+v8U7JzMy/oYGg6I6T+VOaE+fX9i9FHIn3rbKe0uHHVnIL3LvP+IKvTGG41
lef1eagzkve5VlXTv1YWjHwCR+gchyNQpExDEtPWJ91oHAfV5EKm6/AdCS4ynXis1LFHoVSaIjxQ
xnCMHkcDjXkUu/CRJEohAW4f1qQ5c7sL6pXYhju68Uh3yOXCBoTq6IUweMwa0h0wVwx4IyMemWAC
BVUbPd0z/PTumfvwXfpBfNJBgvSfgg3RUXYkilRhkIv9i4tMSVGHUUiM2xlaaC0T7AqD6R4KrNOR
9Vmce4JLNC4siOlqb7h7jZcqkN2g2/HdCR/Qw5PI7nJbXzpkhtMgjiYoF6EJZ3GL0K0uTY5jeI6r
sGaL639PqFmhkVt/Tm2YrzFVemkfIm4JvVwApR4DMLybSZ7hX9vlbTydVY1gn3Sft2IRlW8E/Sa5
y9SjjcJk+zMQEhNZVZ3RzhA+5TERzbi6Wgkcv/n69LYxcQStiSHKD8lTXdbYxxapOg3agNlt5351
Exw2+szisjbdBcYlLwKBs5UurBaj2O/+5VAg4YAOpFLDEINzs/lZ3eVTPs7P3Cqqfj6tK3JCHv69
kgJ42yPuy6ohrMhRXPNPdr9qbzHNxVpwP4cNsA6APCuRgKLVtYZqv7BklzUmMqRp6oikIYvfilrD
SIjD2EhET6QCLuUltBMob3BjOmnPtcPkqpJosi6w1tJzait3EWViRgUs+kTnoq5H4K6er57Wcwi+
zUUc6x5pCOBpd9eiR57HeHlcWHCBzGOw14galq54to1IJ6WxK2k7SabiMuIWHXW7hMOoeJAkLtkZ
/nQjsxlZMOib72RH0Ag5UGeSJZgHM+mxIKACF6+k6s1kNMcxXDBSE3hw0wYA90igCXWAprCJCAX3
594q/ChLFhZxkUZMaBENZpFLbiSJSABXHdOwr6g2QmrxHGkQ4IbSeH8+PZEG8CSVTBAA3a6bB91w
JrghkZdgtzghGlquRegB7w1fjqxfuZoEvXCzQ5DQYG/o5Z5KwWoP94cn86W/SFV+mZ+S4LgizbZv
4LXjvGTi2EELFVwvi7JXzL2ymCVTS0AO39sVMTUZGz6yIXIAWGO3tDOWbqhCI/vrk1ML2Z+Y9AGi
LKg4wpNP8Pu6uNOTol7g/iB77CrXJCCnLY/icv3iwNUmtOJL66xajHeqJstT1ngO62sCYOz5l29z
fE3YBORlOc6+GXz9SoVa8n9auchNK6Fz6ROWqZi76cQ3M8n/qn1vVRdHU8b6BrpaRY8gnfdDkzD7
qtx6JMmZTsWnr2WsOcoZexkGrF871dm9ncLXwiDsK/g75x9Rn679voPdGd2OkeJ01xlDcpBSQRLZ
ygN8P2fCDtaZ0YRn1vnbK+PdLsP36KSya6RJT802FpFCaYJhAWFCfd8pSZiz38uZ+Mc5S+KNJeo/
H4MQLPX1Dsz9Ixbww1SMWejtvuxMyX37gMZHuJYmT749BwRaOqntxXycJxk4BKhD9GBAaruJq0kV
Q4+14E40G0rrENQeWj12GMVgwPiXGRrkoe/QpKANRwdtNXSSiz2gbWJbi78NXSy69f2j7kt1UjN2
ACp0AnBrGvR4c5yemix4dQm2UjmrEZgUfZqZ+OPV8N72MfEK7bre3iyCWXsdFveeRu92Ysak5Rj0
6LngEn2ZptjqgCH0JDD0mAuVqBvVQtZmaT8256mzlcgNZn+gE1WzwX2bbz1BjSPVwezKih7b2Bfn
pNa306wJqhb60sQMLSUxJdpvFtbN+uK0ztjHPtG5kQ3ACwmS8XHa10vOk9tPSF0f0/VnYIqIxFuS
mik6DF8EgodbO6AlVeq4C9vp0WqrgI/eikbB5x5EnuAWvfwPRuNtSxMxwo2blx/ZwM0OokMkuz8V
Qa8tRm4wXGwk9PMXntakONjRp/1gS1Zec8Y/P8xflehN8+6mMNSskoAgXkOqQ3JHcPSoaScPufh9
RsOO/XIm/70B+p7587eZ0oox0w13g1D3rnYKjuhsjulVwhvokD9EC1aaVjN7Gj+sxHGIo0YGAF22
pKNpau8L8Wq7XaQ21rypy+4dUn+CVMpROVvwuNb6VzdAunE6VZXDo6V1cVxdSyKQp7dd8HFomCYt
pKgFm3MBBA+mejlCsbwts6CwwTzmy9x8yImuXmDRZ4zCSMlVnU2w3I9Mq+YCDw71spMyTchD/LtB
E/nKZqdjPZkx0nd8NhyI/j/DASglM3KiAZcEJEmp4+cC3gKjJS7Jaq1TyAz2oU0kWUHCNsnNMT1N
316gZkz2R7/8AvhtiZkGvZLgxXB/6sYCsMNWF3x2VGTLHnsvAHcWHSpuHhGKNyXBmme5F7XekK4k
BHvyTYS2/SVsGCkThHdy7gy6ieNIH6T3wLm2meO/60Fql5wAt4AXwqPgljfYgtC9bMsZGDRwoVUS
nyTDypipgER9REIXaM5IhrXYleKtsZNDGS5yp9lKH3gdonj8CiCq/qGoWmjHWDAhEt8JFzjWC7aG
w2dYk3TgEXk/GCDul5dlk29zPtGDrQgOretmB+hpDu3QxSawLWybMutWatXnahjQyTjeyNIkhXNv
Wp7ro+1jU5yu5N+OknHq5etvcsIv0Qc+IbK/PsRW+BaD3QcuP6uMv0qSNmT66qXm4/91Zb9901E3
u7qAazLATWLQyxjBTUNLqfBmRHyYs30b2l2NB4EOWVCcZJQWlicO5RrqQX8/o2zdHEukeeD+JtMW
iC6M+OLCce+/61yCSdRX6gS5cLrSaTcOisM3LjJuJtFxeUsUfCSMxynypkWzNsqThRgXHvUmiJmH
So0+TJ5NU/cvkevOuehbGuQqxF1y3sxfUPWWSwz5z0k+9CAOCApjzQKNN5/2ATRqAC9PaUB6UwEs
tpWyktWipAs1Nn2GcQQGZlxKsjn9tDjH7fxxZPi7vit7hNbyFhh22veyjv49+REAtYnWmmGkyh4t
GxlZk4TFJddHm9Eivlq+65rMdyHdxcd0zaMaMXvhoxMRV/nI2pgWlzH52OYPhgALbrW/QjsXVd7P
LwdjBJ0e6LiyxnflCR0/Oj9cLgY9v0jJyie5vFAgonnjCr38Q5UbIRDqqzfEZnCshXkiWfk3WkNx
pHoZwLF8TGsFuLXU5hl74Q7USFxZm/pdkjS9yNlcnLwBlgnM4UFIt0J6GTi0n7Vj1+hwIw2DCk6t
3zD3XBuZ2pX9Bs84JUnOtiIE/XbFqdfoNlIdIbMwclA8d65m8kFWyVtamwO2Z9UmEEzl9s5u9YnW
JT/+raVmTX+8G0wuVPottQZzXvyp9GMbWrbm/1d7Zy4CdKKr2eKBfBVWxCadswJBVSCMOdtg0cjB
F+/0ruXF5UVczy3gsGLzMdKsxpxIQqScZ+lz4dFTNyBArlWI6HomYzy6NAllHpfP8NRMxEqZtW63
+kCLFTGUbY9YBIct/GXyevSh2yfjFLPhIkmZuJs9jrgxCoeoG1EibKYLPIXnUj3dNysPEawYaRxi
nHajkD1dHxKw2sCirK3l5AoRfhNhQKSk2Ydn0KunFu68W2Ktr4c5BSKRH6d9BcjDmAZmfHagXaRN
PJsoKmUY36WaHCMBGIsTTNhnNOMxXBa9HuARomdKt1ZQAkChce6Bn2LFwOhYpUymGf5h+Teeokib
lBC1s7rNmo25uUr2Y5Z+hB4Nvc466ppwccW29WTsGizCM3LB/2abZM+zSaqdB+6ePl9YT26Gu8LG
2MHf6NQR8xMLnjhAROHWpZZr39JwHmXaLvjri8lk+2zItgPUcLXILajQnQPBH1chHg1+UiwbQxsd
05WhB4mE6D57JfyHEDJr0crSzi8FccIrUEEjg/VExS2lB+jbQKkdLyJcTD6HhrxATP3wQ+N380Qc
huen83d/AMyXxNYQUO+31ufPx9b7I4x3Htk11gDOSZ50DDwbb+BDHY2hu3lPnsPdJgUM6WwjY8Na
9lAbveGs79S2BOcEeSz0g+CIwDCGLgacRj+Vgl7mfaRGPFZTOH0TCQfVKXoyyV4pyDPkVJP0Zzax
FQ+9XkLdJ1mywCzYqYetmCfUA0GODoj5C4wsZvS07lFTiqvhn7R4T/yx7T9TPtt1mdZ/FHEKbxGS
O26ir1MiwNdEhhdGesh3Ul3RKdRfBd9/8+jy7n5AN+ixj3LFk2z4x3PJb3fpI/+8iscZddhsV9Jy
9VCHTX55zqXh1dpiu5gL/CbW0aa1K8mHlM9usqH1XDFBeKEV3K9PNDl8DHeL8uNwZlFUiqlr2wqV
HhTq2vord/+FBqV6x9HYigJmgAAI9enN9aX7YVaxjNoIVRUCuPUryw2Tw0Gpwgyx3Tc4Dt3lvyel
QxRgdNmLTdOhNutEkX8YVhGwz99I05G/T6VtOtCRZqrnAxWx7LCQc/o5zhQhSnxbFMx+JnghNCT5
qSEs33VUI49bR5Ybk9o4EyuVMQebGgMgNvWIrHdwU9YWuvdGkusQXT8IXorrHHic4TjhFnhCiHjJ
Vjg1Ya1eSo4popHHxpXt+OlsqwHe2EABe1Pb9OBSmeUGALvHom5qMNQ42SOfSmNBAcFf7apT4ttQ
82vzjnN2y8ZhuVuvVGxAwZNJvbIDOAGEt93Ya5/4TI4vkNUm1yPi6hb0A85EhoWqR+qcHjDZAIcV
RenmCtDuBQPv2+ZOkO6IH1Bb6q4W1rS235lcuwH8lFp5M3L0GuTCt8IOpwWWUD6hDkECb6vLdgc4
JITe1YDkBtqQAjHGnV0FMJ1G3gLcfxhYkGTD4QFlEUDboIAaPg8LcTHy0Igx3hdlipjS3K7HQsNB
3608L+eGed3PftOUpJR5Xznh3ULLs4Qe3/1vk/ini3rm7PGJhDYlqONJ12BJ14P/5NBoQVabiSzH
gdDGMcrW24U4t9wfJHo/59DDhGD40Eeb87GUOFzwoluPUmGEW8+8Hc2hVz8q/DNwhGjbTmhEp7xp
ooOh4TQUfUBAHzPZ2mt/k9GI2A5KbrAT+X0re95Vk/n21950C0VVRQnq4KjMUVumRnpm0JU2Rep7
90hTB7X8b9LkXaB3P9BNVC/TkubBhCu0BskRhRoiM+FTeV3z9xe/43eptmIgBsZkF9QXSU9HCOjh
CbUD1Aq3DasJY8jVubBEpIe88jKrEGprMcI6U0M5XObMn5Yz1bcnn6rbA1Sr4+JIL4qiHZe7GSUX
nB9iUtRhXuPyyoioU3W/9s+apo15oXuZzlGaWr3LKOG/OmkcAmZhQGvnP0B69N2F8x4RWnZFdmfk
RVt421YzddRCCePBXHYrrS5UXXstVivJieniB1VRq2TE9ABxXIbd5sRka1Ru+fQVD1BzXKPMtfL1
J4Z2+YfZmn2TDCGqkzU/mPSEDSFD+q+IUQ+LtB4FniE4ieAeclbFNkg/7T8bNZ+6pT/BdGC+6SIe
PBzpvDwgUuuslDO6TcOqTynyxzd03SERNLRNu4u7iNp/wbHIc4hU9cbull4jyfw7ux6fonFsnkCY
WitOyo8ZfCqpmDRqFSSZsjp28Boh6mHrNCT+NJdDwIz9KLqFYtzxV4yxDVGaPozhniwHHvBCiAdo
QZ8/z1pp1vmXNYYLxTQijxsNM9CUJlkKKtowV/NtIDZKV6RPPS0nUWzELB7TfcrI8wEAnITozVF2
q1AjWldH6yOYLdNtgJLgYEFXmkgSfTR7tw3irPlaMCMn41gsmZ7zvVwqY12nYXlDSsmeqjmnV68f
I65o4kZ70hfwSokndNyV/LgcPrj6ZK9o/W/VicFVWw9QLSIi35tjFLTykIYDVquR58ofWAV+rsKv
WWjUwLAOhUNni/yW/1BOB58I1vHxhXbTYJ2a+1WdYGoo36gGC8A3oXJTYg2zVRgwON+F3qnFyb2A
umcphl4vHbOYxo5QeaQkdSnGtUwMoUrMBOosIXVL3tdxKwTLoeRl/rDmw1cLYvwnOUnBM6iOcqOZ
cXKCCjEMB0piVD7VeDJ7Ba+i7MGtmuURrSmcG1n+tZjD5DtfeYru46t09zm8VntJEulc9Gi+zgnL
46Vr8eMAVm7JOJdBlmfhUUkOZNtfZx9Fu1twRPopZ8TpS8+kXruQ4PEpvO55KKgo7gfyOHVyjbk/
QA7Tx1sq7SDAq/DVmmvo3negvYBkyHkw9LzIwv8itkjDnZ79eq0PfDv45iK1Jv+AwwMOXux6b7gn
/t3Np17nS7E44NuipmSNTq1gve9SDBLUHm5FLIsT6U8JpgpmnLHHJZTOnmV442v3xInusOmvufwz
LqsnWIC3C8KBvTlu5eYoDebuKUq6ybvtiqioeGmIaIPazMcjb5mhTan95zaSiTFJZ62o3ta53OMd
W1CrOV3on0dHxETHfg7wOZZx6PUTBIGTX49c8rGMgzSvvePFRg4kuzqhL922cT+Xe4xK1Wan9BMC
cZ007452/KwSRMDAlcvVneP4vrb+jeO6Hv5RIF3P47dVEI8sBVqIIgPkbgkhkSu5oWf6EIV00ApR
qWBg5/miYHG/wbqP52DPtBYRTU0tMsUxiLvxbeqcGgZXL7+gLXV5BHe80A14JKyB2OZ2D00nPRaE
QBmgVofNXzaCSUonJl7IN3r883X9vDysi5rwVtmLpbgAyITpoOwA/IzGWNLjLbaPForbvKtUa13f
JPwtv+fI3ZWzXtW1xOi6j7KbaZelqofbBaDuQJchFLkq3uLz4+I6fGAgt4Y6tSk4okfsRYRktvNc
g6YPLJl+9nUqMKdK6YoAozf7dX57IpqlFZKl0JiKHn6dNjuFeckr46jXiHb2Sz394ts1x5R75lDm
HROelPhqoZK5LxGvDH+c748EIza1hVXcJYmxWzMJzKWeaShAmg/50M4iqCfDuGpbOLoCFmFGC4WI
hVLrfDfNPm5g/ufa9lIjLHUk4yQEXbQ0wD/ue/c+NyoBFUANfkcz7izwieJAZ3K3aUCpvtWeOZAz
N7TwTTMMR+wQpMsluj6b9G6VY11Ul96cqW/GCrq//234yZQalZ3qsk3zLLwnIgWFr6qgWHjx3Rzq
oRgHYI3Y0kY/B3at5h5mixJKIYJ9h+9CTFBhiAnTQNHdp/KdaPs1rZgalEvbYVnr8DucCd1BSyNa
/T4BcZ7u6GuWxaKk8Quub0epveCKusU5k08TzPc6MlKmNey/xMGDEwgd9jJgykgsC2ctOt7i2COD
x1WBzhkD2E6eRRAhMI3D0iHOGEogNaF39ov7XrIZwzAKpYtYaLmhc+Giv6VzWhFIj+3xRVR3R1tG
p3IAHxK89mBFC4Q7h60EV6t9SzQmOoE1Sa6/nBHt9DKBHdc3mUHqqs3DkAN/kCSH8Kng+HVb+d+1
OVP6UakiWdUZ6VmKCNUjGPfef6ZLvuyqpwz/CxANQVQmMp0uSrqq2Tck47vNDIa1h7NexOgr8oKW
NLOSsNl58c6H6BX0Dh0KB1QHYnMBDx4i6U0iv6UE6f8LpJtJ6wzc6bwhD/RrHI24yQeanzF8hbGN
GGRK8BAtsDuX79T6JdMFdJhzft7zUbGwkHL2V8fQVZVpN761TjtJKSY/OTSzy2ogx0qbQVyeZpab
zfW1OaVO+893vdSHuhn231OinOvs17j+MTlFT2ug5urZjW41emji5VAClWYoM3bjxhFrk2UeZ7aP
XmhWLw3xG8xEfz2X0R45i/EzAbSviq27bhnZY/Q9dRsxuIjnlxi4sjeodjCeSerMfYuehcxcd8Gj
sioUMJlsyI9brPBHn5TsFvEnlgmV0yYXfBr6oOoISvvbm6O+ASF5koGmWdWMvwwHLA2c2nqlZaMo
dygMAETrmD4dVG6V920XOV5D0UBvkXizeMW0xshHHM2SM0yfri91k3j6RTmDswA3KyR2pMYH/9F4
mkCN+iOkNZDXQUQtU1hmBmX/kE4Ik7I2/usT7/Wl1iDgkjIisy/c9qrpV+yqxavo/a1hjcWc6GJ+
N+cpfFkaX1zdBa/rGRSXnuFGXkKubVROVIcAUCi7zXZSXANxe2COmy2LtQ8eVKOc5Zy3t6wIHd5k
4dfNkFXEAdBvJn6ZPXLtsoHRp7QZfi12aGL8y/ZNZvyqm3L30eelHRWe1CrMlnNd917dJwepikNm
c36SkEDWNywABFetVZAEWQ4I9EjkVStUg2koxqLNxo0yIpB8IhPWbcrWLTy6koDPSMVOKNyRqBBG
5QWn4oqNSxwafMosAbA+QDFGUN3SD3r+S9rzm+YDxXdqKxcDP09ao440ZNbKA2s6/Pow3ktevxG/
qErH8qS1mCBCZ+F3iET+mRoFroyA6ov6nNWJxylpdKKYyK3mXsuP/JRYzCJTCdHE1B3KqKo0y7Cq
5w1AYgbS6Bfu9GY1cDxrAj5myPp++kDu7y3bBNv9IU/yJW7DyTVmGJb9JX66NqmHv3fMQtEjkiz1
2kyjo51zXftSTU+TxZ/Q87rKeqdMqFtKOdYUw09nwPqTnj2MZORTquE6d0oybUXfWU+nxEDVNaCg
92Ceaf+J/+YQRyh6XwaNMEV8aJotm/jt1qtDbIXc0BvomsgBy4gPBPO3RADYUg+gS/mvL58teQ5i
+vt+sazP23B+jCd/sC1wq2/GRf6yaU8LAwm/RPQwyBP3EqP+pwwHAhptlpiHfMSDxrRlk3atY7Tm
V8ODouLY+Z10H+hlaOa8GUuAVbx3yVEWicVkxhd7zSN6BnN8iq/17+7qB5chFWQCCGHF04mgaRo2
s6vofQ4SkqPR6U13eYh0ONe+trbpEyrqMZ1aCjXnPvRdFqq8ZBkNaA0cY/GUfPx25n1IWP/Vwo2y
Nkz3caJw32W32lG4AYdTSC7Rvkc+ftGocuCYN4dN2gmjrl4W8VrxxSo3yhTC6avghP9ayyxDdZia
7/2wT+6IKN7jvqK2AO/sQBARqrS0vJ0An909wVi8QMFTHy0H37FdAEXjFDEsj+lelIwnQKPQw66B
8bVJvT0GBZLmct7PnEfRVdDepXcrMF7xnBLKx+EE8HI55+qKAgEf2QA0hXn1K8qxma1SqSL3tpzF
LUa2g4tKvsJBEheVnxunEnCZGv6SDIYlG+3zfiv9tbxn+W8pT0UWbdZR3enkU7wQymHw6r1NLMoI
1jVLR4jBkEuOkodl09hbr03GG1Gc9ktXA+9pKLRLjnZdL1wZHQwlNJ4Gk38/Q576p3i70J+Cf6RQ
iTkzSLMStzXjYgCcp0+4xq6q0aI+dwM6oa66Xk3dnnVLt48e+k4NECkc6jDadCNayagWqCxCAD+t
1Uff58yMmvqv1a/AxC4ybgZVuhlfDkSfmUFSc4dtKIbHZ4MHMEBYmJuOxuQjxCaQKH5jinPyCe7L
C1Au9pp/e6HysICEyvaOBOleQ5mtYuGPkHSI2Ho1XnCDNeeCdKTmwA9CmuvDnWmw+Yz8o2YINo9N
m5xN5M75i+IWPlQrhIBaBos1SZOIqG1wskxODucLXMCMHqWoiwceYNcH8Rpn59Z/7NwF9lyYdMae
GbxH2Lcxgibh1xylfRIqT98c7izqqa6Mbc/KxAoUHH3KTspVfjFwAKi/wfjD4nAO22TSN5g9E3HA
tL7lJDS7VW6ECFdyq/ln1czmrijPbECL/mi4F7txZOs+L14gjEtpl9d26wH8IwEJiDul1D5i4GzO
eqQLXgT+OxAlsyb/AC4LhfpAZvAvGQLs4xmIdXETB5/lPb0MtC1ffZwZpCNQVRX5JFJCFQqS1S6p
d9L/a2gBJghcnYquTeHEBxDhEP8xpntb55eC0eeKgDS4i+4G6uNsKJ2v0fZvrbQPfdIFGVOhYlPr
D6Xizb2WRaIZT0IUx0nxSV2bKOSdD8gEUqhmt0qwI8ds+XikNg9VYCnY3J9/Kg/X54UCLkzbTIhR
pSbFnaL3nTeXzU5uiD8mfNOIWmg30zbzafWCViRX7k96vzd7VtopspfKsk+bXTlM4MoHTC4nTV74
OJLUV/yz8wNBbxACFFo29InC7DyWMD96m434TKZREumnCsm87yJbVQPZRDfjnXiLHnRFbfnOaCGu
mSbL1NXFAtxaDAWFzq0o3wE0FyFPg/uew/qi8+KAruoXEiyeMOhJidzdYSkIajQjV6HO/hARUHlO
PRjSjBj9Q6CMsIQFBm5XWz8/Ew9SXnI7+2hq48ZsfiYrh28qIfC151Xcu0FIab41QlCM9FhmrUC4
rQ+6hy1XDDIaDLrZFK4tV63bZ6PVuEM+Fu4XgYxCD2FIofFnYG2YJlUc1NPHMLHeiRESqPCEuwdF
1kzx+GiwahTOL/gR7kHkzB8cB04IRH5CvBPnJYgXzGWAdM/OYF/82INv32vJgV7hriPDa/xv23u9
ZKVuSu6s0iKzMHqs4N7yPeOQ77Fo0HpYwIWJgSL/2NFI09llLDrljg+BK/92vlWVH3RkppTU2f0r
Np2aHaCdXyMZe8dRWYt1Z39QIJUsOIDVIWj7es2HjKaRsThJNpaklK1OS3cMXKXT2xREd3dbr9nY
kEKiS7DpSML/ww1N3drLuPquJZx0w9etIgu9illrPqEMLopNBmQZPLtTzBMrQuh0xRnzrp1whcxl
XDkUbArnpMtOBQRFgPh6GJn8gekTqGbPosCeVLy8rSRib/3+BCdY0KXRV7dk6Rj3Fq7Ogro+hmaK
xUmWouJTdge3PC3Jh6A/wwKz3tJSw5ZB6z9/7Zt95/qbDFBpQ64FNLcDxASax6Bh2l7nHgG9eJbS
UrO78mfWsrwzgzEcdDkojnPgooGY1p1Xb+DXmbXhvmGnZTFALa1x5wKF6AZSGXjiPU8x06IzWFDj
GgDRabZOQLxZCKGtq0xgVYVtET2ksISYOvdnTnSQ3XkUWwieyP3YdNrpCvXQ4djnyXKTg2h3rLi5
nEG1kpHrnwN0H1CNV/Fg4rfv+r9ZfHFwuwQuwexhdDIADDXpOGwxiYqq6b0cT/Z+6q6V5/h8cric
bdAU0RKTn4Otlh3gmzU8PtPdm9diupbxa8of6DLeoEPWQnmkfPRqWCGS4vKlf22XGcaWNP5+oi/f
ouwYY3saO+yqD5k9IUBCj6U8rEafU2NZcUpy9Wst7E9D41aQH8HzzLhnOUrDg8QHCTcU2i6kW4n6
pIfOL6QisVVTU4OBjSPS2u+RB5FKgC0r53qj0p+lrEROgw8RlofjrLdSAfKGd35POmTtM5A8StQk
mVWVWKT8dxvIEkliuraGPrMomvNCF3UYxM5AIQXjb+759VnN84AfEx8jFI//rocMe4/WP8jidPhn
/wRJZFJ5GXxgcpKABQ0XrXvR+jZMgIDt9nBTiKUxSNzwDxs1tRjqgq53twhrZUovKCzN1Im7uD87
MlXCLFrT9frsLWlyS+Xeq6L1/+gvVoY2+PpgX/8J38j9O937AKFXzgR76csAMcRN3SfBVwG5e0w4
06iHiLUto8byWE75jrBa/bM2joLU/uipa2j2p3YScfMTspYzbM053kuY21R6g4VtSjc0r7z1jEan
z6vcFjYHy7akS9EZPkaQpkk2gn70x8JEP81L6UEKG2m+U6MxCrpKtoBwfHkjjdOW8ULaNkO1rda8
WtO+XCKdQp6fHcHo3EmRsgOhDZN5QH6+Shc5SL5NNUHX5Q7EGBf/LVjK02BMhhYApRYoYgdCgQWv
5uPVoLgvBKPZ9HM57wFrA5koOI/M3qFME66OmXvQdJFizLl5N84v6HUSdjXoTLLOVNsSiPXCU/BU
XEPCRuPBgvRFX83fwididpKER7YADTuG/pj00vfeIVhI2dIQNLvgK7d2+mEgfFhdCnAq4IEL4/fo
KOPWp0+egID5pqNmlTX9gIvTZ0+6ZVEqMD+sTbMEU6ikUqVE4wu2OkqqKS7eN/xxpWxTCfnK9mIy
yzorf8j9eiarjq7L5oYtgP7iNLuSmiXXJ1CngZFKZpy9riqCvdjOQytLbAeCJYzBnxYh9fwh2Vm0
beKndz8YDrwdm51aOLX5QXe9ofixk1OtcLMPjORU/xDYVzw8EZFqGwa3wiv4ZWBIQLg2eUKvbBX7
kFmn3LvPV+iakHolkNKoVs69q/l0NLDKwKLy37Fw+Gpb7TvOq2690ZDDGWDlhYNGrXJZ8TndeN3F
obh+bAU5inmwjcatfgyZ1JCwmZbDywpYxK1bt1SDjD+CYne/ep4SesZ7oJgQ8WJsn2ifcUeK/on0
B/wAqs0TDs9GNEfAQIi9Jb9OsZPOH94ZVh1MYpKY2SQj32VFSo23PZP4tjgU4UfxmWGgyLGd6Hyu
sb6XSXFxcwG67cWLtuOSvIYK3Ot9C0trYqb7kdjmoaYRuo6T15wGG01OPYSXgdulusV+bsU/ChXd
O9LTg4BLVO/oES5wmsPg6/welcpeF+tdzEfcbrZMlZeN6BsFoNHNA8dpDQCZHc7JBGbujeaPJHWK
72gYkfl+eDqWzLAGv5v0CsZwQzPW3042Z4ghbufrtOBt9nZ5eCjg+2BC1WulFVtIMzSppE6fmTjt
Yj7bBwf1q3xFvE9s2p5Q95wozRnCK4SR0RT0Q0lw5Nk6vERoHzlm6aC68XNEu9fU1L1O3JXQcgnn
8/Uja3siTOwyGWVCmYhAjcTYV5PiyA9PVwBfiA4/+mRKNIxkBmWiaH+WHq6NEQEVoSItokWiZ7y+
727b7qw/dV+8I0MZW6zHdODI5HkML45/kkppkA2ogc1q3PIKZzW5MuKlr+c6Dv75h4ofFe9v5ISw
UPMplY0Cnd9LaFtm15yOt0gOiwWx6kUrB+Hooq7MelnM5ZPy5PDbemmCcck6mn9eGY8l78GmG+cc
RNsk2YQ1jEOd2Sa0+oYjB5DtfxKXPnR4y1JbhUQOHdG+1mseW7tGtYZJoFaSIprC30h1oMBd4Swy
6RDog/vSkUw+0el/yn88dvuDr08t0ljkDTF1uuOk8e7FOSObVdqKq18PFq3wMR9Un36ZKci1TLNb
EePk3LR+5w9RQqvVZ8IPzvA2RAEFvO3kbMz35WRg0iBd0Fme+sEaxCmWCIltiAtfV7yPiiW4Ul1M
ilLP6E5M3cDNi9UCeeHAVn6lruOaH9e2k+PfR9psXkR2njkVYiN3UiaBq55u7+k3uRdzGYkkyUto
Rmu7m8RvAx/Xdf66zHW3QUlI/3kvPyPPc44YMJy6Fn+e/NwikHYXxL9s9FtikI31doVbugWji/av
F6dZAJs7LktkkRT6rIyB206+hxR1du1kkKTHmr5PRN2stpEDDaiDJseolYcvwdM2yfwBUxC0Yo8Q
ppu8m7/hN2iHwZV7hcdrlQta2gXGRPDu0jkeyb8hHqEVez64osBffIU15J75V7tBuoKmaSBB0zdS
9dhJR0prsmMWH/5N76TnvlQlsfT+wY0eH7LA4Ep3NUFM0yKWKe+gixUHzJbQI4afL0cIFIoq6vzG
o310NCjq3HNB5mKi1sD6JJf805TnFnXigqNDGWYm58PAT6gpOIHd6kcYcWS39WgMHvL47T6uynU7
xVXZBisKV5qxBN0Y56dKAw6KFzVqZEU8WhbxqG0caaJD5HfjuSEFpp3qEi5dV6R74hE2dp5b5rwg
6kGNBMmdnzz6eH8BFaxli0ZoGNP4GxOJ75ugwXag+zssUmcDiijuIsAdmQFgdwzDyALCgquF8iix
2Faalreu6WAiARM0tZUwKVrGtw962XYnkB8u8ZIFUvPFxcrvq9IasR7clUVzsNpT7ON1etupzJtD
dmQ8Zq5XALEsKzMOny9DV7Oyj5KHTPpiIY667YzmqJAT6cjWnQmnCmxgbx6bAKNvuOPBFCAhbRZ2
v64U7gABlzCZrOAxt6Bht2yt8Xsjcjyhq1vzr9Nc7Et48UW164+FW27AlI0yayWxJTHicsr67vFl
R7U0yFb6sQJ6aoemfmkAYhTRZoNwrHQDJv7l2LHw4hlbkUrxhrUiaBGtRf3rc1B+BFxQSfEK70b3
i6XwkCVfD18mCLecHVaOBhST8OS3zQmeQ+nlDkCdeccfp+KaZ8uLBGqBowG5Zjri6qDU/ZDuWMQb
YH+mLKYu7kmCNxilwS3VEHdZ+VEr0RC7EGmkrP3sbdKM7MAnpVckQ1DIF+YHrW3AXMV59n9RNfnZ
zh5/tVtb9j1cPNoB1uBRA0sQ54K4aDNezEVW+TIZjrqfAHIkHzStmGDwUJ0FAbaloNDNcnufBtxu
m8Grz7SuMqeDd1cyTMgJNJ8qTeFC2wFMHxkEJaGHx4ZMtSvzqYF7vM/lUYleK3lhQF8etUlWOYvq
1/QdcFwai5/ZjoEvGtWO0R9qrdwQrvubIWL27LhM68E6VCHL6U80j6yEB27jjlADr80HZ6QGNgW4
1FhYvVQuOZwlqM5DXxD4g6fEwNMSMT903UedfKZBzF2Yvc4nkAk4WX8rNDTuRxGozUxBotyN+Zpx
1oZcLJE2WnrvmIbEtOwWIPhhA0Ye1jtdg1L1WtejHcNZNRKPBBVUpZ5xkQNyGw/B06gZi7ThaPkI
IT4QnOegQfVqg3ayMziz0qYyfEBOAutRto6DOTU/8iCMMLzil+FjR9pTW5NEAeMEGIrYjcDdon1b
l6XAU+U32w3J6eNPE0OJ4T4VU909JA+KciReLwUMPQlwvRqeSHE4AVtsKmwHoSHEz53hx5Bn99BH
yXgbqKIgBbIErxzO9uLSigxfJZML6Vdk4DHGYh+GLG2Q6NhocGEq7EsT9WrAzXRyGw6k78tvzpBk
lCqo4fzelzQlHHHAz0GkbkuUq8iWu1ZAiy9+nZySKuc1RKY3ljjMbck5DI7sil3/kiVb03H8G16E
2Lio/erEq++af+V4++ZoAM/3yKIMWBLPcrly5xJqCl1mpB7T+CZ/em1rGOJCw6Wrerm+3m8GkXs6
upSpAxeC7+rK8pqw384X25Za52hDcfyqAUD66ZfKsLEolsjY3gGdstwPkZ/HKRt1mBO1u58rTrwx
bJPk8J/racD19Iqx5FhQgsW0+L7MUqm2VEdnfjTPbO5igy+moYjZ/6DjQj9+8witFbZxb4unRnul
QkhAV1YiWYcp5fRyXnmUYgnVTnoKcrcbhw733ILuxfUv3yBm036tx1qrqjk3nFucMSx3cUkqVFxW
FWp4g1IFtdrfeQ6VrBPvKUwY9k+mddlESAgzjjg/SrWwbw0lv7mskbx51iRLGXnA0/Zpxh1SNL3U
Gtld77qjpnyPcbs+zsmRqL80WImxLhK00plRaAlKyN7rrdPIhggNidqtFnOMW124Nd6OnUQVzxTT
i1Y1z+eEZR4tUxWPKwt9s7xf0d8RxRSPF6e0KKrGuiAeS9MZyfNhvaxY9TNQIuwoYNGDUvQh0F3U
hcaLk3RIyZzdONvMX3i4+Ec6+HdKyACOgkf11gpN3FBIISCZJAVlWDBFReI8DXWCzT0MJJwMFRUv
pCRSP0cK6q+26uzHrT8WEeuCZbvX+tArOa1C0ZeiAPYUfI/vpnIB2XVxo5oHsO+LBAcvyHwxXCaH
72UP2yaFj3TUXnryTtgIPy1cbIPJhLjsIzJWSIbmUxs+xTFLJ1rNvTRw96PpcQ0aPfYuxBPVF19J
nIWmfIePgePtCe0/QvZUkxyR0pzXFTO3Amu25PsgFMXAGNTjbjr4SWG5KoGxSXJlFjaFnsIYX42n
Nmeh9Y/ULq7fprmUDmyvDBME6nIqPMZ3qsC6beC7Pop17RGS4w5572XrNETrCfyldR3dGUd0qzFb
KK3hvseCY2D9xbvKn9W1SVzKhI1VyzqcMOQUW7Ya5zD9pHs+QE7WudfuXWbuaqFsEyEYRR4uy8Ou
kkTLpbSTutd1hF0tGSM+4deAwIbBAoN5lcvwvJGcwVa5Q0zOWR9e7U46oqsmmwbrE8EgIBrGk7vV
wFogP0exuPwu2HXHxma+DhXlkZTP5ycHoiW8qrK0aaLhD+rGwG/TPYJnRkT6x3dxITgR4E92te3c
I6d6YwQuHPDwt8exlqxaz7wedmlq52P/nxbCK/cqD/skJBKgAQTY9OnqzozwCrCcFaMP0QQJ9MGo
KhkDYr9BngpaifytZ23WgF+/CGJjSZQ599lczqwKsNcw/7Ne6ZP1AuBRxeeVtc1up6WhxzDU3c8a
bXvt+LM/ikHQzRW2nDQanXJJJHAeE9NFuxJ6EvpNMVD2XJZ1BHd8dSFKJpurSXQxvp2IdBf6wyMI
U55PA8BUsULCkq7M6zRiexdx7FFM1mk+cFLJWHUN0FvkdcDDEjuqNuWu6gL+wCIp2g2c/qmRDX45
H9nMmr1Ilh1tDQbOC4mCZ5qr+vVC41IWi9yMF308gPjSttXprGiFNDw6GqfiNKlANoW3ERjxUTfL
fuPPdJkAfPiCSx/Qa2mvgFO0L2/iH0lg3vqohibxjQNlxWIIGcz/TaupS1Pq+O99wDvsEQP9/0qu
cECKAiryeGKypzHHAui97ermguRcmmzxdDq7TBgJtqsTyhNnMSvCmPiGWGoCTLzmzXrV39m6yVTG
G+TNCGHEGDs6tORDLKqqAzNfXAOzJPP+jsbtk9iskvt8WKlkMZ0p9ha77/LW/q0s5icGbQUs7aQK
F1ojiYXmWWbydAFkJ7tQW8QBZDL+7wHmiu4+RchapTNq63od2oWrdnKFwVJKvDWgT5nxNGIZizLK
iftDLfybV+nmYz0WU3oxb6gsPtZzCgXIMPxIafymSlK2UNDvnlQMmLs1xFTaBFVEc828w7oRLYAG
5TSFtcJgyuLqqHgx4K+42SOZFRvJBERY7BZyMIfCYmlUcoLFv68n3mvPUHAAPI1a5BBZ0DC1yEwL
umSAg0lNcQCzpVxYPQKb9XuHqEw8SN3N8hX5Y0PM9TouJdof7VFkEzw7SNj3IPcFO1ws5Ut2qmLg
BaTHnHuEN//DCNFxqqccOxKoxwV/xGTDPbppRbCWkFV4/p32/PFtiKxC8muMmanhLQ7LU+WkRR7B
h0mc/X712SCwa07gzkl3b8eLBydnwyuwQPRXrZGt5V8MJEktRaOPtk+ioAwquHGPjR9rFfLAkapH
FoB3cKdz6m+HMxciQQnm67zUOBkvhjGGYehs7nW61AR9yqfvtDpfvWtgc1Tdt1oGquZKIAc9I+VW
5zONzJa4ZKxe6ArjfAgJPxexOVBqJnFepXb7mhKshKmv+x7UI+bGEQO9CLGYnfas6vBP+WGYfWjQ
EvUcuoOPWygAIzdq+N0mb1nnDV2t4nMGfJS2OqaJvVBs3XaO7+DNJjKZPuKA66CT9RU098N/nAVG
ahzxm4mHt1mAsia/UNSrScicuoyZmWF+EsSiImiNvNtMP7kSocTMcVip2IkgyemUjByznup5dDO3
Yx8Sj+SBDidB3daHERzvWTOWP3mdy+DEolyunqdKL9jkzMZwUf98yAIC0c2HfxB4Z5u6u2GnGqNt
zV595o6oSJslLpEgNL32yBRXLPGsQIpea1bwEp7QbVLimZWIx1WnqmDmKdVJGPfsJSNHI8nysSzm
R5SKwyWXgG13ZBE/FO1wAmVaGLOWrCUADHmxmcdpFkX3go7eOYNWJbtC8q4tVYWDGQ7OrV3Gg2GL
mI+nK0fbPmqiOnSB2XZ0p9YDGHfwRq6FLRkPYfYgA0AkS3tOLSUx6wGuNpkl9fTsuNrODVJM4W+q
9Hq+hfID1DGGcr2RuJvD8x23m28MHEWwtv5WjIg3o8mUBVeJY9W1Qr4lrViSBT1HO+MLDxF346ht
1Y0rdlxQ+pOr6GosORYkX4tEDhPImlfgVh+UcvTeQxayj8/W/C70XPXti8YmtNRjTjd6d+d3dSsD
X1quQJqkR+sx0DjbGNbCQFesSvZxgoB5NHitNR8l2/ktvwBlib3tFCPwKG03T859hSltzRZYN4Uo
061BzgG/AfEd/rvxnqUUNxJ3lPXkXf1YMaC6BYRArC/3jaziPI0vLrUNOx5FkWID54ALFlepJMjM
l75aZciaXkmA5tZcFGSG5wpSmfWfE33G4gJ8f9D1JvgRQsPp6LHXxm2Lel1nPa2qudLUduNwv5V/
i3QhAtEa2T396ZvIvB1AIQfIQ2yAJTT0q5zhdJAvEfOjuUhIpvR7OPuWUbBgTs5eEtiJRu8JGSHf
kOtVflwsTMXwQpk4dU9kIc5g6z4Ny8+dRXyOU1gozZ5C2x0kqGi7bJP9G9lRxvG02n7qgMQtipIM
zDIEufI0ryPiJWAsV4GkTXvXVTWoa873MRSkSORLwAYQdM2Dc6FtIKlJQiomHVLwfent9TGu0NaG
w65gNZW4KaRtlGq9XRmahbswuMziOLxGmqerRaBvY03eKi+PKiWZ1F7xJQ2UP4FrL5i4KbY2Pj8v
l2rlLQ4qvuBMmkwvq1OUm5pml4gUW+ZhB2bzfNEYR3rUn4c3LHVRgw8xAEd5c34NheosAOAFyvFJ
zZ7OGIhaKmWVHfdagoIJry13AZdMAnOREmOljbViNXlxFUKX4lc/qdyaLVzH8olPu/AzwKQQSt16
xSm0Zs56vwo+Yd5IF1K2/IswthspMQ1tqvbjuuR5PaombyxlliOuw93qq6A+Yzgor+hLalLzeuE0
Gia17tw4AAgNVX+a1IcZ0iV2J0oGtI9JyaPo+omrGv6s5rykQ6czRjaER1HleOAfgE4vTD9h1ZJl
Rz0dPCfoybspEENC+ILysWITVCCFPZ6pVCbM94bxrKm7MdNub+r0BQ64sirxjQe9FgwJHhfWcNgu
rILqF3XfXoA8ok8V/FpAiLsqDHjRPr0B1x6IPNPuUKVhqYAn3FozwV3aQxF9e6ELSIYpkcxSVwwT
1777o48APu8BwD9xzosaBHE9PR0zy0to1DiiSnoOcQjgeKRKvM77sJ50VXV8tJpBkMjsjUW26dZ+
GHM07wYiwueetZ4XsGgPUnmEVVpyazIqxW5J1pfgAEg+Cfw3/Z/kELGaTpNRCLunPH5s8iqVk7QE
Z2b3oJXfYsHuqaIoBJ/Lic3OpAyaHCGs/YHqEf4gowlwvAydId1fOI7Xc8jhyASOcpUqX2UgvnDa
LNZfrVeZYqmlVQSFikXh49xxEL2AGMoQZyCm9vwK7hiIk4MH1WhtUtexBE8NVtFfB3kRPNILDWDw
P9HXc5jCHRf+GmxcDNPpfldjYEjIuWOmyiMhVONqnxXczmfIqNiP1BEQgF7Km+6qYx/miDedmb4q
x8QzQfyggb5YMEGSdaZ27Jhj+9eBLLnIdHVIN4qn2YgA6u4iObbl6KczvvKd4g6l87KseEiv/sLE
6mIXV7iUF/mdALkA6Wt6x9VuKRDxn7vluzbQ5QskiNlyetwGRfRyd3BkKFPhyFTruyMk7Sf+H/J1
2YzWFrv0PFteW/gXYOinBtji86KQ76tAiG6E1Bu32sVWYzqIsSuwVTmMF5NmTmrQsUCAFUFjB00L
MaeHDb/q6JrofO7M3Jd59uhccUv3w4xfu9w250pDgZyP3rCFpBCeKVsOpffP5Tvluf/+6Pumkq0r
UdDGhPsBJLDp0ZOOx9a0lzFpYR0U09L6rVMogYTt1vuwOAXN5azBJUBm3qVVlAxqyJus+tvdU0gs
uFz+hqIjRpu/3h8SUCPGSWe/lTP1nstyXAwJRlL9kUlPTb6WnYd+cqYwbjtPljnduPVHseBW8Roq
YlpZSwFmoygwpfLmayOsygaOrqmgHOkp1pKRicduifay6nL3sUbVrY0zX0n/ODIDgtbFAcJem5cZ
dQMdjA10EooF8yXYeuNjUJQ9xucTgCMdH8wmEZuXkIq2zpe4p7bk5B8OXKdt3onfVJBncf87rijU
vHZ7Lxf7J2w2wAFqHmo20NLCoV6q1hsso7DY0mXmddggto8l1KV0wdJ0pUPiKCCvxCSofQqTGf9W
FutgJisiH4FILhPgFhG1XmoHFjcSnVSPOKf0udib/lTmlcGTmn3aURC1m0Gm3VPSubXw9sppDCKV
jy5j+/sWZORvupCoZJQrO6yJALu69yZiAlDghW/laiugQC6XclVc4GORvCxL7tdNnogmHJkzRYUk
PKAwBe/oF5P8Wwo42VBRuKA3Mjr26qfqyTrszlqWeySqLmUX+Oi3rJMBPqNSUPaGo7T2+HI7A5Ax
RJHuZFIgU1lck799d1VBFi5mo8JQC675uoeCZQq/IJV03T4VCO2w/eNbNRCApytswIZN6mvA4hJE
Wm1Xz+gLuqCYejq1RL7X3aiwWyxYfXNUbsMdqpRakdDsJur5OIPcLqa0Ap3X6f3ClQ//FRvP9aeC
AU6NJRrFl62NSR+QbBOelCe9K2ZO2flUC+Zw/K++74kEn2Dn7I53Le0gSunS3GcECUEpJcOhcm3S
t/hlMVpZUmzmuDtFj5BxEQ/mtpY3PzRX5a/kenwcb0xKC4nM0c61veJ6MLFz1DMw2WAp4Lcm/QRu
18wIKeGeY5HqPiGtLGinrTV6j4/fSOpye2zZWXU8bCg+HJC7v+o0aWRpSnCwi5YaO2kimC4tQVL8
MePYknxnzxoTZRCNMcazqgOePBuOt4Ge5PtI4QmtREEvEPskB9hpOSjD17RQvjd7D7HOxr8QbfY5
PSlA8bm4yQw1Na0f1u78O1FXrOaLPJbr50BUC9YdfEcHvrl7Xb3yAOuICQgQKyCpWAkwAFoCNJc+
GqqQgVcVaADU128ff8744b7e0Nx18QnElKId+iiJ++Y4FFJi9Fjerbv9y5GLPg6izD5eVMlv0Bg6
uf0LuU3gjBneosEgTFKmQecqKz5v5C4VvBfu7Q7EkQJTs8iou8cGUv4fovJvauvFM1oEFyrmI/f6
ZoZC5HxV9rdxfJJrp0hftb3LVVbiyDdKmUif7g4273yEGKphnh2fBDV54jmFpIlKUp6PKfpqqs1z
XlDCeDTp1AONwQ7dNliga9ZSJPeoPQIZ61MVZ7AM3lT3wtP5HqLlVSd29y9tLGrFsm4gYwl2LDNA
gUGs4Nk8QkBRtNveFEqaV+hZWpYHnSBs6Ua15XLd682v7v13vxcVYqKt3fVYzv+VVSuTxdmAu7Og
NRLPeDHQxLQ9vqgy2iq86vLYQ2wtitx/+ONxm9YEp/PPh0/8wL+3o2q48z1av5v21xE9pH5mU1M1
Ko7uyfcGGsaywnZN9HAjV/lE64pjLDNZJoGE1JgjreYj6QcaC8hQdzZ/OBYby1Xn5Fk5by/Rpfpz
AXTJaMFv0WMYl1AKuYR8GYBGrFZCm6sDI5xubyXgMF6ZdI71zTuSqoJwteZ77B5HVW0nvjHZjiOC
BdRgCutNfkcEck/YlDMpqlKQVwy1ngHiLcvfeAKkkcWkeh6ieWhzrkR0kLX0p3/pmSNlaSPYfFUr
fGAsz9SrRK5Jfb+i+ST43sPSas4qqMaa6txcDFjt3YdrQZs5eM4bbPALg6gPlcOeTEM4jX2+Yq1g
4yBxMpfbXcqnG7PqyrG5AAzqvOrDzTmFKrvLteJH0Ong7LwRdBaUpuyaMoEvxPvKx1K9igSWxF6e
e/Hh7gTrsELiEI+WNYsMUsHsCK1CFZPN327dikoStuvhFLC5NArG5d6gK9LLknquzd0N0y/iLvAJ
lMRojTNFNZfz93iLe5nmWDZy2qqbo0dxpYl4uYjEXkyIA04Rpdpr7MbbVxF0PF/33kdZizIlTkAA
hTndmbz1DCpWUtOYRGj4cXNr3Lgkj/jZC8/+7SCMYXT78ellWPu2yx2LDD91nzdOAQtWGDuRTBFf
vXBM7hNHqA3X7oBVlFatr1jbMus19MEC7/y8aInvTOriCThoJXNrGG2rSfdnQkHwt7xAL6/xBA35
9RShh3oN2qHMkvhxndpTuPTb6jN+SSk8za+Y7FVNwNOggYMol6J/qbBCRSe0WKVXk9rIigHK48r3
v/mCCDB5T8rKNIJ3zQ0LzLU8NZ1bFNPOcTVGjhVf5hozUrOO4E/joEa1DsaphnAsVUc4C9Z6bd8n
9ePlvcyXVspBpa1dbiZfyck6Xd/nzDe4i1P/EIe/pq/nONhCCkfknYwZMSfhy3v+hk/sh8pLzQoS
Rk0FlkxQ//MLKhec0pm2lY9SlmC7ikeCmG8vNWgHGjskW8Qz0X4WJ7k0xMhZAH4HbR6MeWjURAO8
8eTZT5WdSA+OLLShxSHFyLXmBMKac9TGS/pOFXojGEHzYFp7UT2UEZ4vKoJNIA3j++YxM7h4ENMV
fP95ODofRRc7Y+9pLQKmjNaUAaHjV5DC7h79lvOSk45rbWCt+5TWl4NtHouVOmrQQA+ArOhp4Y3U
eSdRQC+rohUhAIdju3wOqn2Ux1ip8+SSm+wFgXZwZvQXRPa99W0eZSH69As4PK0regivhRTpzRq/
6XL/FU280NGQ9bSoeGII6t6f9LWdLA5I6FISPa4/DlEca9M9fKO4aMUtSOg+FZx8F97T9ceJiac6
qF3mptz2VoL5IHuc8/dRYwapvUiw7PR8gfQMpmVnvzU9ZYqvZpjcUHmwNkNsM0F1Z/leV/e3kgxF
GzKrLcmimHkfZAMYoj/cZufdTCmJPS2VMXSKsIU1bwYj2sOROxYWfeaoukb6INhz9M4fXDEMqTdK
YzdjuYUmbdQ96cjDNGFm20iRbbXDTl8Ed45O5bBUMuoaT2uJhJkFh1mPuLGyXA6IJvP6j4/zHObD
lqFUvWhWKNSrTU9RklUVBypSXbV3UaWwMh1IWgdHfZeUSX+MS4Xxpl21/E050tQGydLXO0I0gRu2
CKE1NExujTbgyrutt7AnoCBzSCXBKSZyZ9LkY++1gL4/b3AMILgs5Zo7QUYz15C8CgEiOchzrSsn
u1Z1utuUNlS11M+59PSgfiM8dzSPyWHtEtv5DZp97XBiHVzgTZLRcclOjS+/QZKDxOfHZhexbPcY
rFR3SpZ8FpYzY+yXmK9gDONmbdOb3VOGMoz+wScRiSlcEJKFjpgBY10G+CSOKyPK1SWEp0q1njTs
9lylNbMmWhjkuJtzZGc91nhe/rn81lMuwvY7p/uJ1Q8nvM7ySyCJzazm0cdeaCsNdC1f4nNXfAg4
GhataUzcNjiB8anyl6Y9O1qfZo2+6oXiMCa7I6xEMTsSdw6sTjzo8bEqLeleK4DfQUq4cUMIQo4c
L/NvqLMnbvGtn32+MrK44wajfKsuZPGt4l5h4nwyjbU4M7UMJ2dNTJLfpOVyPpaBhCr97auMgN9l
DHbuM3b5diFg5bGzIsjH5pI/AW9h3qqDBmUT/CJLTkBHGumkQ3KhhpWLwUKFb8iopWX1kA1t6Ee9
mro+NbGJO2PrfeZljUJ5XIESMg5x1i9tefyM6H0PutFIxNr986u6l2LxW9DQ6+wOr2atR0C8t367
w005SB+IFNzGEzqo9B5l75DPg8GNgdGjN+0oT3dh5pBPpPPWDL8naSrz4NEwUgs2yFF2l+XWRr9N
KGnBxwFnZUvlZuudNCojwYBqHB7mzTLIKWkJAP5x/OjtYoULCRPBzlLuRsjY1mWMgj3VL5lI0Uxy
gL57YQtT5wdHYjNA8Pmny2xpQe+uQdVXFftWYgWmZGNLHgxFK+ean507JeLqQFulAG+L23tIZUXG
2puWTTVSg0emedbX1yqw18sqo4lNLE1AI/Qc8LyI9F2fl79pa5idhj1gzoHlvqnrUa65alAmjnJU
oGpJJDHPlh//IRBEjhdP3DV0TjiMvqfBLihoo9gaW/nVnd6GuW/E2++k5S3PKo2dj16ZKUI1ModI
ZyjlB2a4ALiCB2wQGYk6qWs8wM53kAlGLVS8y6JrHlHeicSNsKZ/kMllpAYY4qsXxXlUlc6QjHk4
EJxUDOtLXOleQEcOiF/twa85JeKc9H/qFWyJWj7MEng7NSdvDswYCGE7U3WzrorD0GnOZzGBzgUe
JNykDqXqkLQR539ccVMpCowF7huG3sM01yLgoMmvI4Pt3MzkvOjIP0FcoQaA1cjyj1mo7f631Ddt
/qSmDOGzAUrLBQT9uslCXfXWTkU+DFzhRd1NgskhcO1Nk82hfIZ8xYxUco3zRdRcds10lq5JAWcg
I9onhxzYvo4UC/sKpxoKMhHxPSWWjee8Wme22UrF1hJ2gWvotU8FFDlWa5npY6Wh6oJ8L+U9ODXb
0Xw7bNkPCNeehq8SzyQhmQJf5WAxZRU5kVrqubLBU6iMDAdxCCcjuuzqsI3AmVauoME3PxBUShK/
GMty/7REdG/xOfkTCpDk5CrY/LemnJHaFZBRq951cn/q57zUos4yA6JEGf4CcVB1PCnkPuME3WUh
wq3OD81rfaGilCBpPyyLKqRx4t9VHd7gPmK4MYyk4rQXnuhzJaFVRWd5iZtfjob0mQQSUYeQMXFr
u6H1g6xXjI2GtHjsFWTSWGqTmFRk8M0H94iS5bY7JQ4rWY6yJTw9JSfFaqPIJJ//bAOKalKQbkwi
p/ZmA2yaEPfgLAvlx6JAyWOVNNiQC0U435Nyy9OA56fMWb2/cHhUffIfx63/M1uA15fH8baFCLuj
RxO9RIEhuBWG92tQKZtUYAA20N5AMfH/ksH8W8LzIy8JUQjAqfCBGpYcyf3Yy398aixEDMbG6IOX
eWJ55jiDgTuiTCQqtw75pZEuMX3YJPdwCrPLZBbF6FcLFtc7uO1vb5zYcFDzn24QkzWCNHUTqgQw
9n0yGZytkjLEvf8BIruzQ6hmu12224QUS2PPfDhPZ0ALMhMq3WcBNwWIT1qWgETyzkTGy0ogAkx4
iCNfIiRr917GQuYv0eMPvsCcgAIhnlCWAsyyN/fEzTvIu65kFF19c9v3ATJk+D3GLn/FkMFHUDjR
/EjeeLyweusu0Nv2PCz7O3Ae8nokkoReniG5OrfASKmLSoP1od2HvaclCkFRBf37nubYW4so2NSx
9Dfg84qaoA+BumGj2VtjnkT0GHreB2PEg988PaF/1lx/qtQ/3ZdAbclw9Cl9Thyd75uXMGgOvUN/
qILwxKgOJzb5D66yuwi0DyzNbOhcpgqqZ7VW6lM77awTjhT7moOzran5sqyTJ2iK3GdGkgMDnsXG
/fBDpHu68Cbxhb6BHMQzX1deiW7bG01HcvgzKIx9PFEkOygC9crtfkc9EQIukDFkHBhQsNOsOaW4
kbDHO2xXgjLQQdfCd5JT1ZZlgIY+FJF+5eF6HafVH2NrX7ldCZnb4BPfXkXGsP1LGxIPUt9zR40M
dAnxO1p9QZ50jIePSYk/ubVRfZ0KvjqPnVPN1P3RAkn6kmk4bYVHtWYc5Orj2N6ap2fOjUg2nEM+
Jh58wS1DNJKGVxP0hAvc0ioHumaowrQkfDHqs8MpSmkAOXSFhwDYdU6b4zl1xoLqVJJrXZqn5o8D
vyVIA10TWG3u/l1CQW8Fct7pvf+8RuufOBS78c8Qdu5vTI5IgdwriQlU6RO4mKbPfP817HO3LNEm
3XZmrrZGRJuDcKP/X2YQzVU+oOnmaR50kZ71rTwZ8tgRmio71rc1iA7OafdEov7Dwfb6nQzVtl+s
BLikcjRL7hYWLgd6x3+KH4lnqgJpi48WE8zuOkdS4A60a8l7EzpegP1I9lbFRzowNeYmjDtU2jGW
5F6iGkCPqcktIDxkaGJwQm/OAZ8nq/kk2Vj7NsFQCEPAckHU5mRZmzBtzSyN4o55A1zTfnrG8DuF
sSSTtJSxk613n4b0igJ3yH27ixwOvYcVLufQGOkGrCruYLGoAP1Xq861KuTmaj5L9MhERQEkRar0
26pPI52+McDznV5UqQwxswTc+f+qO6trmlC5zlq7yHz7G6tAxg/Cf2Ln83omSO2dPJya8DBoYeST
NceyUPR0ghRbs31nOQ+zY7uzg+JoMuH2SW2fUnvpKWhVkR8tUvytVUkbJNn+0fFmo9TcuQ4Bx8Km
+qfFrIVEo8pKJVvq6z0bEmyyJHLMR+ZEmH9Xw2eTka49pKBLRiQoQdBW+YnvOC8vwMzuRehxMysO
1yvlLr85CUB73P2fWRFByUeWkFrJDHaO1ee8QUi/zdxRurogKkik7KMROAL3auUP07nCUp4LtLm6
eR6MqzRROTdNTYXwZqDcgkhswpL5IwbD8l4yVjr6EVHpnOFSt7W9Qy3kf9HMvAcII5eqHkVsDXdQ
z6M6cJ0plSv6fRf/t5h56VoLE2T6dErkYhzbOlbp/UD9V5KPsDoOn53tnV3V98qvQLZhivi52PY7
mHcAlckwMV+TRPlpGnhk/sFxbHBFv0cbrvIKwGu/udMvEMoRWlgkbdGBCosQdZRktOrnO/Q3frfY
/zAl58A2Myf2BiYwTpyMlUOBilOrGlL59KH/FK1BZAiSNxVdop0mU9quyJiUtMULJs9qG8+NxdCi
1DvEqOxtvToqWBgDElyD3a7KkLDY04l4xKU3Lxej/3z2yBeImZsW+IUf6fpmMTua/oKCR5WeIw/x
aILy/fvhY5r1UtEgfbU9TWwPoZrAkWtkc5HKf3ZV9L3f4x+XRR8z44oIu9NSDG2cjI1z9aGK/ry8
c8Yc/75bpSDPnnL5iZBYuuiyGsFkjJwwTnRePa7P8EQ7mBSOV9nrEc7O8qUPMLfotJSNloD/YcII
4w9ivwtLUDM3COIEFCMc041lecLJMmbpdlWvfqiUDPH6QnrIkUFqhDDWORLImxPny4NzvXjgFNnS
tv9QyiTtI8mzPlW65IfWQQItKTHAb0XiTjOPOFkm3Xuilh+yXZu/d2FmVm5nQ080sTiqAZIKhFRF
MMqwKZsZSGhfOrtvkf1V5+eJmnMqU99NS2visEQr2f2pbD3vPFHmB5yv2c0wJhug3mGAWsQfXMhm
ZadgGB6ggJRKlS56dmkOE47Iw3WNdmF6y31l62mUm/yhnd3wwUrVIQEyjreYVyfx7DIEvUgiQXVY
sJ3f2iTwoIxfrqKk/pGpkjtGJIDBLOccAGrg0a8k0naEgm0GdjKYvEyqALv8IcsBZQVwFIIioT/9
llqKt8n3jlVY85Xq9yvMYTOFfVYbhZqbwYyS8ByIuuPD8Qv6T3DqD51ctx1bacXhkPABfXZ1yJ8Q
iuLMQ4bPHOR3atdbKCoQyQvQxxc5m9MyOUL5Y6Cy6LuPDRROTlZBj+0rXypFkEm4RrcMysfEJh0r
lU9Hd2m03Ud/M5nh6bo5lNtAbyst4+6J+w17mZdCbB6l0UWMguzRLADHWxBqUf0x8cuKcvXCTRuR
3u0HMQ4p273kkyK96uc0WrazecMvm/f5PfnY576p3cf9dodm2DQpUSOkSuYUJrOvK0HQIqe2L9Y2
zwVinXvZCuvzs901A1NhUNK1EDEOZLAx1BrjVAB1fSRF04k/wHN8ReQsq65TfXvsovLutP4pPEWz
jT7YqezXmPUP9PcuhskwpSQqrLeiaTE29alTMOzxG844+qbT5ihuzvp6KBPpG3dVvBETBQ6ggeAA
cO0utHNFtHrY3PWNnZNsarDUm1wsV+8k2TpczfxXSfq5RavFjmByX4XdRTEml1+oFo9gJZKvscXt
PY4ZoE/NuZ1Ytu3B6h+NegD247kO1Rvcbpu4HN9tFVeB4+ObOPw/iyopEv2G2PUQ0FrfTQT1u5bi
vXQozcDJw4vIGBP+Z4WXa7JcOOBt+MpPpEYxHbDZhtJtkxrWxAskxUZhDNfbz67PNVD6tj85nR+B
FPz2wraAh56a4msSPEeHrmpq86scS5hdd14to3Rc4nMt6I1ep4+O/U5px7v5YKESgksotLJ8UTGb
ad0PjajeiWPhq5qf9jDFsqJySTkDkyxdUWutJqZG0DWrWjBDnt8O0f1Z/njyr3OE+7yfBw7bAISX
D0a8W7mCtYB4LcnKlfc9A7uVCweAd3keen2QdW2vXoTG42qy2JLoCiYbYS5zS3I2wSOplvBFHKI3
1bGB07xo2+SB1hOa21OTxoOsKXBkXP5kVpIbbh5lMvHwYKEZBZ6QtYLHI4qiYErya+Y0ArAlugYj
C7so515O/rIWqyyEYxQXnpv7lV2+3eWqw3A+8EMqhvQXJ11Fn6EjAvN5J7QWAPZFsoXnvoc05d5Q
EgAfK19dktlXjUnPWGu3Cs+WanxIoYUGUqRi3ib52606FRpq6VhojUC+OMjktdn/MKWuOeg5EHgX
W6PiV+MO5gZm5PW4UliHl3oYexnJfPBWT22DZn0MnJRhhG9EsD1PNlVl2IrPt1aOZHdHEX7kPKMB
dYWH+l+W79rLu3JuSGLNUjMyxa2GQ5qz/kz84MRn4dJhWqlhjEzIhmywOoFjZwtx8GSyczZlDkWn
+WVsnEDqZHWBC6NNpx70sOy+feMBcXDH4dz7Hw2KvPaDldpaV+6vVXAYoGcI2Vtf3Q6+v8F9vda9
448Mku+9JMweAWrmB8yHGDM96vXqiMmRO8dOqHk+fUTusI/5Fx0hRSRqzpo3T1C/45o58zQJyM0o
QakvOvDCUH5YMuudA6vCoIMhB8j8jJ6g+Pp3l/NGB1hj4/7JskE+Z/Kqsa4yd2yL/arLxsCxhKtF
8wEKr4nUZdUGzkAYOOaEkqOtHtQppqnEKUxZ4T+1LROnVFyCam26EO/RqPXUMXRh3XM9UDFzRyyx
hKQpIvn8lp0JR1NHq89etPIkdXF26rwaEQ4u3ckMS+N3ZlkwEOBmonYuS7kxjP2pOXO9MK7ZSfwj
pfVTR3p2FqOvFXY/jV2GU6wLNQyoLSSDVS2xLdAMzdxoy62ma1spChVTjHJWaGXidIIxIt8vlqtR
TBSMyvGlQPusBdaVVjrBv80O4U6UZHyyb4iUpO8n3fKhxexCEyMhhk+ZreOI5Hx2T3/Qel54GH8z
9NKnuXLl8KBhOMSqShgxwNZtE6O5rW52ivVCVczckOdwLfga1Twjynq4Kk0KXjtUN1o5RVwnvUxi
/plKZEefMMa6n8lLeZ5Lunm8ruTK65LcjyGafTdOh/Ef6zWsAc1yDvSGSFd8vy+0QxHMiBlHcAxO
+wBZQZMXqvpUGGZMVj46hUKlpdPKqj/Ej/pzOgODyOw9aCiAx42nkcVQxLDn+TNmji5XuspVhHs4
SssdbCiPKohsBSbbyF7ZnNpbx8sHCMQmNKYxcnaPr5rk70Ep2TyD0xu1SovgsSbyKJLTOuhgCrjJ
hLbSC+cEJT8XMF63bXLD3BZuZ2qrAgAly1QBVNIANLlXxYRs5dhQMZhXeMBuDRTgpDhpE+FYjsjo
VLrtJQuNmS1dErHOKlNu7nTlS/jxqmt09rPfnkexgGXT0VrCPSFMoMqo1H1AHBNmSuvg9SYk9VF4
SFntaeg835AngaQ6+OjHrzRLDeaq1wWeFbFrFg8EfJCmL+dpVOnBOwPLHGvJZEJpA8V7mOOOVoE8
7roq95zrkBqcvijR+CoqOn086s/rq91oq2jXvypZqSlArj6vHixJDo2ztuHV0sg6rWmnUe7g5nvM
4c6+CS6ljgGFTb2p5jfDTICeZ1LhV4woONncqL7pVlX7OLEHIE1m3+5URDMqSsFArQGGd92xYxtL
bWz2Uora5fZfoCL7xbFYzhAhrtSbgnjscPxGjY4XQ3UT2abHBH1kEWexfKYDiUsAEdjwgNJCJ5rJ
Zk4k41xaf4wcQD4I7PnX8k4m3xCDi8jdBi4W3nhtV5Q6n/IfajOnhRgitzeoWT7NdTo2CIRga3ON
kiTeteLR1XdFDwL+BhOVcnWHtFyhYvKP8YV/FFJs3rIhpRTRCFN2SboxmpOoPxfFM4WAjLE4b3ho
Ip4A0Fc7uIOLWTOLbi/bR2cxiO9xY4nv1yCMVxB7OT5wVvEd06RA5sZAliWs2ZX5QEOC1F+2O79U
PAKOtM+MunDI7T92Cm1DBnMz8IrHd1q9bNHzt8Af/GibeAa+rI/Gybm97KSPlxeikZs3KNgUNU/0
DFo1YO+Fbh2n6B8wQ7tgw/Fz8Sm3bMsmeWhIdwf6bXmw9a04+XaLcUHaGhq1N0AWl7hD7PfDBYyY
BkcvHXkGuQMtzFmhB5fgnZua/oGh75JA55BBqV4LdcO2RzDxBc6nLjgv2ROBuU5sbhq1RMYVUH4D
J4qUlkFsSw2nADFc14DY4oDio3vDN9g2PUIiFcr4WteVwmgH+W5E13ID+5HIBZAkq6UTV2b+KEpg
GZc0n7aV/lSB06FRXq/BPnnJrG7WcCL4FLtTgkO2B0xjw4Mge01nwv3kT8V86ZWBPYWtQhVSJsFQ
6XWvUZZbMkPQLssQ0DCCXpA6BH44e4eQh11pog7brvVbEnyvKluWHChzPbGcJNHuNTOG0ozSC5bI
l+DDmncgogyFvW7vcC7xHIU52jnj84k11ms0mAWk2KzupcZPv44IqDGmh+tmd6wrPI53F9SAxNwQ
SqBkThmpZ/0W3gIVQOUbpW/esZzJHtYLhNb3X9YRYa8VYnomvj+Xq8JeHZHbbyGmUIUuL0qapT7J
r2VtVvCizkmPNcptlKXLrQUxjahAPI0YjeoyTLruXFT4G7qtfiR4vnjWxu7ACbWF4uimDP1Oc7tm
tE7sg2eKjzgGY6vK2JF/26i6M+B2GTVSLn+r+J9jCg8cWQbJEPE8kF6eHY36AYx8W1AjbtUEtOKb
XCzoETImd7K7IZ8J31DW/uNM7dFhfMgTfSUeM9SC3dIz48gpHsOFEllFAMcz8A9x7iFomByfPkam
la2KSSWkHk0S6W3vAxk4Bp9tSlfEIOJ+ZO7otOnMcHpwYvWU7rTCs0ezgvR0P1U0fMj7FjeyUE+g
NHu7LoyD2Xomb5hCgLgjfFwQ5Uu/m0yBQm5N9eqtsMeIpdr6B2rYt2rbWXX2S0574IK1I3KzO2wf
Mx/kKtASiBK9F1j1SylcapBQ5oglCwQkIu+xv24YbN7bBXaLRQoTYQjFfssXXVIEQVkuJWRBxSER
39lR+j82OeYLepMxUDX5fNO1Bg2KlG9wbUfjU9ztcn6Tb+XCuQ1AuJshMbzPq+kufc5cazz/CVan
WVSOL1xFJVPAuz6nZXP3JvF5CRfUhEX2KuyRqmMN3+dAGLBdzB7VrOM2LWoOM3mhYWwwEX3vvAD7
J4iVYeTZvBHsiXlFNYFmd3cU2p+0fzfS1E5DD8cIOq/MsdKJOMwf/OoW3cf0er3wn00C1r1LoLy0
R4UXzCntfO+rO+hymwS7wp/GLwfyvui2vre+iEYO8WTH/CyEqzSbs8MT2L5aZpZmA9c2GWKd5BsN
BQnqQ5Q/bFi2aIp2fPz3TiZUy4iolFpYxDg7EjrH7ePSD4VpkilcCB3iPJr6WDnoPrXtGy1vp9sG
+dbAe+H1VjLBpKbcPFiLyA2bQisuTgbIrFqoU2SmuYWuPBeusXHosloY9qR8eiX2GzjpwY1A/4qL
/d5NXTXs8t6TYjQGaLtcagHgWGuvQp9NXm8BOU1mlQ2N8jz/zdqXBaqJPtj1U+6X6RzdsZ8FWb2f
4Fq4xYzH4P5WA5uUX72/DA9t4nYLTuMOL/rFegbF/tm472O+w3kjDJ+arre9cB+b54/nU94fOcYn
AZtCEPkMeKn/Ccoq85gCCx0Gat65su5RsRvboBHnYjAk5+3FtIMhdVr19URs+xXPjtCkDjI1B9Yo
sLFqKRF95K/5t2A6rdAw+a7UdWy9SU9m4nVofmhyZuwlbj7S6eJbnwerAYOsXJoBWK8b+f+LuxaO
N0wDDEvtUDq0NAmPLuQ8A5C7mw2R9x9TROQEEJUnqZkLLpg+jwoZanzlTzFTZ9Qqpd74ipXM4mnx
KeEGdtTY1WhPazbD2AZax4aDCSrxOCMuNysO6y4jxrYDoUXX1be1LvoJe1NIh84rCyqAbKjYhEg8
jz3TFDe8tPoTiajvIgYvQU6zS1TYx5l5omfO91L+L6hUQpBNFPS0ta4ft1yM/3r/py390adm5Hxv
o+cGBAB2ILbYUxpOgzu8aI5FhryJl59qJcKlD0x0b2RN1PcjL+1ee3slEFmMTRSz6j0x3WAZNT/C
jZyjJlufXkKpsibnDoRgYq8IAHjyb9l2dZFdmETJMNEBo6LehJ+QVDxmHM8tf8xx4A9W+WONAl70
BUf1hZqDuFXqN9Yc0nAyCeGWEXAvgDIJipPZAj2K8JNSczGnvgDmn0nQ7s3gLeccIO81oWSR1Ghc
7ywnZB8iALYTyQ2cIrFzcfGI5OGaGhpzM+vtxUEv3KcwdJ7RvnNfCXzagwXuNvarnEazg5/h6ZoY
zaVXir8ynEGnHqSXlIiJgTnpbsESbDxC0Co1uqrD8nMULe8KC5QVZ2Ge2V8XxDp4/YgoPcdknyti
mjauW3alu5+nyUsXJ39HmqY2BGY0Fb6uJ2tgBgDRl5Bh8N902LMj3lp3m6Nb/yZYhEFuFhH2+5cA
DhNmbUWGwRvlUkUU0+yAENib5ErHnyZPPfTM5hFc0AqBrCe8wL5qTwY2OT97Tv21fewbYqzFmn17
oBtCS7R5g+VhguLJw7PV7D8s2FF7dAAM8jlgrrYb7UrXouc+wqwxIXwxZqhmMpaxjcC0gjdAr5Wu
cJlcTDy8s0uTViTk3y3hS2vcG/env+Z0JAqPLp5rb7tKS1WSY0h8sttuhisjZUpS5NDct1kcD1LZ
4fau+YB1s6slfuQKQfdnWeaNQ6XAa9u6xfRCZQIFWavEN13Z3ZTJ7+JGCSuusmC3DLO3RyVcctUu
O0I28Gea8eqHtnojvG1CMnJwIES8iLakYebygemct/fpYXIt82yUC3AhUtZ4sFQcZNWZucDahX8Q
KkiyNqUJgs/kByX8HZ18Fv0IXZuAbEGp0iAvLa16kZBlvqdQflk3vj8NtSYZdhPw5YjrAIb9OGIX
BgTbs75PT8LhG9Hkd1Ba01DQR+z+c0WMzbCqwztPEFgKTIf9i90IvMkIA5qf9uoeOqZRWWGzu2nW
MGjQZAK/XhDHhReQy/HSgefTk2Uvazep3S1gh3erD16uSK3OnHyvqc9t/nHwG8yJWTCnK2PWAhkf
zd9APwv+NdZVPCR6hsK1bt9cATMRdS5gHBG4MdO3bBEZz4y1kdDc7eGqTXizd2R2mb5B2dB0oEq6
WpZ63yQD8RkxT6bLNfbgGqzTltkHTytAgKBNsFaDyqXwbADafLxd4aEqcCcDhXE2xqaTcgD7wgzV
l6E/6WHQt9YnqFo3cmmbMu/mtysVBb0rNe4iQ0ahzEA7WpLbNQD8OidzLeTc6GMaVUyR218+z1Nd
wYPiKM1my01GZtFlwaXqpMVGJv43Um9YqN0DDgLGYFerR0otvNExWmt66CNvAwxBWsQ3J2L+RrzA
PZi3z6xFT2l+xAwdl7n24iq0RjBH9g2aMzLH5K7cvbUAheXOt+9TgHg11YTGIHFkKeO/G7OdGsli
xcYlHxrBy4nydD8Kc0opf8GQMwJl1ogSkmCua7+pAw2rsL9j6WRE6V1iLscq3DcChi6c9DTjI1CW
aOpBXsszSIrktBs/VtqDkDq8wFWC2fx5u8Y70vjAjrwAGAakHODL/OZqYuua9ZsfI6JyLUXwE4Kf
L/EaRfVIIGVBX+v1g+6zgE3+l0hDo+WgVVJL1mR5C3PV/lqMOkcb8K9zsWYdkb718uuTRp+Kr/rh
ZYrSLcabMrZILKaVdKxAK1SUwQ/ttlQYDYVxH7kXKwVQz234H4tPhPAqDxKW5YQss+185OgmXMmy
cp6yvdKzML8mAaW2h40BlOUKazI1XrO7Yv1DkUjSNAU8OXXwFZJ8t1J1GrhjWA+Yl6ZgNLNsqBkq
0rkOqsEUzbReJQEspk0mxPle3WnmfefvUeaVj+W3eJkI/oU87ZZWoc+VRpvFzqtyLmuZj9HAQhwO
a7OOTZBHqFBcXvY7P4UfE9gOjHGFKyliTAvcLcGbWAm7SmjQKYHHbYZXW1vpAMFxf695jhEd0RgA
mqmMVazzagYwSBWUwKqEpCMc4YfFpy0sk3GTmwwW9OnijOC3P9D77XDNusVOSFBie4EiYJmQAhul
8924A5rJdbKeHKqcifxjjcW+fupAhRniVS9EZgWyX+DSlQCFtPgeIEDtnb/IM1oY5ZPPN3myTUMf
RlTX4gSynWnSWuFTnWeNJA4sFdnY8tm0Y4Q8lCs/gcSb+RU4ulD+4BS/gSnnXxWmVOAOSo3XdN7L
pFv7yizlj3NKa19Jfj2nvUQDCp7Zv+hpMeIs8VR34Wm2Xj74xaZ5V5yjLI8NF4kWPo+KqPXnhpnD
7lH4ekhVYIGNInb9A+D2FWMRkw5TgKDQ6q6QfQVkB+MDPUMNq7x7InDnPLanBuX4ChzFvOHRwTQJ
srLiumuz5ppG+QBaBg0vuk/2umvytOjC/5R3n1mJXdMic5bNoNpkYbpIMM/EYDO0KbDrkW+uMvjf
Nv4buxFrxm+Cq1Dev8N7hcZAEZGn9nFPVJcv5Id0DC/Nhb4McUAoUF9GYt/nPAaKyE3/8mGCwsdW
5Xx/mkXLkPj95ALiLxXyjTn2MbeLmd2x1oBn0D0IWPHAwOlQH8Axz+v5y5Eikd/9CqKN9lyv5rc4
s2JZEv6ajf0fsYsGkPf7yc06GJo41GkTX1cQQLCGcNPO42OBt6JPls+LAOL048mJffKlAuKc75tG
a8aqKFpEUpzbWUgysKm+LYTcgMk2z/ZLjIoS3CNn0l1V7IDEoijN/YNRZ4vDeqayoQ1mTvUe/aQ7
1xMH7rXlRvYJ0WOBh02TXTlnidaBiIzZYUOeavn/j0hzY1KYEA/kmtelOtp8o/2UmHK7UNvU4TzR
fALihtmd+k+FM2OGb+byIT05dfC+g+Nj+iU/SKPwBYfY+LkPv1jgKwOnUlVsimYldtfSjt5+ETk9
76sym/CvncexskVtDPzICUSh/BBVv4C2T6uUg5VokDck+isXQmZ/0S8nrNhGNWwRDMh79/yPM9zQ
sgQFJgyIY0lkf29Homr8x/J7jE/anITbAqmtAlfEGN46gU7ePLjFPwObF3n2vMCfjzQD+5++tyJN
3OLaykpYLeUSO+1Sij62lz9Tji2iSSNu38UdFOFEtLEK+gbA+6+14W8RSBf8P6+xxVAZ5FLNb6NN
T/XYABw5keYWY94KYyMY855vmfmbvr3NnuRWqY+a3ejbBJdATnuzX53Pt/G8c17iGv+yncLaTtKC
OHOFRtj976LeKGx5Jqr+HmDFsyj0GRNdBsZci1qIuRfYsb/5vjUCqEaP4yqJePvnxsrr0QbCde2V
9l/mkyfNos2lhiWt6UOPXxH3jPRqUSqDTLtSCvjo5eM4cUnh4FhVvU3V1QSxSWNv0FS1WvnCy7Uu
7Q5FyrZneUflZ+iyjpo47r8wOHdQhJ8jNF8z3DvNoyDr+dNZForej0q9WhqaBCu3W3yzhaX1dsgY
u5cR2wYKXxll9LsV8YgtXDmvNXv0TowIXBl9l2WiQcq/ZqYKxMeap1Yi6aonz3evtG8ni4hk7z5M
NfihgC/tFRDDtbn/2o9vjE90SEud3VJDbFs4HMWThrs9wVV3YV7wLhcJuHtbNfX89mIPtAZCsDLA
eXPjsfauSEYiRAVfpzeYB1Rbbm/Xzepj0KG4ZfCq7svzIW3uYu0XQgoh/fdBynu3unloS+5pmq3M
DkfxV0BYHuca2ItqSfzp5jhGCLowJXvN5GA6JErwMPB4exOTBvCuhO8q7Ussg8SEBayQsVVJV9dZ
/HAKmbpqgxT5ffVoWwsK/76c+arbfbdAAEFgg18boRYhxwtcChyyuz2BZ0w2T48eH/WEq+TXwQSO
gZTD//KYigOQ25iiBE2wlQNzEY5t0LlfE5vgWrpmsIdDSPUKjbXGBFmt4wd/YSmKybh5oCV5uGhT
+ACJ0DhNfv1fLlHPvw/dakro4qKw/JdxPQDLqRyZ0VDDGgkJ+guhmbY46U0E2odEwaDqgeOX2wUD
BrBeCI4vkFGrjOgMJGNpeLwNuWDrXpGjKnUqTVsZBA99e3pDdhUKQovucvvBPml/2myF/dqhZ6UC
MWI+aGiH+VkfE2pwKBFB/n/eJAuQ7VxPSuO1ZnD4ueVO/9f1NdgJOa72bJsY+fnsbWnRn9C9m/Gx
XzRbto7NiOVp4CNt4u7pe/2lYbAt5EGVhchRMAljYMMHkVNJF5dquf3XLkDmvigKmYr0OdtUGzXR
+pQqz0jO2TlGGc2HfnWWSL3XFyZHzb0kNZeasmH8GJPk9SHd2WrVdLcL2iJLUwOUEOsGJDTmbowq
hftln4V0GuyBUwo8o3OmDjwDeOmjL+Rh7j5mYt5JYQwh8q4a/5pQ8YviZmu4yvPMKroSPUNfiAYg
X1T0DDqpLamkIpEGWIx5YWCprBnio5bFliGb6vejx2/uevI/DO8D4mdpuEGwqoQ85o+RPVtB9K1R
eeHWp0di3jIRnwo1CEP0oVsLcVr44RwGbn1YPVbf2B55iHvrxWKefl9BF5Gs+rWbEdZmgJxNpyKb
xXxMAV7VLIh4o6Fpwr+0Jbu/t5yXIxxBLFKDTzJ7tkcrVDpGgqH/6j8Fhq4FT2AAQo2zJJcWGlH+
2Pbhg19d6BrcX7l2/EfqLtoiYieiu2cnFuoVzsmaZKch8b2dZPn6akA+jgUTECn3Fcx5fLRqJuVz
dMknqNQ21YJp1sYcjlfZeylylly/ZbRS/4eJMTWeMwXeheQ7hh24r1uRLXnHAX83XfwCEbUexTiK
bYZTj6EjfNn4hfN/zbMWhdcjyLnzLBWwbsYxJ5mJVi0L6lMckbsi/Z4haBLvJZ7N45QuFxPaFtsO
WCM3kGkrNl0lH9Bi9IqB6u8c9C+G2t4skGRLchJka/kc0Am9VEmFEsIHF4D6AikjUfwjDqTnP3EQ
5cRCeeVugSkn2e51T6sXjcwn3JZWuF2tzoZnAA8jsaXsRx019VRt8vKOnHTI9DQK2XVLp5hlL0fn
jAoOk+hUcx962Vd97ujYftceqQ/HnZVx8Y6fM/8iPrldSuZYuud7CbhKAOzCjfIvfJxkmNPJLLsh
DvYD+0rShgGG/Qr6nZUawjsng0FCZ7crMt4XtBXfCvyKmJrv5Ew9fLHXAImsDtAVRUJpHX5lFZEd
Q3/yMBD0eHr+b6Eua6eai4DN52UpOrWKdxg/5eMQQB1ZSmB35ci1bVAbFMfkhOq8mPkFDNpZfFwo
A4shFE+lzdMBRvJcTelC3O1A19Rscpg1uMuvTUNytk4di5PD2wdXSMEHjnRLB+2UFVncMwL8AkXv
qQP+yPonAo/wLm7kQTkmMhoIQP86tlii610TP92PDzICfYp7gVkha6FVeQneyj7lQFQyK5z81vUc
EFP/DeQyptaooTt83wUIQMBWn1HHXqYIs6B7ByRR0/b+VulMzG2KveLKA/C0GLCUKx6Io0Q4hiC2
e4YZRGOGTcc9B+QlVFRr0DQHuAkY4VNacHyftIHrbNFmnRXl7GuVJ8WLRhFZK+7m8xlea36IFKyt
0nuNkAkFoTmpZQev8taFf0jG+ZEEyVLAvxvP7S4+Pu0eUNrTcpv2j4t3oab+/xenJU8SJpcyjCCN
MyAcCSaReVQxfC6nlLjtniXQcqsaPtYPIhr5O89Mjm3rm6eEX80hGubX8w+mR9aYXcRdwdlXpcLB
OGqi2Ut7C3SGr1vHUif/VCqOk+U2FP1mXrXz2/9m7dVaeid6hDgKr9vFaT7pw9H2/ERWQPS3cqGl
UTd//XWfe/JxJvVFj/PgoLeRfg6bweAY28IRSuzsU8CZRp9uuPBcPtOISQaMbJdYa9H+M06eCmGg
uFPbCv45MFdO6k9XyzQu2AA8DQRTR4c12TCUl8mPNWlxW8oie3x35mjtJv/CiM41pLkAPgLzUx3L
FAlW+xJKoK+/u6kJh/QE+lQFl5wvtErKPS/MmjHOyyZQON96hXBmr+uyGFI9zeJFTyyManD5+PDX
6lJgzIfZMo/u50YQok1y+kdPQ+to7X0U3XmuJtplvcHyqEYoW8jcCGoCYvKNiRqpe7AneZJwwuF1
Y5uia+KQ779uWuspM0LfCZJsOhUHPtuxN/a+a8tf1kZjG1xkcy84FPMsrTobxgE0Da9DBh57qNXG
4AYExiuFPme2xkfGq20fBLOBaSv6kfg1T/g3MnXfcfafuhYgwcWM1SQYVZOaWrGJQtwOy5O5ckZ5
+tQKDEXGwtkg1kuAlSfPC9y3Fg6YshQ//Q/8U13KNCG+sXwKfUt108hXsdC4SrgI8Rmf5CnbA1aV
DCWk5747CLvNFPP/S3QVwRHC4UqMP5DlRShowPJ9CDwtVzqv5Bj3pa0IfqTCEn1QnES7RAE+h3K9
oxo+2Z5fdOYq+jCaaWkpalSvWIfgD5G5ylFfDWoXIA3JDiTANm5rzYGkFm2bKUVJJXoYL2bG5td7
RJ9WFGoWR0rcszNS5Vzhf8xbSZqQKguMfa/+kc4IMrIFowFfKvQuR3eldxCnvfmyHeHVEgmB1eeO
WXo7z2mL3HR+nOQxldqSmyKdG+6gk44y0f7JlEJAjKI7VbP/JSZy50xDXAU/GcE4X3dbQc8QD2TH
J1FkVNyyZCPbjovXuVhqL/pWq9DygcrqPiseszXu92ph9teo+vBZxtl6paC6UxnCDIInp43XYtRa
EQ3eFqdhXEgLW48iCtWfb+2Cb7P1HnWkaL6TUwX6BFW87Je3Gd2GrH9AE45EklRA9ByejB0pJE5b
xtskz3JqXDsTaD2uoGuybVB6CG58nEx7FQ2aGP8QFUMjGnq+o5jFCzBICfYCjCtdz0ezJ6yFjmIK
0RsA9bJjuZpNP7wPyvd5ToKsfzFlp+Otosok040+a4N2eoDn38GdjozBN35UnG4n5Eye5mBz0Qod
6uyrn1b5FRvr3zmunkv57OoNjQJC6E9qUv28AntSKsFvapHtVrOvyVeYRyF+qsIaiX/GL1tgjHwQ
zyPvik2vvsAKILWKFs0a8LUzGcWXVtOys57OsN3AE3VkJeIeikj/ZAYbHW+r1wONg5n76gyb7jpP
DoBzolsH/9Bx1RGSoEwDKrg5A/Kz3wKZUjGeLuqShEmUxSKQpEiX0AStZXc87MNq18yM40q19zYw
6ax6K70ewdstkGUSM+JxfZhOecvX8E3CNyKRNSlSlHKQwy3721io2Pp9F8iMwTf/JIRgDOtInj7w
DKpFRSZJOYTLQXNFdS5r6XFZj/vZwzcx+3zv8jiaZRT7wYQMXEuMSibVjIgHGNASfZVwztR+YDH7
OzFu0QgL8T+kngPBEkDJphqa/reNhY+FRtn46eNH+u4yN0qi1tW9h2gxTUP8hmy4uEOUqaDE9yFg
8myOBGjAbvziDerc3Yupd6m55J60VqBTwo3rYBIKqTJoSkMrxl1IgK2aW7dhUlezyFjwLtphg0q8
fz63RPzZe3KXNuLpjT2DX62KxLlIPpqZ8cZEJNjEb/+TEj6TzBsdUVOkSDrZFLml0h6Qz3arJiM0
iCiA3RxKhs7fZnslzRVsgmYKu8NiC9tdgeXvVPOgKa9NdfEQBG5nljcaf55NqEzwxIr7U1mVDK/V
fd+6e9dlA0WOFqA/Btc96v16GVwfrtEd4ZeRlPrAlKsua7FHwPNL/Y+rs8TI35NjuGXNwpucDiOx
xqo51CkhNQIIQ/WXetaOp/i9C0tQsAj+4I3VttV6cuOg72fD/ROe/PW1qslE5kB5RS96Gck1qR7W
/O22fNdVesWGFv3d93kPOtIQBO7Efj/RI6LZ16HvV6+WQs//gXbkfVbgB7UXUTDS8CMmz7OkRL94
g7Hax6PpWyqDlv6jJvbUHaLWpgiOQog58NOObs2Jg05ZHeY7+aAf4vlM+0P1Ikcct3wFP3OzvD/z
Rz6KhSrpQn+NeBoa6A0D5SppMAas61BMl6hPUs2LZNOqi51GHXQII9e4joj29Tgn1RTAyhWuSsa1
5GEI9JSfMCWsYu+m6O8v8+B+ZzZPEtRjmbzS6RhW0jaN4FVcUZzemVl8Kay4aim/va4YqZvX8gcm
564zSuKQ3bt7uRy22EgsOdFWg8EGBFhyWKF1b8ttC8IsOwKpb/Zi7ZpP8PjGVZIhrggFQ3aCsx1Y
pzagmd0/d+gs+bMccj2ThV1KfluOaNt3vvOmPlQ7f82qhqfC0ySUDPdq0LipZjKoplXpUpjgE1jg
Gz3r5aRd8Ux8uhQjcCk2G6C/uLhl2DcKG3k1faeeLqT7THGbR7sMtWt8Vfkx1A4zloYAkPYPNmUw
Ll3LzwcOtc8Is3AzbufJrG/V6P7NUOQodfqxiUDHLjMZbe5qpo9Zz3RIw//oOJFu8ASMlZSAjAWw
AoJT8ouNMYJ/XeHMk4JowzZdrowUM7UQzfE+uJdX+VCa3EcjFZ1pw0W4DGoduFPqraqg8KqiFNxW
0MCzf9vJ64yipBLe94eAQrgR7Noh4MpQoRpDzHcguRccR4o8XhszsCZ2Fl74qcCXjVJ0TL7SVQ2S
E3AKG2NbgXVR6fwhg24oxIaoaRMOEBczYRj8ZyEZDfCxTIGEBfEBpAs4qmaZcBkeGRI8ndFz/dSm
bfZ068kXVK/Fo4K9Nh/h8FFV4LCyOs6UqlU/NdG5NiQdE0KsVvGdHQnmAxzkwAOfsgS7f3KCk0I6
PEIvX4X9IAJq22wb41x8JiFwlmjTSKrXWJlZvaiYM+W83in5sMe1C7llD7oH55zNByNqtg3G6dY4
Xwd87HV8o3fdR1ZEJR7QAwyUvoUOppyXsWIo7jq96qZqJ2Fg79K+E3v3qBQiuU3V+7T3TrMn0ziX
uM+Vv88VIFyUEHRSyFa0H/dAnlqjZULohkLXo0F3V4Yw5/EOjSf8nkiSbI3jRXJMcm6iy/aG120S
z9J72MsTMt6BOwCYJvSgBLnrnTX/cowu8Z97ZstX0Qsot9FfWG0qJkSQePPGmZcK2LW6jXNEh+zR
ajfm0RbsUaz9DI32LrkoiS+602mgYBxaM2RnJVS8lVa41FJA0Zzt01LNuBX70/l6/1prreuuv2OB
/qaftz3LaCS08uE5jMLjW7sZtUPUFPjYJCR7B+f/0IjWrG+xk6AXYL1SboppEdt2fcnXUd7HVJnW
v2J+LBZOxTooheE1sLCOZHWQbxKbLW8eyRhaUp5F4Ch8uI2MWJwmKq9g6CJHlFp//qEoCS1paZZE
UEbzcCs8o6dDkuIz/v6iNrEUQ9wWYfGAapmb4RVgJPgeI5fAgZhKtQ+rrrrSDMlungOhO+1iLpPj
DqW1ZkgMrkxNx1rFpHDbbN7fjxFhqm4F7JJtfRdckJ+DFIJ0bOaPPvGIiL6cshvjErVX1ah8phxw
p6w9Y8Hg2hTmVU+TFp74uwzKjLdNMju0rOg6i5nOD39EYnLmgl0xmEElhxv0EkX0x/vEtsi4SD/V
saEgF22FiLojP4Wu60q3rUAIRz3DVQNZyITSCUwg3jyFZZA0NPr6sTJ0o8GOnUFf0XQSlGqjlRFV
qb8T4vly0mi92RXIPy+yqGgBQfba0sVfVBlnCiD2mTIxpGaK1dqJseQSr5r4WoYqEBoTTyCSdwsM
smDJNr60T5/sbkxFvm1tFQ65WjLgzz/bG5cAiHmrf+joKKrgs93jIZwEdoe4uEZ0U3szJg2v6hW5
bcTFzmgHKXW4yMPm93XVbRr357t9aWtpvVBGm8KLE5yLN09ngvHjePPg8Mo8ZKjqbPBBYQbMkoxI
1o87XURdfTBbAWEakyh4aqUD+i2KjFDxW1+XQnVTJP1sZStkwE8oZUekXF2wK3k1RTiGTSORC4OM
7jqRruTv25+EonoqgVRlJosy4LJxuy2upr0NC3CPO/RO7uzKXO+3m1/f8mMgeUOuNXuOk8JQsBi5
9k6fQsfoJkmwOL3wGZsKRR5QATqnlHPqFJCVJqbKMhtZvgVX+saq4+nkUD9hhDl2LrCKUkA+U5qy
mY6Y/uQvhSyPYKbEaPDp6IewXSx5H7RN2cV+LbqDvunJwZOld7msJxVs7Z0br0lCizRi1EcAztB0
c4VkHMKHnm3ZJZWxksYtt/XsQqKw2aZtebyYSsNYPCb9+2fdrMg4ydFr5H++vPURZ7OAT8rEr0zQ
lXIWEnWQ6yYXkPAgPbPOIufyWu4hRxuCBW+L/XBQdezUwCsbITZseWfvlFN2fvLc9CDonebTq0E4
IoW4nx0z+kexuCVA/aQY109UqXUGfNGrz6Drs4oDE2JzQ3MqvmbpnOEPm6rwW21Q/vJca8sy3ebD
aEMrcapWRNQ493HiZhrKS6PVkU7jgIrcL8OCb/mFhScw8K3Fuz+RqQRbV0sueU1IQoEv2ji/5ha+
IjhcMhA01Sc4jUwauyY461FL1MxI3SCseh8nFeLcvEq6MT9i9MiYK1+3owSI/7cP5Q+XOEP126Ek
THTyltalkqdcgg1/Rd9iG2lTugKewVk2Wlod6XLjx4/UkrZasZSJ0e8c0H9C3Cop8/4sHAQW4Hx1
t7T45cRn+5UY5X+QXOitj29nmH471taLrncMBX2KRHjfcU2KDfjoa/xb55+bXw2mie0ywGX8dOjK
lQtf2a1nVJ9bOxT5IrZADi6ZnSK/PEvuaFrupo7SUNEshC5L4zkZpKkFXmhSz2vLvlQrna5P+vcx
EzFlbqihURFy3AKWNN8MI4wPpHEr7Q59Cj36rjP3So8gS5ED3gBxN9TPPqwD+Jx08S5Y4l4JXzIe
r4lOb6DeWu2WOsQAXJpQFUbNdmOm0o/oEnP2qZdS76pMMriluB7gnNg1AXQd9OMtytQXBZWDUMYc
5nXqJUGmDE3vOSMSHCT2ofjQwResLbP00sLysZCljs9ViEMyOR6CnV4pc3+bOwyODMejLbTR0GM8
givJ5Z2uJeHMEE+/x7dPg4KU9a8+YayapExUThNS5BE6V58Mtl74L3Sqw+T/ilySFIFWtFXq9AZZ
EueaxlXvPZByLsiPMhJ4TXFctv5Uc+D7CaXbPIrRuCwdhqzoPDchNXu3bU2vGSNYeiSNvIHsjino
Nmj/pWCs7n1lmsZRaT1KuerkeQWQxkU3aDtaf+rQZRe6Rbh8JVPTqk3p/HTeGe4BrDUitv1W3XiP
YXinehy0o0t+Gh9QXFECIT3B9Isgqm6Bi1akTpq3TTNxCxHEIOfe6xSJikuhFAeKdBfCHmMnA5sa
Up8pIywWB7rHdQ1lRQKr/ulSTZ1CzRqBe55nx0rNcqwGm/iUZGEwq7ntVovyw0EQ57y6K/nLMrcf
Vn+8qp4aZgkSuF0EFQbzesmGrROanoR9rfluv8zFN0fJHV1zJdnYI/6O53y2ISr0zHTOvONRIw2j
KpU+djPolLcoKg9q5pyaPYFuuDjPvoCWMGW+H3U3T7pOMvosOncUqouJmKj5/dcg+7yW0jDJXBlF
HVBKUsV4g/xVD87S9chbL2TvT9kNkMKAUSf1XZOoAaVZYg7H91kQxVOwmkruJOi+7M3Et4LPYCVa
DVfgXteT2Kd+I2sFNkuzWuAq646dDZHLRbHfQ5BGAD1qexS5HdYlxMCjMUQht3bcrhrLyrvDLRdM
Ljjq0qmgEF/oV/SPbMnYJldRB5TrrRWU9Lqdll4sdvmU3Vl7UC8lHlP2ZV+2eW9cqMqOBKrIvjwK
0GAJIF8PfofmleVJoAm8scaTwN/nruKF0QrcVNEoFZ0DBNDlfXY3SfKsoZvIywypEeQFnDoTPmkA
6t9ZHmrwbnwUwZBZEDL9ZRIfM7EnnKeHQih3ktHkt1KAw/w2zUXomIHyk0FpAIEtbL6VU3CUMXZX
sYkoZyBbfvJJHvCagwz7MFt4H9eeatkqLT5Hgpi9WLeUTE9tvaO1i9NIRIj7xFsX3VNXKTFd4xf+
4VCsrH/IQfCtZZ+YjHKHBQMs0NunaEKeoKxqUy8osD7TvWeaPk1IJeT53DKrYZZ/jsgDz3pBnKI2
ShbOt8LRJCJoPcIgtDyFZDugEMHo99YxfA5kdOXMccwM1uQcmnJEzr+OfbbK36GPY2EdY592lQOD
UIxYPrWFoj9n//NPIxqnLuuF0UKDF8+w8hJzfi4qSxQP0d8HoR0OSQF2lLYXqBgROO44oP+GObH+
LZsNvBeQBBcvBK3TsESw4CuqC3Xt5v0gwtlOhjXEjLELbanO113UFDnMznlLYYjndTwNF+RaGqpF
OZNlbAwpcZWHKhmTaJntGjAoccMI6CQTEsnL3JEo5D2copzw5XZYOBzSDHMhL8bmQxvd1L5988jV
FYvEYvTekGR9pTEZbKUw82Cubfk5tWf2pn8l4Z6hZwlmhG/QwGxvvvEg9iY19TJDYjHmefh8c7aN
Q53dUKGuj7+FvoBnjVSBiDHnnoN6zGAIYc5VhUXooLrdLcveVJOT+yexBhPpgNTooBpljYD0fk/v
TcKL3m2kHOlxMI+aD3TWIr1/ZqZrch20YrdPQsemNeDaRg4kIEAVlwL0owVyp8GHPp3V1xsvRBuw
Btr42CFfQXLx2sIygdGh8ia48GAU+a6pbXKfBDht5bxEHKOncs+43jubl2N3ScE3ywodfls3D+fz
Nh8+uxr83F6k2meSmvO7s9+vp0pWxzyHavyPKT1c/MWMhfMm7W+oJfaoUEDvTLjSCy49sQrGIMxt
EpE3V8Fc43pqQwTJFTe2iDMeP6I3ZYmwPJXGrERGhDl9flhxbgw2nhLW3kOFnplUfgVQsoGWFZXV
/9+AXBM/zHE26ZYKDbIQNQBrY6OiBCNci0tKN+igex/Mkp6Aknqhx8KRG+SGGHT9j1qKopu1Mc8w
XnQQ0yUvlv26MCtE9yej0IOLZI/+LPyAAQrn3PKjubRfnx9IhYyCYKY7j/J/OtEmd/4lz1w65H7V
JcxbFgNkyAbQrcFx57GkbiPUjttacTzP5teSNg9MqRVRD+PGStx6MJ+fVpvjfp/C7gYboSjpx5vp
FJcUc1ynfOYn/nxm5mcQYg9oSEKII6SyQPxG3X9RqzQXdAstUuVSLPJ+ZzSGOgAmJ27ymugLgg9Q
EKH4EUUyZcha/O0KgTTKxW3i9lcRSofMQgMeVszr8/1KzBZtDdD3iUd+IR2MA5E93YbazpNbkyVb
o1PSioX9COnQ/+w++bhfxU4oxetpktDJpl8b5F+F8lNw2b14HgFtNDH0HpNN8ik9Lna5QnAvscZA
oIxpjxmBGxN4XZWKG6p5vUfl5y6nXfpzUqXbW1nnilNcowtfV/U6utJ5Pcda52Xo75wAsjhKcQ5v
tS2756uwZKERi3503Nk+VO/8DGINjSGIbqHdgWLxZNOaxzaTNFadQtZTHSl9LZProLEkKUM4tYix
w5RJy20wknHbOaVvs+5GL78AFlKlBjkPy0AMA+3Vjs3pJ0wgQMKiMGYgWykIoNq8IXjNn6gN74XN
f6Crp4KR4oYoh0epjNQa/11HFt2WAveVjXwXH0Mm8E97lD+vyoh72qJ/LtFaWKmHI490vNQ6F1vy
5N0itm9rMhH4+Lg7CZV4+dvdc3VdJZBbPYKAHZsox1JA4BZ2/WkyoECBQNf8YgdNK5VKUyEykiW0
IGMiQbmjnhgZ10W9mnpIryPCoT8uMb7fZInuFfbOBU5ifGPAwimhHfG4Nd5VeufiSgjTCuCW+8sS
Cvp3lB5pKTSTKNMakGeS3yqJE5RuBjo96FNpjPP4P6dcia+A2Iva5WrMdGUplwdmzWaSJ/pxmDOs
9yyEeBBita3eMIqtm03DwPbkFb3Nc5cV2UK8airYMc7jkMhOrIkcWMCBtbwiEcwKuv6hSV3TC2DX
AuHDbfk1y0vIzN2kZIH5ud2MD2wo26mKG4RXjvBvoA+K4CC+ztn7U3+rA5Ps7UbImxRLpBFhtuSx
usJo5KxJY4gDgwhCVDVSnbOR7oi/xZ1vlikdmGvl594hoeQXljqYtrwIMBf8j53+XSnLid06k8tj
rsJFAaAMbF3DNj3pPd+r6/BRjr/s2o0wAzlRGjiWZtkILzUZR7Ofd8jCkAmPcUOxliv7iQZMjziF
kx3wlHnAcYU8RCQnIh8jbRZ2NLX3FDcodYgxa3P2u4MUULUiBt6x2tfyNzxX7O1NT9l6T/gERBiF
EIIBIW0ymCFrmq6Fl3XL0FjhLgoQzCF7UNSpoG+Jkpy5KQJDFO6Q6X6J4BYlPlfUwN8JWRW0agkt
kuLWlcLadbEoo3rUAnt+qNbWxv6e2qZg3HMRhMV8lYZXyGUWwKgbptk03x+IKT2lb5hG64Q9rj+9
mUNzVYGN69HyVBhKNfFx8H3MQCJlfBhmHMR5xaKdIrplHw36zXRIo5AjkipgPb8CCJ8shFEMhLVh
8BJ5PoZh6BeS5CO69uVxa+/Spw0RSY/NzvizdYIU5cayM/RM50VZLlO04+m6jyW3G/dqLrpw+5gc
6ehIudWy9FxggDKrmlUJa0RI5KTy7xo6ckhuZtPju1mtpDXYVVgmQTb/8wY7kzVr5y3Z7Fl0mILF
mY7vBmUFWqR5jcq0qQDMD9zpQuro8Z1ZHG+htalP1L053gUpz4kg9T26OZHokZhoHNpnZWFoS3J4
SQBch3EmjJX508xUVNv6vEac0lCvlaeDaTfj2e96U/MZvY+DtBP4Ae5emphlmiQifZEXUhum6BtZ
PWX0F+XkmkWR34pL492lXArTepVfbKMUZsORlNWTa25aZvZvmPJ2XtFpaOHPpCg1AZb4kW0m1OCz
ky/u/tzECCz9omfDMmeMB8U3WHxNuV8dd1bakQUaykCe3NJ63B6f635UegHwfJOCwwxeXYuLn/Oy
G8CA0dfvbQmXy2sgsoqUekpT+VIj3MD6zswVOhv3oPhec82sSj5oJjJrp4HiPVY+o856jHvEvexN
jgt1lnHqmJ8qp3YR1uzzNLHOhIzVOiy6B0F3jG8XxeS/kkL7vgC90zCnzxB4UHze91Wh9YF/jkvt
Wh1yR24Iz3FdgieCc09LW1D95nuw8WcS26/N+6Aewi0G6fm62msixUxnuFy08DQZDW4dO7uEYvns
haKuoh5aq1y0Qb5GMG9RXuCgGpP73OMz7W1Wwh/j11PUtYfvXFHNIEeO2PAS+pwO8eA6f4cxG8U6
aywBgFisOyFQ/KWJP+chPrpQkzvc5KtsHsZIyZabtWv0lJmV/KG22IUYc3B0wSBn57HXQJA7Q8yS
M+IlUF/8NKJxd0SXJ3yhYE86XmOWZEWJXSZfTGVHJq1K1K74Op7Lty2EVQwYHcrKPEuhICMDiqiu
jqrv0oS68ry0Sm/0ryLC05LldVZpuQXLj1ZIYikDqZTRpFMSBF/+c4prWn1DpHWoA4vKLW8nE7Ci
3XGgp6S9LzgOtgVjtn09czFJL5kwsrv+/IWhaJ4biQHSvM9bgTW5GLNphvvqY4LvuNDt5sB8njV/
kdayk5J95cNN+/bXGL0cwOGgTDzV64Tj7zOFHqoOaSYLmXA08W4vWYlNVI2/KrErGlzUzsyPEHKh
NCbErTjoSQQs0L9KnTBT7kjH8cz13h+IzeAfqRGgN3X14ZY1ksUxDraidru6dMrr/F1OMbV9MFUj
zUReN87ZY8zBE16sEOsIsrhmXFK9j8/1RAQyyHbfyBUfVNQ/7+Bt4gzXzxfJZE922+ntONYiaGOw
Oct5A8urxrmuqj/ulYjkDPUpOL1bj/QM1el9WkPEW9j6O0VRMd/A/fq0kfASi1I4EZeYorvhpgCm
JZnI5oebF4iiJcoKEy6O+hnL8bKd1EWqzS9U9xAsCkTXPh/xeOOOVRTdiCAkSGE5XhJ3SN9TxKZd
Xc5TIZQ+tjHBw3BU6LeLz2GJxSNqr7g2hMPnvLvftE1F6zbxzZqwacfNBWDScxjLaP+jI6mGS2rD
mtPbd8WvAqgpIY2ZNrKK/NQgaAEKG6SMGCyidyGMVfuIgZeQjHEIjrAtEwOCo7lKGSWA2g7TcKzn
GLeUO7ezpDWQl8x3yz3y36UZCJ9pJzLm79aFK6zDaYJY7w3qxJ/JJxal1qGohFXolhMhzrTu02CJ
kA5AIaxUKaU0qtj0SAicxy8yiNdixa80faHEiOXtlXXD2DlcKP0Hu8sBIuO2x3BJN9yQnZtBlYxk
74yqhAxp7ZnL2kfB9Js+Chwnv2acK9KOU4t8m8rkvcvRuQPbSUo0YMm4WJD4P9bq3tGp4+EAJsmZ
3Jta2QKJ33uQac5mBOaZzUgehpvrBaJVeVj3r3+6/px/0CpAhdmYeDKhQD46gh4P6hIBVuZYosvI
UV7NQV/APDIGhRx9wqLvmoEbQvbdWUbsqLhb/QM6qYHLjBnI1MNpLtWvCsgUy9RdSxL32TulL/La
WZWgg/wKV5R7aeyFUsdbsLC8KS/ft0PhdxV0M9XiwiSulAuQv1OTHNUEoIoRIz9smHZjZJZodkL6
3VGzVsY4FXmtTgDXXeocG7aqUC9KGwJ/qSWOC6NZsik7ORVpId5/7q62VnfPAY4h8EQ5fyg1scIw
7UirVDxoH7feL7Fsa83kX1iPGCUkHmNNGbzveUeKBMUNoKNgQ1Zp4amF8jf0VZKfW7ixynJ/rNzI
cY4jFkWzlT3yvsRFGs0b8dT7HJeCDMyn2kgOdeeIVa6GoLrG32AILcI4/J19GT1iAwYObJP3wX/J
nPA4SHu8/7cgKKr4WwazHNBfsGfaUYMsI5R+0+O101ToJnr0yoTDD4HEoN2EUA8gpFrecF2zyVeE
tyIkhqoE93bsO1bNa4HSRmWGAeoI928DtLbLy71oVvidPlP8oFjd6PLAnAoblVALVU5bFP4zNC3q
JNcmXiYqPBJUCGUztJkCPkznYJIQwzQFxzg3Lgxm1aBHOkqmBeyHrHUN3OvTtarT5yECjCCZC46E
Q8QMbuRZS+0j6JBzfio0t3PEGnHMXvCNjHgqkMZKw3VZUUYHn3MzRgtHgPJ0jJqrnlP+/Kavi8PK
zulC2JFlH6dtYd4W+FOuPbp9qmPv34E7MdZH1YKWQqa5etJi4qPy4mThB6nuY4A822vCnCdB8xNQ
9pmWNdMqrfNoFWrRv6jKb2f2L8Ixm8GvMDYXXFTLjysjtpOqq4JJEOyfQsKGiNyM45R3NpNR91XS
WDYLdY4t5r/ugZgmg/G4E+2g4tQ+eYLc+6nqyHZbeM7mdzmBRfUfa/pHHzttAPyLlpNMjuvXLHgU
AU4ReSWoDCUjTnsI20ZLxXJ56jKwbhjlsfZTEVn/884bCtp3XQfJtthEHDT6xGoZjleQwlZ++7eS
OoMFj7EddWtKBRVfRrJo/tnogzH73gO2z8l6+CVagUIUPaGCSva0E2G+hk24qt7OpsvzAUlKqhp8
fZZ4HeDtjgfSu4LGJABvFG0vsrqwR+gpQnY4Bt34jamnKgX3dgx8uL1fSYlBi1NT208ThWPZFwiY
sWQqUAt23fz14gm2sqCl91yqaup9M69Qc7n2WAWJR5sVGXLzmJq1Y66gIov6yEp0XRGKX3YQ288g
sg6s+iQVrYrb5DJ4z2xQI/TmORiH42zdSep0dX/tyjoLMJEkrbeUfmMjlhZGSakwnAi9UOcSvB2f
F3Qvg3FpzszhknHNz5OOAzkJUhCdz6JEojeCOZClxZoxBInP+tV2T8s3Vq04ct6N3v6Ezdgj2pyu
g+xm3gBGSgFvysrnPg2fNxP70/ZrDHOqJLt6y8T0V1Op+U4vBtARAjkt4Yjdc6/2ZU8pNOeBwZuL
vm3JMFdMR1xAU6IJ35oXuMpt3tK24DENR0h/zJZSuzHQVns7e+H+y5ikync/+JvVLlnjuFm1FGJH
9RZtQ0qlI1Ep/dEyVoyOkk8+trjcpQdUktytAf0fvjiZJ8UFwVUwwN63PpToQwgOTV2cCEW6tHqt
HNxHrv2D4K9oU1LKJ/Fsor9NHy9x2cBg3CPgZOIPP9apvN52P2Nx8LKV9abRGmXlEiXsn5a09jgj
Skh3RMCwdmLcMMreOFdf7KAQEwb52rOaelBG8E043iS3sfKzC3UKaZGgbXybPgR+jjI6dIm6+m/G
CPigr2hVv06fPeVsSAPMCgtN+csGukcN+OOvpUcbp9XFw+qFHx1HMRSTO86qHAG1BLl4BkBd6tmO
gGNyiMAgwz82rOuf3NY2svA/yfur1NTFZnybgXc9rDqWFiF5vFwQRtd4m/GDpYqQJshdGmAuhfDU
ErDzqMmQhaJyizuBmf/JoiasbLg0sWxb7v8QpE8eo+uvQ9x7StYjBQzUGZsE0JAZ9MtEybT1wOt8
gI6DpCuZSYc5WPEEkGOHJg9KzBhb87yAMNNYlST4/JQrqWF6TYf13JnO5EhnNiBjc6AUK85zwBNf
taGbCVDMmvTE227rQcGOWZKLGvzh2fJq8xXe56PfdbRdXLP0KTXeThkGD9ww3xK3bPCZC5tuK+F0
o6gR0qEWj4+nhxMAQpcss4H384X+vYQu3XIVRMGZB9yPvpIBAJcv7vpI2qiVZw7hHksNOCKJzvBV
ZzJ0edAI0UHHlwvr0AfDOR12ceyf21FT54ewDqmXQw69bni6thruBbs2pYmYAyMAtk5N9LwCxrKe
k8hAMnrAjNy6MwqI5/JqAZJshdpIOcQzqCnwCTBaoiDBfbc6zb1mocobQOec0HzzSOlv3OZQVvjP
PgGpgkby/x9zzp0gYXBDyYWOjIIdssxDz3Eci/icjg2mVCXEjq02G7HCwp07D8MTX3BNWXCDS4u7
yrPHHgbh5F9Cs2KlqbpZ4JKhkDrgvppIS02x0n84oRzL4Sq00mwkqADfkomjxP0Yp8B59qylBEwd
hPQoI6G9TBZm5wPzvuhxYHsOiK0SiUqvk0KUJg6rgwz0IiuFQdT0g+EgUo4QXIAfvTQgFe/ksQX4
rHp1nMFyd0DoiIvIux4Vs55TqfTZzzp27QFZcvzVJ5RQ2kxV+7iMw67Fa9ygm0+5m6XyRoQQlP3P
gL5unTB4x+sDjEXsoJNIQyq6NILTaQSNeZsUkkmyqIqaW1LC+YP8qGuUlr9tCDG+4Rf7YjTcOlZW
/iga1+/xh9YNm41rYQGb6ZQRyVZPfngBrlBO6i0FdFoPQ60smhiv0gSoHtXNCMJEG4wy5tWkePnV
wy7405PR8scRvYzhacSpBH/uzUuR6OnamYAf5UOPoyP7xilOphla/yPgKkuqHolfj7/xfDVqDDkG
/eZQoYb7emV4HPpng0a6U/aT7dt72A7+XNGEkDL0BB1pEc3+zjohS2VB/2SQYOFXPBhnaLmZsrV8
bXrzIX3uzBDZJu4JsDJ5LhSXFlZ/S+IIOBVmwfSorBWl/ZbuWQAZgruYffBVOZc8xOLaZwC9XolN
wRy3eKM63hW2UXLi3YspnXLrr9If0qTG+Dip6xizZEbmzBSsLrltWXb1J1/6UQXZpUF8v1f2quVz
jD7ipLZjOQldhzVv2bNn8aodzabmPQZXl9Ibjp2GBtUPtKKqeknzRSdToSylvb+7Qzn/q9nqcM+B
02E6ZKKa19As2wbKYj+04dgsEoC75ER4MVqL9dlD6dKHXAOSk624LZCiFSBEbEkGC/T90Rf+1KFP
l/1jcsM+TRemFR6G6PKl4a2GK51yJJU8ae+qmBFSufrMfCtzhv8gV+JW5IRaQIG49MTIMbi0jhvo
dvz+xSe6XIUtdpkNRr/T5FxES1yeO2fYep841PglTpGTNzCDAk7K49YQVZAyMG3zJnjkytm6pTXs
fuHRkGFJa54V11KyZnhFt4JedrAsO0nY8zZ4htkqkdDH9nlDIxV/ZMYt3cVgdFEdbBQUa9r42cD/
X5ias9v5U2cB/3gcWwljtTL0G4I5qtPbd3MrzX6uSurdqPSRNA5hFD9b05B6K6YXZoSs/fpqRVMa
2/EVbcRJ3NCnL0fhCoXG4ojDLlTFNd9559c4c3LrevC8qJ/o3V0lL+7i1bpB3jWI16L+Nz1dZCMR
OWdpxHO+5D/cI1Xor3OVOmHVMYayPf8MXfzISnsTnuwpMkP+5a/DV2saCYzJmBye31FaLwjfUOHS
l7EZssC6dT5Z0z6Wig1iA1y9kowDJBDAic0oG78/mr2Zk6Cjd+h92rgTuf00dtTaIxIykSjtmZtE
jZPaVoO8NGURz0UIOa+NTJP+cDXdg5mb06Z3sL/jVLkgm+ItAyFpXg02CO5BaOQtv2o78dasE5/n
0o9qE0NweCLDMDW5anhELd80xW1Lp6Z1HZW7Y5wNAfYcFBj21bIdkLdxLF5QWrp0oqZxvjjYOjk4
+mMwbz/QHXDg11POMJfZTY0OqLcgHl9dJyyPaTjASf7F0VXR2Fw1PCu084HKOkqVcU3wwm+aWd5n
gV7yKbmcv2ybEMFVx0IjBfTHOqXDxx6udIyvaxFYIrvY7t/jQeQ0NuxTqn8I6lx9nrFt6o5miAt3
sJg7iqRufxjvyL4uIuCb01MAq6pLC7TC2aGtBWQ9dou7mqTDCyIJpcT3dIGeCRz6VbRkC6j0/yIj
R3cz9L7E41w+nkYX5Q+Nzmpiyigk5pg4VTALgyUtoeDKfHXkjs71c0To/4u5wQg7at8+0TZe2Xhw
gVZMj2Ggag8bxMQz1UdDLeXA2XJ4uNhj3f+41zGct70vbgit0H56gQpMALdO+6FjnkXo44nSd35I
XoipCeZg7QRep1Ez0dZ69yKo5reQ/j+3I5ThYgTVgNqEY4y1K8EQKYKeFrVihkDhyH5yyWDxAo6X
HMeEWjT4WIMia8XgeeBaYgjCDrndKKiApu9LL4kBqJYxcPLQgDsXhKs0N28217Sqj3SQQy8geWeo
B6Y7A+JtOFoCxr2ap4mz5nBH3f2zs2+2V1SMvCBJe3/NZXgRI9Xvijq8ka8S8K/YForG9duVFH9C
EWehUNyJwJPzwB39GHr8+v0I7k4btax6cw4YAKGJBqcrAHWdEcU9rpGzU7I5QDWGQf8+yiqJe9iA
8fE7Bq27JpAGyjAnmJZK++QMhW/UmgtQTkqKUSSE7eaEwp/sLIMzOs89kdYM7fiu7UL0SGMbgl9x
sSQ1OQNpYR617r/v9tO+ys+4n9wuyik8PcMCBf/9xujkKJf+ax9YxB6ivUmYNFsoUKhqP3/UydIR
FgZcVZZ36MJNubSbuz1cJds1no3CFlg56cacXj9k9798+MukM4qhb5JkP2l4c1/9ut9LIfHTIlQU
IEYl88sGmKT/R/yhxsmr01ptE3o2D5NJv6QpbEDEH5ZQCnbYnWmsgVtq8ZjYmM89eM+/QqWHR41o
mS4LDQRn42aU9b0hMZqBkSNv27Y2yRMjzBrXglyfXUnxzXcShWQhQV02B6oesqv6BR9gfsfAuH+a
ZUctIvqf7GL5G0CRGS79BkQdMEWUq2YDjbM3Qq+RmRpsf7fEPtycKst1O29DBTcZJGLOPKc9mVYd
P+ZGx6jR0O1+ol9ZesoJIz+wPeZs2trKgcpDWUtItMF97Eg+RUIXXfqMXuOsbUWxIkqszOo6Tgqx
gviZxl6I1z8LQgyw71rRST7FuqkfnxgTE/wUuBt4PdE00D2WDNofzin+qpl2Awgy4ROWjNQ+RfCZ
CH19L8ZgzWQb21FmdIfBI2jO0FCa0rHmDrhrofidPjBovlWQYt/lwftsN4+nS//h1AbIB+D24WvL
3gfqsV6/l5QsUhuJqfgu2ZFhOkr8vI5ptAkYSOuX1ypsiEe/xteNeV8BmCt2Ljy/1/ob7PUvmvNs
yMr8L4UAg3MUxBBcV6D9MTfOBMcJ8D7eiIuJLi2vf7Ii6X5ZS2e0HLd+Vy9T9Og4mZTFmOnXUtNt
KC+RNW/jIvTp0zppPqtSETPg3VLEX3h/6Qe7J8j+QAMVxEGAMpRYXkX9VMfeLnHVtlKV/huQjQGz
qI5zXdGxaf6kPEAWtD1Ae7E104sz0MVavKVkhbd0gTsJCGj5PnlskrZf6CI79Gc9hsGQpO6hud8Y
bryc0aukaoSJjw1WIh4e0Ej7jwTc7+3I2S+rT5oLysGol80Ts+eshMxTszpPP910O7o1dl2/T/S7
xCrJf8Bqc4le0Yafr0GnOBBs31EjsACOIexwPtcW2IJa9uhNgRnNDHMhV8e4g5x5TGoNyTpAKe4U
7U0QFORK3cWY7RLzzDWhcQKJUpI7JqVRAKKWp5wf5TbeMOfzk49KrmoXW9Kk6rsYF4rg7ZFzT/U4
hqARz8j0YrYEQ3aiBuUZbm5D5CC03xlsLKJmTt6waPW/h8alJLlaM+zfl9KfWjzYxoiBkRksa/Il
4FMI+JDpdK7fZg6OHrqUi5+4ZhsCXURbIpovw61NN1x+fiRoeP6TddaWsuG5NAXXvAP/GqAT0nrC
3DziUGL3OeK1kKXb9FE2TRoJOvgh5zvsYH68CjORVWtYJwlGG5T/QXZR/Xl63D/wmYE2I6HaECnt
qV/AZNVHD/vY+xTOmW0BKhQpWhHsSngdQXuHMLqS91GqPfrA/wpjU16MSBNlgVDu6y25BUsDM79t
4QdpAZPOKVAsg6zOXRHfKRBnl+pJ8B3qx7YOUPfQjiKZBtQqbOTv+afHAlDFwURlrAvqP/lT6Ujg
UZ2kUZf5NB/B6BL6RP9Py+lfYSyW1wTujN3/QQyNqaBUzpwniD4uiN78pGlOa3/m6B8f6GDNw/R9
RvjpLAaQuH6OuOjg9CV5iT8zIjyO9Zghqfh9V6iuwXaHNd6y7D3nhnAyCL0d4GTl+JEE0E+rk3f1
6mvJoE9dDzZMAd5MPNmSaCiVXEU+EUYnxnVjWHaN02V2DLI3fGUq8UP53Y1zk/IhgjI+ZyV/g4i3
lDU+/kODzGhuTTk0ZS+qg0Crx/Ynowj8PViRi+ZB0MuIc0NluowVy9yU3SM1ijPi0lKJQnfRgJwU
2yazYhhJCuS6VFIpAFZHs2LsSrjBoG57tNMmn0qDm2J39jN5+pRfnQGyTZywt8zd2H87kKHiehT9
69zyXReliKguQh0ednX6yZBqBnzlukquUSURYrfulCXieKjeKBIk4T/YHaFAer9X6yTwklTqSxV4
7gNGpO0Fw8n2BdOGR28Xa91acWfin+yVOT2Q6nv8wLEmqlbC6hu9QPMgGdK3zWEX54c6A4jOsWp1
TVcFzswPCZBTDUejlIExeszXUJCIIbEkgElOfO4Qi/pz4RWOo31iE5NGi4qyLPyEo2pb48g9GRif
jftLTxm5qmZSMr+3/RErZ1aklGGJ3L1mObrfH60maiHRvotNqfYRKduG1iucGITONtg/O30Y9vBy
fYBt7lOoeiiAUxnVPLvlIXL1Plyll9lDkDC9NJdeYdURCkcnLGUigw3KqJm13mLoO7dJ5dZ+cP47
7pLEYUO4irCVWS/vAyZ/bxuDsNQ5DvMgCq8RPAGAhpGiwBFqvkyRmNZe++Cf3sqHYioiS8UyQjxq
FnTcBl+bkOplwRFW8gR1y2Vl3wqZ/xCSqclvoA2RwIu9LKGI36feaywILVskf717JWUXgPd2ayMe
zyShD7xAP1MMl82OJdw08C8wsk68jTp4TCRbGGjtJK96nNQPgF5VvvI0elmN92I22gavVK/VKfES
b8tB4CFJJn6ITOiFuGKiZZYX2KnxQj22HJ/m8M8RzuQfwgcM19KT922qaJMBYgNYRtIqGZLZUR3U
9fDt07QNtCGHwHfks9B5KbKmx1VuxDBZxaKOxeQhk83kqJTzybrojSkUqrmfTErKWhhuIju6K+1T
sWYUhhDpMsVmTNLk1w70VSjzX6+ZJdqXheAxRoXVgWFQo431iiCiAe+fqa1UqOB9R5SPJiR4CT7x
UEknK4IjW5MwP6l3tYEaCGR1Mji8TVyjgeoWo1ybv2CGXmPUqfOte7nzxOlGbMar0zMJg/yEwawR
HM46c22oQPhOGSpXFK3tp7k/FgFOqoenJcQ1UKZA8DJM5Bt8XejRf9RsM5wEaPVqyQlWwaHUyxjX
t4zn4QEuxSZSoNR91TIklkv2XzFmlqw9K5gr7DoMNfEmpCTS5tPmMbrBVUsPlhW6Kmfk9CGFD0OW
weG1V2mALsOES/1Z6y47VOmr2c7OkMkeF0B3IFjtNWaakI1svAWbLM+vXWAwlP+MDD03M0aq94zD
JLavj8pi5pxc3jGZWmbfa2ZJXb7wx/5NIMdX1F0kl2eepTvAWXiClW9j1tlaHN0sxdemfXhYkNpT
hypIgAzgRhZv4rUjlRL+WagM8Qx2wV1fwjXgej2NoXghMxm2QRLBOJpjNoH4a9j9RVQtZTQgU7f+
DSi6zjKyVLp0twXnO14Me6QeVf4qZQ2pW7n4dKPsDoyP6fxRHAL0aE3o8jlzYRonvTyKOaoASFTd
W8WR73J34ua541rvfjdgsF0VnJS2kejn8s2TnMe/pU8lKxQXTfC1vVS3YnsrbmQoOjgPfYoWn2JL
VUKPcWlJgMUAXISkdScSlWLLFjjLlV+c2h9o1ujwNNTVaQ7FMSaScQcbFKpMjKc4MuJiM8pZtB3k
Y4//cpzVzGyFn35klCFd07GJpN8fKPaDJs+pcLm+ehuQcmDzt66GkXHkedgq8jfFO/MDC9mHVPMM
eYgj7hJvLEBYeICEcFuPQQJDpKWLSzEYMpHS9joSyonOH0NAWdlSUOayxVFQytCFbSHtUDHKWuqw
ix9igvOAr+ako3hC1e52mNLovrjhYe6y+cjnyQro0F6bWhitoG/8fLv6Xp6+F2EFOBmVLuSG37iZ
2Lp8XWwIyDGwiVgsJZm87/X2lM9KzdqMI6HMErt8B815uU3iaPre0shoOygqAYVLS51DwrY+ga8P
p0W9M1cflpRV0RZnAJWeuffqQytM+I3x8gRUgqXi0V6aTopF4to9SWFPPN6MGUm0JEGOswlRjL8m
kUwU0QX8BY+HLY+f0sZA9JsXXvGhiqoYEP17MC/lzNhrPx4+f8eMff8ZnM4JOlAXhDvCvFzcKoUj
6Qgi4HB2lYm0WQioo3f/eoFBPPpDsbo7ogNpbFqCrerGvTPZqeMxjQmXEe25nbRu+5n1HJolMBUx
cbCNUSDpEC0JXV0o9WO/OnLGQhbpsdj2ae56n5k3tA/qyluXFrl7BsabVOjmzPb1HJNMweC/irc8
9Fk6ZmWdOZbn2jB3AtEC4AJVOPqtGRDrMblCAy2q6AFiUuX61hjCMPXJ0RfKFknI5z+0lG5j/+9t
PCzeU2mRPbUa+yvLFTECeMYIqbJApKbmNzAp42h9b+4kEcgp9t4+E25GxHrB9PNIpZzaYGtuHarT
bbsoXOLC+Lmmxh/t67qsP25CpYwJ8pZBWbtgi8aVtHi5/LLr1zMKqIgoCAzFDtlyg7GwGMLMl9ig
d0Rf0dAx12jbrV48cOzmtMnaG3YD5sYRP8+QV58SsUOVp77dWKdj8/ChHsAD5tukcJqcvT7uXE4Y
iQIXPBlHb+o/DWW9BOEDAhhyEjSBnQkMipuF8GSaSNYPnGsdl4DloIQyKNiNSdACGj7QfXsMEPf2
EK9ycrCiwX/SSvH83AX+zxJEsqPCyXUm7dE6oWtrZClxvDylWUhYr+sYp6WbGlvEPcLQjwGz/e+a
vSW4b/zMX/+j4sr8C7w+Veltz4HW7cR7pLibxQvnBJ1sdXmOkFgVLO7bl57D69CDiRVrd5vXBYdY
K4MCPUq0TFcWTdZlkhswW+jEwGiSEFechaiFlZ3dZar5UDuxZhL0wzr2/xjV30bW66bHMQ54MuEH
cG7x52xogvTHLoWrDcYHry70ZD4hz1uL2HxmaG+Ktq//Ru2X529JvKQcMTqmTHvHZIoGzQIsmO8y
DW36ExJHBXO2hH0+n6uXLoSqiJKAxBnbRaMX+zPet/woNcaTFx2JrPnn1ELa+OdO4z6mRqiUL1mZ
a5J/b3U9bV8w3MzPRT2YvPu72wcYJplpG3ragB6wUwuatlzqO+GUDW7+HEPxIf1h/mjV4gsvZ9ep
QP0Xn/soiOhOrszcf5HOsDmJh+E20+IO0LMHeI4B+SroV2qAnqb5qBCga1yKEEVZnYiHPB9oJTc/
YP1r35p38ygib4IgLj+t+6Ou8I7rE7fv9OQ5yBVAyaH6HAPxX0COQjtv+XNjAXt3gsK7dLR+1Cxm
rbK7s6IyFzv3WgXe/Pvh+p7STgt+0aK3asNT+ImjcDIVl1FQjeXf70FVvXIRE268sXa/ewwcrdp0
NsHikOFtldqW8EDsZQjLfbB6QSF0lfNKjMHoyWXg2zDzVl3Ik3JXJEHuwSjYHC5my13vtPTfMNGB
uxbPvpqauO0BWPmnn3acrCikOGYo2YYYTQVjOpgCeikUtnJNe9z55dSXa09Kp9yPPdHnh5jPXYX2
1pULKYt3lWEAjRYtS+UFxcb7HWqp2dVQJQNLhWDh5YQxvfeeAaVjfADWE+BeEkrQlESKkG4r1jfE
8riawktR5vNif+if2uZCDFQiBhHS7pFcgu7mTjqCSg0PpvyadsIt966KcwugXQy6Lvj1g5u/Gp6q
DTjWYxeDWfw++IA07PauxwZneJzzht6s2AdmW6OAWWMBafKse1PoqF7TVeUK7QNGTSUOu3ciukEn
LOG6AugmmCAF0SjebqJlDwps+Y5jfdjGSU6NKaGZ5cZoBV432BphdLVXJXOb3aSLWQT+AsPHk+lV
6qPPQ8NZoMfQZcbnuespNFVAzngJbQx5/JrNdhROazJSdbEjwVB+/vnoRzFHVYjV7EGAu/d+NLxQ
iEIzHcWRbyXI01YDwi85EQFMZSltO8UOs7TXGIAJYadlltpOz1LrGI29lUWhSOmPwqqqsneDzkT5
vzA0s4BywTPknIJzfdw3S9wUrTnY60rDazvoZNz12XyUI4J4JSGYrU1+oXNr+hALOOby9XcuPexn
gxW4VbyiAKC2Rzi3BnDGSZ/A5RhcaqeRUEtoJNcRz+INNm/AGhLMLDRq/ylaIjZpLKxLVaYnG2Jw
WIGrhCgS7xWDSSsYecDZpHOfJeGG/lzu0woOYiCz2RqWZhVwtgasjYYdVs9qbTUShuszc5SEHLhK
lX4CGosSbnYW6Noc+uSdcjLoLIKvtrvoOSjxYEDrYa/7rJg9oBbv2l5eeJRBtT7slDI1NI4NpjOL
eu+D0ySTZLrRWIR/uvTXFnXKr/P6zEo4/PN72010p2safPN3G4V71ShbJHtnOO4ZjcV6PG2f+CkK
9HDu24aLk5YpbHGE+w2G3TCOeJBmEg5IFtpZxirfL36l/9ssuAthUEBxOlm5vXdEaBd1ybD5VPVi
OjjRmHdDt/1Dyh/ljUH7s2qaT526T7/iEznk9MLkQie0ji8EmUBFIsRbxB7uZ+ZQsApiWl+Wivix
8k1BHRfs3Q8CB/dywHuLsK5bi8SE8R4Xl1kU2n73MOaQdvyTzs7hejphSuWJXGFrTmz18LuCAvkt
HnQnTZYI1eH0iuVQcu3nP7H0UfFqyMXuYBNgIK2/b/K78+lyGQlwTLR2/EPJMqKSNKdaY4Awwbx+
kB+FUilZoNZJaiP5OGPX74Du6QcHImonQRYOUxMk2Ys7/zKabSHJAc263QW0Kr+vmGF57jCQDTMw
Ek6U9MLbp7WMHO/4jMuR7mWbdbynUYBVLOwzPtSQZwxr0EMUQ36XpKc2htw+VuC9VVa65sB8dP79
01GZ+vaRhE7Qyv4n5v0bElxnIDS0izTryGjKa/PEeef+MxuDtBAd+Ag0zlSIo/Ng+R0oIlVCwPCX
K70a0CaVfKK2zUT+iGCSpk06DRSc+JFf0MzLry9NxlMellmIRIWs97TWPhYbgBtwn/tIGNz/YPOw
ZZSw/h7HRpCFkBTX3L7ERwReo6XAeW8+R+T4UH36os8xGNPt5D2POM0+wMNQk5lSFfGbLmGTPwyD
o8D/eq00JLrQpzYHTb7ggmDuvwTi6hzbYODNASKjwD/jcGxuky/16ba0i6cRVfUGPKaRMCXNc+3h
8ft/8aQkA8S8DNJgDDDSOlI5DJq4iTiacEwwuEF9gHlux8YERjWymfLBTMXfk1Dtm6r39Vd2NbFK
wUUOxHFansF0FOHmx7SUC8MiTw7LhrY1VxSBINH9UYpVs41Y4HrB/7q1TE/iFZMDOkI/OzHS91gy
MJmz/QoWhtXajgJFyZ+aW6HFGvqKq4LvrmLDa2/5ZI8uI6rN6PFpaljHfqA4nhCAYzsfIsD1AFSn
Nqkoo1gaun7SZtpWY1l009Kq+b40Osbg6dbbQEU29IWIm2719d35sslnf2DzIFzqdKhYXsdeYVYh
+QoXogmcv3E/Al3sL8mi14LPmf3rCGPws9GJ7UFJyIuWxRJPQTNXG8j9qK8WVb3KdAhaR2yac2tK
qzQ2AHCLMEPaeHy49Pd90mCvRh3sbY+4pkKsL9i0roZMduIJng9xtHeSJL2/VgRavTPurIikAAKl
irx4bB2E+S2mP1K50W/yHfTI8y/9ev1WtyUVfE9gQ/aZ8Bmx6BDwI6ZfymvWWvxzPAszbzuiZXU3
9oZguaz5LIJC6zosZYxWyIuxiRAwGLHwwtSV4uAnzpiVH3NLQRHzesMaD+xBjNRgo7dgebqH8B3P
VvE6Tx5nVsYM9Gnqtm5ovaZyfYEusHcc/e17dzjdVFx9KiR46ZUTX7OprU61p0J9rKl59rRvUFaR
pdYsO8vBRFoEUBHeMZWvmFrk/bCb7P+X1furaVstxGPoLy65KXLsXQ6dtcdUfWPFSurR8vt+pfRa
UHupbJlUjJABKm0GWQ/0+21gLFF9l/Dn9398IvRVymjMIax/quLK/do+FWXGHeB/Bp674Z92y7js
X9bCwLDxmtWbQKhZ+MIzDdMGnfa6cU0oLyqZfROsCb4omavd004EufGENx7e1P/sCRYd7mT+Nduf
N1aLUoO63AFL2GhGatD+7TPKl9o6BIllO+a5fmSAI2muqZToMfzQ/ahiasnnwY9bDR35KOQM6IP0
DbhhtYdWR7vuH42jkjd/TrL455F7y/VcXyk2gswbrCGYF9pEbCfCzUpp6e+2GwejIR4MwI9BqDq8
/pYpdgdk6w59SoA+S5NmafGRPYg9Eo+mUcDAK0eSJqUuevUV4TcDowswGa7pDEVP/dY4PaBjTG1n
vr/sYs2Gv6ftYJxiG/U1mFZXj52SIGYSpmXuvEriJvjXzkRCujg1FWGSw9tBP5JcIQLtNJSwY2uz
5Ku2KGj3fJqW+DcnB4NFYtoL1u/bZo9E59HpLd95Ap40rcs6k+Mj8X72OqbC9S/OcnIWUfXEZ2s/
XCuC/fgrpCnDT09hQrl3+MWJm56x+EMJqCvMN6akm10mqeRa5okf91wWqQZh0DUWd6nCv7bwgOAk
vaSUTypdIBdLWDPb6cZ1eVU26AjLv3KkFojT34ol7T9r19lG0R5ZWp0YtbsZrk9n2LWqrRit4dPG
PyVd2NHBheyZWg7kcbZSDn9OLe1VXhIxE9TyGNycUoGq0X6kME2sXGebBU/78LMb4wkYMSOv1rDM
ZOCwWcTVozF7257EV511A01F3XcG36vKQ7glMrPq7w9FISi9G3kdFHYgK1c7vg7aXuTpkbnXbxAE
qXewJAfXhy6kDSef0N0l9rM3X8GNcDhQeJ1wR2Lm7qLX2mI1xxupu+PltlHtMy3MZYVqJbsFO1Ln
ZwNzbYBaOm2Tijl7/1gu1LtF/2ViJlrNvy90pxHvV+7ZJDQ+fvMTts5zEdfpS19QtjQHTzUGGHwE
RztrZn1V+UbpJSafJZYVJ4P/FaXZml2uJ8SWeKqh8mC5VdtYI72yIEB36yI9JYfYiXEWz8AoPe53
k0C1IViD0YKAIaGzWob+L6STkkTI6100Uty2dpmI3R36OAel6gsrAwBz8ds8byqmcjIHFO8bohML
6wldtEq8nSSJ3YhK03qaTFJi7VaIO4ih3jzHtWnvJWQFbjRLUgYthxJlzeBInxlW4qxNh7Wl2PCA
XfE2YNYLjwECnZ68i9XukpHlg/PVcVseYB3892dKAWwnfmR4bvtaXI3HiUoLlLT2667kTfigNbSi
lpvgskSr0T/d0P7WipbW9hf1MnudgZFpoo3XnAV0Wllul9Erjp+GsL+qq3HtE0v5oJGyjuEWwDab
ZnpFOD1YWneQQNIKZEezg/jHBc2wPw/6vzU69k3j/sLc/UFge0apRetCSFVcMkPEgKzh5eEpE6M+
R6oJ/hDzW5R7sV2+6w+hac5p5DzL0LofVUy7DaW6qBnd0cHIcsxO0l9WRvl6z+V7c7uAnD5BNFCc
JWtza0IM70hbp5I5WEPoUcA+tyUUbrfztdiwwyh8yF1gW2+5tEI31lA4mvcZUqNs07ju0f2FXxqY
IbXHpQ96AU9uBFJ10ZhZj4PB9fSZHqpbj1RHSKHmPQNt+fCblhhWoVeT+LnZlOZDDcNN3sd+wAed
eVzyqNsXyTgioqcmTWaJ619th3PFcLNicbT2rY4mPFa0UzmJnFhGnzj5G6xnj9lxz+jpYufzNAvj
Hlf5KbmXA/MP/9z7HTk3El25x26KNAEuWLPSnyXi8Qc763At5osacu2MGvlxR5uN3XcV4TfcsHaI
DwMLdm9vpy5qnmXXeCQ0bXlPwnstqxgtv2UQ8i+q1z3W3pScx70OPI/ovPFIkn+xdc0ZE4tfGWmD
8l3huL8tf0s3PWzw8v99d64BvQgsyUghC6UarJ9IiGmhsUJGVCCzYu1X13TSTdOs2NyQYWKnaoju
G+qMPDLcy2FCG9dOomrDtRX0RdgRvkRnrnOibo+LvXJrvr+AfgQ3kk9+YXUeHIIkCMq0tfYoc5TI
MClz3NEB6EMyJCtvC2/Slt536EKEz5dR9gnecH+q95G9Ryvq4mewaeeXsIpk+EhOvybxKFsYjtc6
EAU+sgG6gQS6tKPvpgYCwWorFZD3vnOb7f4Jjlr54kvIMEBOdinXejhV7XrbuhcLW1MV7XqBgHvd
Vd6FDKA7WnQ9CNSyHF4yZC/u7cw/HYDF7He9bmbNXpABzNdkvFmHvwdW0aJomIqExsgdCxkCuSqW
gRESqCjI9ay/GPZfxE7KLlVGMY9s28jFdz2B5GAgUtnOum/24gck2re0L8CsmGYRjf2X+sxL0G8U
IwZhfhmSo0cTiOYLA2L4l7k/5yGsDtGITvR0W/ZxfFkJZwZSOoUJbO+1yAO2njkcFZUPkU667FSr
5Jrj6CQ5PKkMBgmivChki0ZQcS4m03CRgE9YXDRBR7BjZsp/vtqS7TLhsG6y35Gha4YCDguvUNw5
dqpxmJbVV6EndhumKSPvhOA0D7rhEyTOqSiwDuMYux0+Ba4X6ooF2d75ULcJQ0qL0bzwHCfO/IZI
z8QkSvBG8CEQs95HVWR/OWrdhM/3RQj/Sb/hfHtlVarCwo75Xf/DlU8NLqpjco+YxmNxN4/oMks+
ZT5LmmxHC3/cwcLwJ2YLOO3RDmAMw/D7S7sP+YroG828RsS34k+5DkcctgxupK5DZwWnUc5MKsLL
VGP+zDdxBn8LJ9S1d4HnZyJHwqrvpceId/BZVjELDQ6GMgpT6p+/pQ3pnpTKoL8V6yCewlorZFxp
hXMuhfuDjmmKgKqJvqFtpdMj9/SeMr9HFI85mq77rbGVq1MQqPXmS3WUIyYSwB7M0e5jreD5H6df
ff7M0cdz8cm/JmVmKUgbpzTTm9a7qPh6J8xilqhTTwAwh9nUoghE8DwTkxRibQhVtQtrCJgOaTqG
NzykKTw0ikF/UfyNAc8QGAf7GJm2a+inhljCp2i5Sm+JA82SBK3rhxGOpcSFZS5BPyki0GNMZDCy
tdfUOojwwawHSJNPU7Hm7/FFLyMtLANkdRPyGcJYSfmpYFgrbN7e9eVmAIYPGKDSIjq8nDzcqUm/
f3tJxIq8CynMKn58XAJSReVQPHA1IdshzMKta9e/EllXAiHy8a2XQWdLC+Zj8vP/d6dT6CQMwId1
7oelCbQ9hjOMv/6ESkhppa4bvSeMN/pedJGdcR3yF/QBD6HzuF2TXCY8kXM7MdF8xIwbKt/2nOWR
Q5vH9eiZCGt5hqJEOKGkq+ipUMsKbhufAqDiZoSE5A7JT53ZD0A16hCZZH+XujFOJxjnmHnM31S3
ObOlV5/4Dt+oSWMAV+gMnE0jbhqXhbp8S+R48fe6pPN8T59xt+ntq3pmig848UwQb0vByzhB9r3v
+AfLp6mr1mrgSRVFKY1ITBhzbVlh4BDjCgO272lHNLrW9RuuXVVp/zCr9p3QDiy+d2JpR/FHl3vC
CCGgUWzakLqjuPapRezO2QoidvSn/HyRZbgkMCzPWRivLrxV6O0pNYgA5GwT3ILJFlegpMuITihq
24FqDDfN2KBZLVLfAlert1iz9z1NK8oj7VQXEPxToSKCQ9wU3b8DD+p8tyectRtRES+ZXbEFeieD
YfjlrunuPlcQt/GoiKdn0yJCDHBirZwlINVAReKd/zlutHuGFpgWlz6qMta6HnoTbt2/CVpZaOVt
uCVMZWIThwFOwSuIwJPSQ6SohNNek2ymO5NF2sVGinTl1bvDlas6aAIKH46JMDSCOqi8aHpSfszy
TnT/ab2PJq3QhueivOEXfBQ9aFwZwz9tt2hHNdwamo478poH7kg4vXs/u9zq2xfrmc+G/Xq3o9bR
qnpmUuQdANNb/aSk3iNfMsnUBo5G2RWwah2MM72yaYdpz1VaKem4JttKq+pUddNNS7Ie1Dp9/U+L
8v8YeO5nxKLB1rVYqLWIKYQ/G2+3fRCllXk5x9aGKZwXYLWbF9KkESmTSUKJE+h3JhtYxbYII4iQ
vnbnOY8q7XEjvce4nFsW+slRjDRzghz85IaAa93KQf4MDpiSDgxLqWyVqLfrQn17rDCyo5rEfPqo
OYJcNQIgiXdcGpAml5Rkzg5UACtMX88E9BYoXTHxSmyKkPfbFV+2ka8AYahK73n6lTkDL2WEphzM
WHfnirZi6EfwH1XCDjh4xYFgP05/bRr+fbbC+tB9i5ml0iXjwnnG3zyb+ssvzZfJZI7A6BAbU3xS
iTJ23UvJE0GrbXAbfJ4tuH0Otd4EENxj7vrQexjmSbI7c4xSqnut5C4vxdyydSIwkiw3Uje/y7Ed
QFow9jb4v25GZ7k8OJlKTUDwcKORnk8qh4TKLKcM4aNO6R0rnDy/Hw11OWSbLBZqFa+4nViru0fb
4DgFJCvrkyoy5wBs5bEIgtQXGXoiLuy/PO16iEH3seZJN6zGuhlqtrM06TlaI/I39388tJpQFVXF
a0/rzTOlWMuevcHY2U349RqZObRcrgDjsIB0rBd4JI7XL6PImNkyRLZSYBT5ohPJ2/QDXiMAGHf8
NldJ+1mB858pM0Q2Ydh402OS+4jr0b7HOFdQW3N3PGEftbQTTF6uOBo4QVqGYd+dboC6r5MgNej8
YeB3UM9JGE//n6esoCujwH1PM0I8rijkOLvZfeO2K+nUr9qwWPkd08BQggivBDiumgkSuXMNNFop
sbJOl4/8lE8qg+gd8UdQOjoMb9MOhRBuEfmg6ik+Um+HsBaiTIPCSByPt+RvxiGk9LpNnwTXezXG
0u8p1Omnj+Y7ZvktEU5sSda+0sgEdF7+Hm7ZptR42eQ8lUAqfPiB1uPSUSLdXaWFOwokjDGgyqQ3
qUUKT3RdHbCU/MicOHWv7Ayk86CPAnoD71PVBnNed4IEN5gBJkiy1COPjoyt780FnfwIkz8YY7Ts
r/OZCoCI9CuUuTNa426IPowNpOT7LAb5tr0Xe0WcvzQJBMeLTq6R3pIpgA+QsbXJrLJYef/mT+jJ
WjcjTDwkoAWEQGtnz2WkN1iDDDy5NiFn09nmr7M6+9QaioNupOdtkkGTw2uWmFaWv61z53uk1iBR
LB/sSiG1xCbgkLR+mtdT8c4P3UFNlGyfEcYhshO6uXhVZbDH05gcxfoPBz/df6QEk2lp08dODs4I
7jcsNzDOD/PjRjAdUCrngCJgjcvURvtizYsw3p1JlG5dZPdyIDBrpbc6XmKQJP7GEJt7SuWQObwO
Vvc2pyBNFgEifb3ehWoeypPl8tlB0Y47pFVbnZzmDJQaCiEDCeD4lnZGaP8zeX+unUGEilJmxuiU
Lhl+ZRxfjXZbgbj7GhfDgHS4vmzelz3OeqGg5LVkDhMIo3nlwW/GAvvaLkWJngL3CSH7v4ko9eOI
Zx+bMtVQ/bl/Qxx/QJtIVS8SJUU/81vPC5iicb6VQvOgDXSagFFqxKTAnBj2d5ebFHnS4NuNuHi1
q8ei3BPnF7eOyRY9yWXWhtM77bHhVLrLh5KwzXGwfSzYnfOC4K+OMkoM688SrjkB/sIb5bwVrL0g
zWh0rlKZmWV8zu14V7etM269s08lYk7f2jYCjPcJAnY+8Wj9dOY938xnpALMtP+eiZ2ND6AvSoPX
Kb5A0O7/XiiOyakyKknE+d2ug6tm0+61UK9fEG+V8HlGDAZH/hicBL4ApZLPN7E6ny55rrHUTYkn
rdcLe2a7oTGdkvJtUH1qiTVeOA3h2V1/aaGWCrULysf8HPkF61Q9hJzRAafQeWrXtQcNDUxr8nwq
w6V2n9FlRV0qH3JrGDwX3cPKC2d9xVO5di9v7lWMoWZj2iOyLCh0KnvVoUgZBleQ9v7BXNYlLgto
xS82imx5aDbTkgoV8w5KiytLbyLIHwGZI2aguWZZkDh/C7uNTaAHrofof02smdJ5wj3pZlEOJk82
SbnMgHnNo0gbgfa2D8CXp+mVJWx380eCvP8XjEXXn8xJBS8eDrKOzgmjsUq3LBjURKUNvE/7DSpd
wOc7tZHnRw/KgNxoZ7s5ZeuF2cKA5Ga0HhTervtHwRFsq9rrkyeBU8hpoWrliLwJ1OyWPLCoveKz
koBNpmaA/BIQsPOkImH5b8QN6CdY4VwijrsqMBXgCq3jANkOP3nENi8cQM8MfmExT159kTRtn1jP
0bm3JEyBBO4L3BRAn1DW81A19c3YHgyeZVT4EyuefdToRUIqM4p0hXr3qRrVL2cZ7qEma7DrooS8
cfXKQURx+lXqWUuwKljbL7lurOUWrN28gwhwdsd0WfETzKQraRM75rPc2IsH1/1Jtu0NJmTeZvyW
1XPXwk9v4BBZvVjlOzej8y3io6V70SUEHeJUcQ42Hrr9zmmgyKRVyzvU4EI7jPASrhV//jVyetyJ
FYgsuJoP8E4VlqSEibBcB4vmn9P2HJfiCenfkTLC+kxkCTbA55EPX36k2DvolVkWCuhzTM3rfA0B
4yFozNAuRxwec/FvdX/teJkwL+mdKyTdMFkNeHmY+cB1wfG5qQ+sd2tRSRojaqkY65te+QLE1egg
jxsLgPy03fXIau6wicmgzvHndf0X2QhAgdIv7XdrXlm1MOahDGLZI4VZL6CME1uk4rR3pUMZA6z2
nknHxf/2jf8pUq+llY+zDEDlUxufJ9EeCmy3EDNaW9S5OazBucQ9pIb6y7qEvDBhQ+lV6/iJpOPt
5sz5zoNuf3LcgwLWJh+/PN6fTSRr9piRsqap97FWtg1orocrOjREwSHND4/l3yfkZFa7cFYg2jZq
7BiYnfCNQuhtvknrGNjI9Td/nu3r+hsrcWD19I76m1FMZ5mbu4dftG23p0GDLRCApMxUEioFXznR
Snhh7ySd/Dry/C4tx1bYVjNQPXqvOVPEsPXY8SeQiDmJfkNnSHLEYkoJN+uNQUFfQ/Y/K4JusmjE
RuDkRwGmqUCTd2ZNrmbLqviLPH2oIWCsDkXBQCMzSuKfmfIKBdjAQTeyBrOLo2GtPRyt1cLEh1YL
rI0N9DHUEUx1Xb4zUFGtMfKKUYrnxIeIAEVk6FyWa2YjTSMrK0V2fNF2K5lQ/MpaNt9sTYO7avSk
htA8feza/qPYa+jK2IwV8A+HrGgTa7rEEyACATVQYSg/vLeGjbEEq2JUAJr3JnyLF40i0gZY0Jij
YOBUeBYvpd6F0zGBXfp4Tz6nxmKo25no24i2k1B3WpuJSpRYAWCouMOv/sz3I35ERS44aBpxMoBn
hO5RSVt1NwwzZ5hdEVnPs3VhXFJi9VuovGqNWOJxe0Qp78qywnV7K/ICliNn+ZVE9eOsh0lle/NJ
kMOabxCFo1n3RZVH+z+xO4O0mOBlz2zR9TOzf0OZEYsQOhG17kEoMifHpb+OY9rzaT6er+CiqlBR
qMnrUZ24zN21fzAdAdKPto2YTeniahzcRGTtpNJcvks9p96oLK0l7UmbQYhXZ6tJqvceKO7Yu/xy
z29iFTBzu6Fj9N67auyy+Tyg+zr6WvGHMka707aXQMWWI4wLYsKKP/i5OnQYf++UzizYu9SZaNHT
ptlkoUA9uAExB7k7LpCKjfYLRoSt2Q5tlNecHdWJJx+jRKsJGYK31r7e6p02zIWJg/orEGNlO1Xu
lTUT1ETtN1q/wxeNaqNHS7aNfEDJvefdFrIi/hV4MgKGxP7K26XjSagoE0D+yQulcYTssR+tFSe2
mkUTPu+zldhBoleu8sxSanX9bQOQZeL+WRHAM7iBam4MEUtzIjNGrV4bwS6MMF3pVM1UIiU5Zq8T
/qcjhl/AZfHPzVKFELC+dY8xI+pkRtnwKOvWr4g5UJi4CyRIloBnfNiRUFnCYtCLbOkLT0Y6EXm8
wpsuXhLnjHkHMfer/gfniOj8aAm2Cbo90FETvn7XUhFSssbeFGbhYJnEUbFfhKxvLNmYCwyKpd+n
N8r1hjhcHQ79UGll55dd7hbq6Ke1D5U125sgHoJ/AgEkTW7OGDUMD7N7EPtm8zf+nfQDgcoXcUZS
WEQXtxIiGu6N8lunQ5KU6JiWVgjvxwUHH9tXrOxZ0j1o6Qdzeb7iI9H6QMKlk+fon0c5bA/MZ2eh
hNW1axuc0OLnAOdZgeuHPD4NF6O2igszTUGNMmMs2k9f53DHmWR0JzbY9Dyv8hOAoE52cK/W23tV
R/n+9WIMoyD05mLOfjDF0sKFbkRlvz9dDn80dOvslMFNaPIczOXCIGgAbA2LIh7rqkihG934e/aX
fTkFOeZLOV1BpbN17KeI5O9spnUsCd2gO29g+VV2o2VBUJbkv1T9sH2FSby+jSNSutyCXeJQPH7k
8n5sbXH1oxTEQpQBaZdkwaBqp8FwGu/EXa8hMmrG2d45DjGB+4ZOy1uZtcD013E3aoLIUVF5jj5G
dDUI+nJYQwX904Y9MhWZPF0Tlx65J+HplotWNguphpBATqfLVpMzaBL+qMzbXwprEIhalsTx1/OP
RaRMogJagE88ZBRGLBivBQWZTirW4IswkkWzxR0blt+SujDxgbYQJVZrJHc7VBE7rLY6MH+i0+a3
2Km6FdJe0yJtvsph9yZOIFBKVqwaBpI2cZ9Xn+YP1lHNK5wzSGJ2p8vIRqbmA6AMoVgkeh6BwY9i
AeGjpPPLpbc23OyuEqhyKiedL4mIyl2mmpCaEJ4eLYu68btm1vwfL5mrW6ToP+kMjkMnNBt/fsef
cZx8O3prPluHvcwPaH3fCtpymJgyi3z8EE0s+HnXyH5pXKkTIA2qnjr2BmvASgBDSDoZ7MlWZaVb
MNkCwVcqW0flcHZyHrdoz4WcWFqHyN0gR1JAPQ6IhPvC0uf4os1/74AhY8/m6hKVnqo9TQSuKUI0
rCFdfUZnyeVx27LiFTHwarQVxVFeCyZ3kS8FsQspFJAlHgfLEh6Y4QZEidIQ5txXmfobjBc4Wn+p
+Wa2kbP8TKq5NC9W6LQDUqzjjiSzeY93WJekcW74sAKuE4p68rzps4axb16ma+ybu9JodCbq8hyc
OmoR7R/wR1eNgAufCq/mQdXRMS7LmNe1tnoD/X1nQ1MJJH6JEV8mbJpdnbGpcvEYiSknoilwSVuK
wtcsF2pycHamK2zwTQHgztsjnS5KnZ4oTx64jEaRZ9W7cs09OKEnaVCV1JR5ALvOhUJgdw7vOJZ9
ukZxFVmSwGx0C2c3q603QVK2ep3xQSzD4qfKjPVGMGUQ43b+4mSZfHhRgmYSOQZI0703t4typL+N
FxsVuLBk5AgerGu5zxoEnVCmLVZGcOHbx5boz/HW6gXXMXGhX/9ueC0pjIv8lsoHJ07raBtOoCxS
DmEULv4Rx3qowGLFb1vQeumiXxouKxtUQ03zMPwQNBBjITzD1VSPKuT1ZBYxdwvR5nLasiS9qH/l
foIP4fPrScX3TdBf9lerkGYYMkEXBNwNuBMNLNB+27yehOClSG4CpWcdXvacdJvWUw+zPnRTu03R
ciD6fWeWa6Jm7Hi0cMv364lXm1UnncLvM5/LX+URWwZ2uhY1FuoS1MZHITSpiuukyMLf/biT8L8x
77NxRcncJdRI4JZVXjl0b1sAl2NptYqcxZcsjctT6lVlkmbyKsWLW1nMuDXvhUdkTakU7BnezOsG
aBjPwkLdBRN7R7HbIowfJMxtpktStEbv6JNIZam3CwlpsJTTuHdRVEj+Rz+QT66odAEJhvMQ+3fJ
n+Q05/wMQOVPy6ux1lrOfzB37yzud0k4yJGjmYzQ0p2oWAHVJ/6Mty26hlfS+/mVMlu1UBi+9k66
UbgDkrcjr3pcVIsaY/iCaYBLSviD4wlp34ZzGTTGiRj3LLEm51dN5fr4L7fdGvGB+BOKaOz/Pv4C
LfJKKlIVF0JqQ6nej8oQHcwmqOt6UolYescYimUgYbjasnMkyezrfzoa+EIzQLm2Zx/jEnBzjfCY
UCU7QFmRD8MOlvMNhkziT4TyxUb9D5j3MQCe64yyY0GlD5Zdn5MzVYrXddGdzq75mwnoT5cy1TVp
dQm368jZaVnyjwqJLbCZhpp1G/ogR6uuekEpijvJcEsOke5EO0scbkEVCSed9b8Wfw6d4bUbtTkg
Cfw0JaVFH7yC57PoD+aH3Tt8PnQvUb+klHaBEW0fJMhBDptulrgToaKpUxnBtSUnjF+Yp5HHmFYT
kndVvk+utiCH8d4msdYRuvwZvxSY9v6n84kmjD7LMg4p2NWoJcXGBCce20YsIhpDXHZyKAOS1Ho4
S+seP68kRxXB6meyu19bY3e2wqJe0NrUvbt9UP29E8Eyr7mmzD4vnhgxqfgYRj+QBWgiVbscnaYc
gTAQyFRFjDBU5laqvS+gH0XvE14rQw9hu4CIZIjrIqOJ096nLvWl8OXvZjGgiVf8ueCI+hBAiRuj
OUEmmu2O7KLWwewGDXqLmR8xI5lf7/kmftSxrlS8n2t8hrWqaCDK894voEFRzFWerfR4dAZ9YpfX
75sCyPn/SnRN98ZaKsRQdLBS4fJ9kDvk/OXDKA7/sf2+pAczXihRkY/BRnNnjbbvvcWA385EGP0G
FSpOGliVrGF3EP0uiU1NgBJbm0NWaX3kUfmNi1uSCNzOFrlRhx4Jl4tV6KLZgw62LpsLqxNauxno
hUeMatcq4sDDn8rA0ubb9zyoPzbmeAgJ7cXHS2pHAnK4KHWKl05ZPjAIPBKkjLTjKqJvbs434BVZ
PFoo5WkCR4PmxzOgG8GhE997uLjRhOUqqsTpnNwoAi3+wa3TQs5tXbKQWkP4P3Rzoj3Qw2lONkvo
8R5IW5nre118dCXifq+YDU0lnWL/nBxU9M4QZqdv2zSsjNfO0NIovkLTPQ6vbOx/OuMfKtxQDgca
aGfyIKVfSUshUHaDybQUyObtXdx4japdIBdprQqEvMC7aIYP+o23F5UvXWAXwGa9qR5yQnpa9XMX
eGliOnsNlF91Cw3PO7TuM+T9NfY5btVxC5q5KFArVriHIfSvvEacclsCIluQv8nWVmP4dzNsi9pa
1sH+Wvbtw0eedytKQDye6do4KiI3xwwWkYBD7EG/ZiLrgCF8WvjGhRCmFz7YXGgnOSqYAYw0Mj6z
RqGip5DVTXoOwfrce7i043F1TZ44KM1TNo6w78oG0Jl8lMGq3YKWqgBPruxT/uDhW9xhXYWX94on
xMpbFo0Hr/mjgwZ5+Hvt+eaPSs3v/5dmH+npAW/df53NJ9Qg+k/OW0+ucSFpi9rNqWAk3NJTEt3D
orQzZ2odKQUyWO8J1NPiKta2KkxdgCItZo1LZ/QNt06lpYEcZsCzj6VvHXdJ0gap12U2fXqKLkhx
qMqD9nYhLzBilRsZXK38CRhuaYifLO2KD6vEf+cx+GSKZX9Rzv9FVhyOfau7T9rcwVBqQMjQIAyI
ZDeeCCas512/sJZSDbqz2uQlQkQB0LQHEOeNRbG0uDyYes4k8Po2bEYrJLdFOZO1I2fSzgHqqm2S
T0OrT9QRl13k5Dh7gQUIZRaHDhGNuzHuRJi7UhLSXCjjG6c0OWZ3HhhjFczicX1ezbjJwhkd9nBZ
l5qp8hQETYqg75VlgaXqgMKXseB9c78cwOB2txBW0MXhXL0/AVuG8QzXAA08evba6nLRhVCW5Vx/
J8b9bJSxl28gltS/X2ASYfxypWgp0XjU8o8Bhqg22RB5Hc90JYYyXvoF4gR9Lz/nnovPkW0Q5Vvz
+6LzTahOuS9c8PuCwRmXYGzLlzVDpooh0aAtp2R8Be97xVYT4oiG8fO5KqvEpcBTEwfkyCmZ2i+F
gYHnbfdBnD9Zi9n54CiWqOb9kwgc0PH5uUPiMoxRfwifj0Sw9XrQiW3AkjYP/b3YxUN9mZX/26/2
3NDu9g+CQnWetjiMtRO5z5zaXuFuH4ae/TtrRQhoPlDBz49O8gp3zOPnpiDTOt+fLqxUsI5ijaWy
VJQ9nlEbD1v3XF/jQmT5bo4k3ER5Cddl0g3yKFQ6uPEkgnomXi9kmVKMmclAOTn9QFGZmY37f/Oo
vcTNeAEaSkfh4tzi2IZpO5fzeHQm4Re5WBjCOhMKSSNYVEDzJ1SFd+oacMhjA49udVqbdbe/9+js
m4VYCOMmF+BUE3OOGsiuxk05nCkPlysq5ohHaqYhSdq+tTb6NaAOsE9KWf+byvAxtpnGFMYiuvxM
yHZNsscKWl0cy2ioD2ytnOa9Diag66I6Xri1vVXtZpMRcdr9ZDWy0b1h2ebNtlgf4NgLUuqOjFwo
EGyzr4AdcWItGV1W1Cdx0pcVSvq0Fv+g+jYuCnDXawKNjudA148Mkit0g8K7HwKEZTCwTRcmbsat
kzk1/O47GjUtzuF3668TMcEEE0RYn4V6a1q69c68v90NRsr1Af+NOmGMTufVYnd9EGFkcN4LxoGi
Er1/iNTEzrGEYSMoY0kFyX9Ok0FuSqpTZxuT/IRw7J7TqQ6BBkxJaJqp5DokWzIm97ZRKsnLwGgs
UzyvQT5zKCN1dqbMtJQ+npsykHdtCOz0vG4rpZRu0DK5vel+5SGXudS7KGXFZPe2McSo+cqo0Hud
M7tS5uPOlQXJAuR6eDYwl1UlS9EuGvAJ/pkezeWQKoZAXQip3+GO7i7y/jEbHUhkl+IpkT+AGfM7
CpSGMYg7XaQ0tL+9kNt4yUoXMz2Ofa5D3HXSaiSKMvvXOZKGZA/0TZrJM2tqameWplNLV81K8ULD
dfPcZQOZY90D4krrap0WE3A4ds+m1v0mbIK456i9UMQtLuq4yM6JzG7piLAwXdLz+E3Rv8Ao9l1J
myk+zYLMz+tN43v3DOlEV1AMxfO3NhxoXhW8NQzDF8SbVqEPt+Da835GW2MmD3iHcx4K7pa+atrA
Yw8WTq/m9Ze6pUVnONtTJmts0F0wRU9E2PoJ2hm/X1pBJN3E/QuhJfSrY1hJ1NmvQqztBr5OGlTl
UbtveKKkAETlD3E76bTgzMXMyZYoaZO6FEzp04VETSmZ70Ch0PSMvbNz0/YTVD53g/2H1ERyJGkk
tUCUNeG+lxjH/5LrvyZnLS3A/q0ib5WdXQpDPVA26tBfllRTaaxfOVWjkUz/Hwjf6Z/TGS7jP66n
p3G7XrVDZzLsLTMcDHqYV82DgJyJKL0hK0DW56tyzM9UVR544BX9hEt4jyFXbRelpxFj7CmJvSnx
NY+5ucCuSynDlAOUI6k1KgS3Gim9fRZN5Wy63JREMhO3YUTufyWBArxn67OHkNW608R1F0nLOIKe
UWiXYbgmSNG/G2lfhLCYpkYrdoN9VKCrUOcJp6Tom5OM7o4/ftP19BGJfnnDVF6oO+xnlpXOZW5+
G3UU2qQ2go16y2cy9U6GhBMXzi8cUL6Z0EPag/Jv9tOz+nrDfGVjpc/xJjEtHZCh/O9EgvnBp01i
NGXaW0BaLOYwm7M1DkRb3KqONnyss1RaGj9I/Y8Kzpa7FCWef2/Fw7JSydKBrGjAzSkV5iLVXvme
9WzLMZtLB+t967HSRxG5C8L8vweOh21fwUFkYOkt4mnqlvdyUl1WcB+yY9tYrghsJFpbU1BUexe7
SvWuSGkZSGKVIlpfClAo2q+8WftmBdEplQvVObsxb3jlaFkkP34gRLYGkX+V8WvZnY8bDyPLQUtt
3+xbftbZ++UqM9EVwbetk7BJKZ7KGalxhQwD2jZs6LLXwW6zuSG2B0aNpm6LeOQBFuWBLJ/u9c7s
pb7hze1Ht0EBqIayBZXihYneP7GiDgWggVvxgJBZPXnVip95UV2mNGcENxMFCHGWcwzYISPyr/F6
Bf6F2/7VRT20UQysdvf5mUitzFGyptLODT7yyiNNT6p8f4R1NSaiLWrP9SOWYSOOylEa+tUhAOxT
9TmKX5k/0knbCxYe8owE1SccSdCHzk0P/1jbEI/8BOW3fQadehLfMmtzT27WaUR6Vd7+ieBlXNMC
ANVMIGeQEh+OIKHwCe+AWF/1mh8CZE3I1GY94RJRtgoPhJjx9WhaB3EOGWjIYuYuIE0myQGkIq2Q
YGxIadkMvlaiuKs3GElKVqLrgVYeGknT0AK+vq/GKQGQEtOusbYmMq5WhFX5irk4AMOsqrwwzCJj
EOqRwLI5uIARDq9dZ+1RrkC1LfuisXKZLE+YF8lpzAqlcxQUtV229qKf41pV6pO1ebqkGLfwneV5
mjqWjlARtqjPL5s/jcRQXSX+EkDwi6WwWAsXb/lDu2GRaEejnkItPHwPXyiFMhSK9DmshT/0G3sK
qH4kriQ70zNcC9IN80eZC9ycSbWskMZIox5fvI6CNiCgAPNfX3q8u4G62RikPHi/hQ1NGe+iaMNC
MKn6eT1Vi82X+jCOW1osqD8zkIkIZGdToCU5lHxgtW52ftKmsayOxg/ufGfCdfgkq66B49Tt4NiG
9JWAwfeJ8coDBZQ77UTRM43idkUJ3Iq2SaIiRtF4MT8q0uXStwJwmJihQzCK2BykQc5UomVVf+WS
4XQvBjWE7WUYjmEIK55s+aIFYrzE2FHM47eyCB2r2lWYBhlrYUXdHZ7jyXJJvd6GCx+7Bsj0/bp1
PAroUSuPNRBNY6PPYTJiq8kbJFK332piZ5OcImX0T+NbB5wlyr8GLeLeMMNJb8tG7F1BGpNENtPJ
8huAm60U8ah3ko2UnLam15pb6e9STjjVbikkLS0WWu3KWVovUX5yx82rKdZfjh+W3ThkCwIGSeGw
NgjnRfcpn0610Z3P02w+TQANgmDZ7djSyW+6TV5X2vfDR/88xqIMtqNthjRS4taPRLCYnNJ9UHRi
vqVNRS9mwd02VebgqlrwsegpQxhfoEUximX4zX0uRg3ze6qDm5tOxkp/phaaWf16+LeGUOgxMMb2
poC+etV474VhYNDU+2nsB21IumT4n61mvMjbDOiSg4uNkjUvgWt8Hoo/jkou3cUBwGcRmnT73khd
DLOYAGy7v2XIm/gexaLU+m0jPwfJThW5aTvnbH8t34efQ8+xB2OxDL70P1sq4KR4ppJbUCpleOYR
MJmAiz9maCB9Uk778v9pYn6LnyZ3CRF/2SUx/+57yav2InG+srvcMrYaPLnRIXq/0clvmXL/CdTv
H6CvUEhzOsgGNbXVVP9EX5GHHKE8gBxYA3wmwF3Z+JYKGTMSLegLYRz3CoR4hCR4mgNfdJr6f6kk
kBb/i8CtD82XhIB5UEviLzFEzVN5qq2fWcQFkspqGOEbDCHdXjZqtOA/JL4fL0SH+SPqVL3a9kEO
fITAQrsD03TRistmhXzoqR/V5yRqqN/tK/TLAf1nYuo4wi0p678a0mqu0QQk3RkgSibkx5ZEHI9Y
9lilvHmfqRQDfd4gLwLffWuljiDzGBiImkdjogrv4Teyh0gKRCl4ru5RYg3GN90UBXME2M9CD7E1
pVPPT9Luju6WhKbBu6LSm5Gn/g0eJ0AjklT4hpcjJuft9/I+byawyPWvBfRiQ66eLaNvCS5273V9
/UI1/29yV3AUxOx8rwnkT9hQhR1HfDgDGAlIAyyJeJRBbRLSyr7Xs26JfYoqIan2leDBj/p1kqAt
4QMyw/qndkWUn2hCzLBGkyUwPK6f00EFJw2LQXx2P29GV7i7TcTkN7zNxwIww3j3C5kJ6YBq6/GL
MxD9Nz7Iq7c91G/2BAZ+EofVAIlO2n35iGfNJ0T846fBymoLVe8sBsiVWKJ4ccutcRBhsQwRIuPx
awyAYaw81vJY6xHyOCileaSg4KA6rU87JBat3zGJC9oUdhx8hOVNqwG7z445dC6KxTyNDyV1N009
kuDyWpi6Z7o90cUMqD4nQvrRizkGoj5N7y+Z5sLuzHoS5qGFrG/OPjNRINHbcqyqYoIjgg0vgxFG
qBnMVpnTVIBW6vs1o9T5D10Hf0pfxy1axFCBAvdJNSXRMAgZFYdSb3pwyoMNpdhCTVdiVBtvXb9Q
+loUvo2nz8TNzDUJ9cb1ER9eyZD4Qo2or3I3Mdx4D16BUWYzhoKfUpNu2Xv5XqVeT23YheATJbQc
byURaReTxuMT1FvNBXUlJGnK75OoLmu0M9YsLLy7III6LqOP4pv0RHjQWgLa3V2zNgSbW3EcXIu1
aKwwZ1KRMS2K5nxVFfa2WMNtduLocLsnQBRPKq4doktjFcUWt3RhhlS0VQzDyjXIGoeYJi9Ixa8i
143+O0JMuYjdoyAlYS8PEh5Q1/4Mtb8BgsSedwgkdOiojHx2OTMVPAgbLjqXfvrsuQPEV6+n0meM
jCjFLhmd7RrnsiPMJuxvTNLDdNukNGkvt2lJTLmfrqSRBGybrPreOJFpI6VzJnUbr8yeLdza3t9a
1isPakOTJMg0e/viYvxo/5k5EjHoIVWBtMtGnjsycPxeuFDaQ5o/OlT3F/XghpDFX4boadO61/TF
j3/zsQ7q/tnW+OPkkRh3WXN8slGh7K2nC4w/BQnVQ7OURTrt8MFZxk3iQxX2hkdsTCOMFL/cQwF2
oQpQSsJjJTFqj5E9pi/fNWgw+cyQN3HYbanER2khaacJ0dlEdZluOnyILZ1zah0Lq8iinKkyKINb
37PVoV8hBzyAy4W7/e0aOgfhF6KPhhgmxe2OrHILdHpTRjxZlpRzIbaIT804J+IHPKsHqyGuSxls
yGTNmdLWawMDUyvptMbDMD7+/55QcWvUtbL5OTuAEP5Rh5eLjhGt9htiE1ZJ6YGpbDtS5R/XS8MC
vVLX4PZuZcDbbDDs/1qGxeWav4SPrvtHxCnXOMsh3uAaDDnTobsQO0yVpus/ihtmwJD7TUTBxXUL
5kdZ5t6ktlhc/9b9TNEN/ZcdD39fc3VODdZs7y6wcqrmd54WBohWWKyTAALF+pSPlA5f4Vh033gn
TeBUlsjo1Sif66iCjHtPIArQFXrOXg8iGrQNNm27pP0d1Gt74edEsZWnUvGK1KBcZHfLIC01fOHK
T2tK0c18bboOU3PzjHbQXcJjyvivqqZ3HkhzKZumvQEbOo5U1TWfwpFLs5v37SrKkjZhDsLb9TV0
u5X9cS5YmBZSfZDVYGSzyxMzmdmBJuEqFM9gE1LnIH8XswchgqB6wokl6o4PDduLje18txpxBImw
qeDXYQ4xaeyzd2h0JI3k5/Nb0YV4K9jVrvd+5TsP/+m4sC7DVnpQowfS8+OIz91xpTk0EY3TKVr+
TmlRwL7K2UCRzWNP4v19A723f9RbEjHWcNQ3tSn55B9pkjFDepop4i1iTigqRGCHZ5gtPGhcgMrQ
it7r5guNjf0tp9DFqKosmHXCf2yxXPesYO+S8fovhthKClThsLQERHb5XhBK6SDM54KD2I93UjkZ
VjxWadmcrOYR8w1YeEADmTYPkf/onoOvOw7DD1haWInJuOuaNLy8rqBIhrjZJ5bsMSnOJeY5Ycgv
vC3ku5VwxR8YetD9tzCN36+mGqSsmVxHE7WKBU0moU+NanjFaOELSCA6w/QxsWo5UuSqixHjlmQK
TEQkw9F6OBnySKmBrp2dWW30M+Ekdg129HCyXQdLtHTiUr5JzV7ehBLA9flXl7xXZohEKF3GSV7D
2usBsRdgqG0QiTAr0WvtYgL1qaUWdt5fQyoLE8vo3HkY/ZD8j/fV/1IZ5nM6W+RdP/iOFj/qdGpY
OtbOR9GKFRt9s1pgNiJDJc2SaaJJ18noarfoVtksNyTPCLNh2WvWcIUB6hCgmpleL+hneRDzFVFr
864OTnsvse42AKft1pdsoaAVGfknykil8yxPbveiyLLN6QzUNApWNjY1HtDvW3qvO87XRdG9j9eg
EyGDFBMaF4rWXUu2rzsnmibxKV4SVgabq1FclNjLVolXJo1kg6KpZyrk7qc9aXz3xx0dJu6gLPa9
/pkHTbIbBlC85QknwAS4jCXyLQiGEi3LiaXbcHhdaVchTGB/d/8YaYHxOcCpQAyYBEMYMETj6Sko
OwZ0akksxiJFwChIcjXHBpay0OzDtSuLqNsEKrFcgleb8nOrUlsvBFlVnLn2wWNla1uHLi4zxW0k
jhw10rYLlNJwuZCrBYImMuqa3DVqlLOelhhaXS//3eW5GdEBaz+2T4jF1zD/MTiyiTzSnMvkio97
csv4+ooX2HctIQsKFTQNpbp7v3wvEZm7oqVJLp3BNo83VfMNRf/4mrHf4KGTtNUqWzA+SKxti9Lk
31D0g37auzk+2UXqwpTfsYWaQSK3XEzCYXcYFX89MbwADWRqxzz/6uylhx1HaAaLAMbMpFawFc8D
LyzUcgv8kExQsSRB/5onpQAs4HSSYsgFniVuHLsFDINUicS65FDoKpttbcbygUQMJernYfA6mNg6
3eCZ+h9u4s1TO1KM5g6bvS0NShk4txUHSSFMX+Zs46iNqClW7J2NgfRzrLw3qGeSNgTBjg9U2s5k
jy3mtnt9+m31gu/5vI07uYAnrgyyYcM8R9Z1nNx3bt50gDGzfuECwi/B6mLwDnA8QO5CsdTMrKW7
c2iMACt2H01rK7pt9RnN/ZPS4ECila1eIKfG3WFMKwRvtNkgI4JJmxRf1s4mgsgrAjONq5YU/m9z
GVZhBVt40hyuaoO/jbJXYarzOgHuFxCqG5ZhSnWen5jxnMeZJGb07eOTYgHjYlPekDItwREGSc9n
wTmOf3iwZ2vETHvxGJMTbEwLY0Vstpw+qPtO9qWQOEu9G/jq6NzxHrp3ePq00DWRUKO9ibhEXVQn
Ieo1f+37mgVBzkLUdcf8Y5qFi1kSkRjwIcyWhFTSeNEd8TrCF9kEM27kx8+zjurjkC/dS4RncD5/
2UJx+EEp2SFJh+pda8LdpEfTJ2IpqU3NaUojaKF2Jr6PbxFDG1OsrIavotd+VT7R3ev31yj19F/O
yfVDJ98+XS0lHhgpOfz5t3vWa/cHz/8TY0eNo9HKFTYVjGne1TFpGWKk4AXjORKfMz972vGPbvN7
QKAuokH6KGCfXLJB9EKJTa4JoTw+nSkBpmLoO9uFORXE5flc2St/H+jYTHFAgVlb6wWpIgkj8dfu
8W6kcirgu38Ewf5kiecSjaz5Hs1P6xq0VYGXu0zCowAh2zEKAZcMzVVJX7EQo6JJJ/Np1rdaBsq9
ySqnt4iChn6z4y31hgw/mHTHDoziFExJIoS/aW1z4LYlslrJFBqSxStDOSuawkJkbMCe1hIpr99C
Lu5QODC2/jF8p/A9v3vO9JtdSDdsa301NMNwdrjtwTsMjpxaFodzBxRw2r4ta+Rr495k4lvuyFm/
uCPMy8IlNn06Z7dgYgD+i4nuv9dULcls2nzJpph5VLumCaNZFqHg4fbZH7hiScp10eXkA6S76Yji
+OjDuYBKWS4jyYAmwBfS4PQllcM4LnnNWIdCXoKlrLE1yhGA/lNoWnooDXFJYKYhZ1lVSYWDD6x4
8ou5t7qZUJ1UvqYe6S+WLDLHp22KkgUZebGViiFKwNW57/j4ykAO+4hWruNcCP2xmmpp179GsQYv
5Xhzruzv84KPCM245moD2yPZnNn1/58yF8adEEzTNQzUlV0+aNKLDRRVGxPo817Fxh50QsrPWbaj
8sKkRT6xZayCAE9F0kMRKXyI8YVGMcOtOv6F5HLY2sHBjIr5C8zHYoVjF/uGEFAGWQuXfNbp4cVt
dmcFQYRG/w01tT94VxehJC+bAdAJiYM9u4H11OBZQ0YB07nnAmZL+i2USaMkQk/Bdf9y7t+cBhBD
fIyuAZpYuz+fEM6gtw9SBCB7e8ErlxzgKbls669288Iwnios2Gl0lPfnJgbXMX+yJ3yX8NvnFf9k
LFi9oNKmpz8D6MgjclH/o7+8CN99RhGvLue1qINGMuv4a2B/LjX3GiOR63zyLjONU+7ivUXqrMPh
8yNUMvom6eAwn+3tZb3jGHPg9xb+HmYScuCQPT/7NfWyMTs9ca0y3ZGLdBjAJZ0NDvpg3ilKG5VV
ex1wt5Flkm4uNGju/yGo56X32V7ZL0xi2FqlgHjjXcp+aRj7SyKjj6AL+rpABW0pR63RSJyl0qEm
JcQCq17/h7uDiOCoTbgMiF1zfqz4oe5QkO0OM0UKfkMnobqyoFX4q5kxjFbR6yL66UkuXnXS13z8
6fywCg1D8futstk3AWW42L1GjzPGkQL3ObnTAEnQzYMHMLsfC8HPfERNvHYjGQtTnkZvM55/pLT7
HoBrRm2vmNG7L/0+GN6QvK8YSSHr/fhBEGC1aoXYjEBpbHVtx29GAECt8/ZifbIVWW4iu9ryEvqe
V3MFaPYyzZD7RUX/yEt9NibnMedqIo/k41PHfUcy5gNKyLOgtu5++FnGzYkOPukedohUmPWtgss7
/mY7rHnf7WJcE67xFKh0p/QxtQQB9r/ymUbcW0Jw/4lN4RgFzjURhvhAoJQYJ/AxZCa7M2RP9zdU
zlrRflXGtYptAeN19+Dold59Snp+r1QOLzjdNYK+RrmdHIPJ/BY+yUJc3mkWvgk/wY5i1mbHpPyV
VP9rO9Z/dEFZ2gTBsEM1agIHhqyklk2O2yRm9jo5cI1wv4x6B0SSl2pNNT1y28sHrAIm9KaVj7Oi
a71DePvq70rrGQ3mnLFpfxLi8ijpezy470INSHEHg3Kse53hrYXljStJnREMNcW/HmYuF94hMO96
e9lCgWX/xJiwiDKh8HzmOdFAhAIPDB3LabT8+GtvqAqbWokxjB0BFiZYLYUu0ZzRsWjFHxYWstkp
BdIjLbak42zVXcsiw8hJ88cZUP6Xz85l2DlbXKrorKwUtzB5GVjaqLqr/E5iw03QW+UcMI20pTUW
2VK9k2P6PcMv7wBrqGhcE1yl5fuN0P/s+UZI3LRpf1pS2o7EFsxngG8sYB/C4cTDuCNmjFZxW/qj
GhbmM0H95Z4ZEOdicJePZmYS+BUxhA6PFWqkreVOCcHdVqy6A3e8jmPNMUqtT2KgDcvIzF/tUcc8
sKlFLsWEG8V559wA26BmMs49R4qKv4yOeQQOQ14pA+RDNYm0wzN+zjpPhKuH5nYMiRMYYYmg4WOC
ZtD0ibNZudfX40fTdOBjw9V/baOgfKLgGT4XF5+0ao2rc9q16l9EJ3Dv48TIj4j8ZspItI4oWDX1
Skvy+Y9wXgO7lPcyIsWUvkoksScJNockb2O5wdpQJ0VuH3TGMNsj9qYtqVricfiKEcSfgxDwfPW3
LVRz2hm8Mbvvty4jyazAMTG5ULuItfz4JaqgqQNcfseYBxIz+L9Br11inE58WLqpateZHlHdF+jJ
jtdyENQ8RxxjmTxUKV9kRaapRzJtkFIBYH0ZcZDQgjwFSkJFADaj45wtBnpL5LdoZFa3l26qggai
os/Zi7nKacBcIcp580nSjMJJn3znJfI6WMnEIhjVNpwYhXEvzJCIsM4pLwIVRLXVGHfnTFUZsS5M
SnJVtGW4UBRfKjKOLnW8dX57pHcyvYhZL0KzPtmyrw28+cAiJ18gryjXea4Rj8cS/fVPhiDGacbI
+gBpKRm6L/KwbaRd7Oz81LF/Cb/S1xkiWYTthpJmL+6v3FdApOgGDJxflBqx4qG6GmeGPDcGtGMn
hRv2FyJllugd66rp8JEbGYjHiX3e1DKC9J2Bcd5jlbT6IM3Gd5fbgAf38OhNKjow05KerJ5TBpxU
K3w2RFi2D0MnJlyb19iWZRxZepJGagoHoDoGZKgKSt1VgjRI5Khh3PjbZVmvnuBYOfb4AgWyIvcF
LyFdfkLNhGBkfLn90UkFFghWF4k1rzv+7+WwPH5myqmBGHays6UCmLuDslum8KC+sHJB7/vw6F9x
b7pE6r95RlWblrZBOMkXQ/tXlc/kpk8lxZm0lPsEVqYRNjkhmJzL9W3HSqQ73spUxDPZxxnG3kYz
O/WsOMiQTyDQHP/QQqDbbRbtYbYOy6Snz/Hs9qIwwaay8tnXS0hTqmirDEqhDp1+RbPGJ9OXppn8
RLRlUEEsVl4H+IsNEipK/viRRv7jItBwARX6MJtEXGgXkzwx1T5cptn4KIKB+/tgzIrLvy/6RzPz
tt5yukYhupOyTCvkFM28gh+fCYubF0ta57CgplF/10e5DnkiF73WDQY9buZrbXeTNZ5wnmOp8Laf
3XWwVe7KAvoOVW/5hS9qivHsZV88U0mMCFpCloLk36RjMbhqAUCugPoducplqZOPgM5mkiyfAjWj
n2rW3FPz9hmwSuikUHfQElbOhENGOZnKdY+HA3xworfUQRLjbIawrEbehytNXlqNmN7qydy6I9zs
urADNG4sj/C7upXaH7ygfARtCKGkdc4l9AkzUrJ5uQUt9fhW5cfLkiPLk2yIZzTRt7SL6GsQNWJo
FJaB3jhCjg7AWftHKhivTwG3/N0H+3YY9IKW0eRLs5595+kibrWl/T4/an3yDQUXHcznXUYTm4Ej
zWvIMmkpeigt82aNgpBjiJV9MmjohTtNmjZmXDFckdKK0xlu1WKPld9wjoIZgUUqoUjDP4Xn4ANR
kL1WJQigtmniXzxb5jgDcv9qYsm9mIkazRVrimvfoMLnKUGYknZw1EUNjhxk617Gv1xCpT1FhElt
qZPAJPA8yL22gtsmeSSLBPJ1J5A41jyaw3BfdjwrgWl0yyfjP+QQ/C/q2e8iQD9Z7b83DVj7WxxN
F8ZwW/GopliJWC0EvERsM0qW6B3txSLATm9BTs3IV/Kg2uXc/x0Asj9vcUT4PGGF4DMKhafZM+EX
rymYzqtVP0SBhELKUY7MdJwGlJfvsUK6yC01iUcv5pzx1Ku68zp2Z2uANgRswIAo1qd6x/i2ZCcZ
tK6hJd6SRIQRXy6PvpR0fhUeP4OlFIlSARVYfV/E9wtm9nU9uosDqgvCWApFpciLOn6zgMXJUxPr
SwmWQTueCuxjcb+DOw3tIWZ+tZQfpGcsOaWBTMkVWFJFMhAGbwOHLoPvHG3OHNrGAIY6aymUvfWg
zObAFNprC0lraUg9/KntSOXw6eVn+jSiEaIGj6hFZwlu1r13xa/+ordo7rSRxPzWXjDR8wLRvTz9
FfL55j0mWgBfR6Cb8c09HIoVVPUMUoK1bK1RJxvohiR8ctE8MNYHO+t8LoBkhW9ffLVkFgaOQKa1
wTiZHtkUqPyRmVmEoUfOR0J/zW2eAevyFLJ+4KJEqMnkEVTmrFssWv/pL9770NGPt4f9uepYsxta
Pw+HyfqpoIeOU4KyRKyrhneane9TNUGIKkdg8rvCKDQSxKjyP64NeUd0xUCygpqd3Q2SAwUM2ZoH
+iZhSU6LFETlBZ1DUQB3cSdU8qdUGA9A5L9t1VqcDb34o3d7RfZaVwBZ2BTRn847qsgaWZroeoJY
3gvyjQaMcSly4KZguOkECZ4MfgZqNTSyG45LbJimpnBKSqdln4or9RSiwccNENQKo+F0zcaeQ2vh
eZYuf0LrTMj/0+MjUzFkqcMYaBuRcuwaVrRGBIPmRcrafk/Oz8PrIIcHD0ncMb7kKI4odMypENf/
1sd2MSJImae7dNHkGMeDTayewFjBOdOOTu9q2jPyvbm8z0ow84D17ljuWxZkm29q2fMeAiAg4U0Z
7tsDgAKmDWTlr/+koKLM7NaSqjyturukBSkkj6CXNrESNQUWn/LrqvM8paMh4yWuK2GKBDVrgCNP
vRN+EHJvkNTT/8dMdjVGcJC0x5Pmq127IRLnVbQH6f0yweHcXnmDmBJmbWW9sxzCpE3GJCI2bY90
VqOkeJzRw1hTimZ5maicqrRECwDWzge4h+oi70komr049aasWaBvJbfnUsDXAlZmRKc92Eo4sn/0
mQ/K0B/z1joBUECgMVXP04IQhIHYsOXMzKgUOG/qcwYdL/qEHTy9wEzZM4jBn/eqSAc+H+PZD1hY
0U4uMJhcRrvJ2YyUeE8oRUOxtQSTuwfo9U+oxrzq+peyfJn9jM8ATNY4aIErnX9l6ca2adApDGw5
TWtmXGBU7CpXpNJaBr0TeLyn3+gBKr3zM9Hlt0gioklFTaggMyoaIqex2c0iOn8DNhiL992lFFfQ
lSpbUXyTP3WHBgQDzb8gaNEnWyxs0wW4dICapV3aDuH6/hPb3czgTyx5fDAINg1RfuJprstxnd3M
srMRshVck2+c1SUyyZGZSmasP1sbv3bPb6NEqyZwr2etwseMMnkNM4Tczh6DkeLHoFDdGSGeZa3f
71Afr7YC8tEE0vRsaUygHxk5JYawuERUqFdeZG7bU51K6dn4yifsyLMEfGQQR+nHTtHi922UYOFp
dmc6WCOBVYuPHOjExsNpRsqT194bNOTqZdEGwtyoeZ/il8S2Odf+s59yYIxdpD7c6I3j525vSFfT
bo+otlEyjPrh7g9BuZmF4aRYBbOG4KPMJWlLVpxMqcgdAIEPH9OO5qEx6rKuPj686kNwYeQrZMhU
9HzIN+06PTPd6VPS+68mJc168skPT6nyQ+MWZps5oAnrg+OSjQrUIYFdiE+r06KRthr7xozH5gMB
f9oWuXWdNwCZe1IMDp2LjCdi5qjyIqLnWo97FVb6EUGc+LH13xH6xx8bdSSAOfAnkw3XVimpJXel
hH7ml5PWpz8A0740tGADBabz30tzSucgI3/uEqrGAXTM/xFQpLyzx6+6icXvtqVB94/GuYnoaA/9
ygo3sJfW1NJHNNCOeBLTcBQTbKPCoZ6wqRE7IKSaGmXyopnzHibwNUeUWzcbhlDqoUSfA+xFOWj6
1dNzIjbOK40kGXRffcM1rp3WqUUhlWLbLQB7ZYBjmyiTG2BYV/InG6VlS6OA3bfRInmwC7rYhon6
+QOpuwyFRkohfbd7IMzirNb8tk50xHTTH7GtSvFG9wDGoV+IQ2Z9A6xJOD1/QKa6gGS8EmYfEG3d
xbLMVfehtoHq+2VBCnB4zIasOG2+LSEqrepICf49B29tJnnv5f4kkGq2tTH0hCVqmj0CpNZvHlqb
oPDnvo/pCml7Q74iWyW2ipQ5n9vAiVzQp5en+32jgok1POLs9DXhf/GNLGzQgG4dckw4ai1f1eBq
bhR7HTQUrObDvtbXItqS4yd8gkopF9iLeDXjVpwc6HAP+jXCVYstjZs95K92DfmNXvSGWhcnuSpj
ZiajE/SSpXrvIOVo9WXSX3YtOB0gEjykePgogMjAiBW+ei2SgcCvwHm6CpWwrZX0WRyO+9ILuU16
HKBuD20RMwdRG14GrjqTPOEsZuY7ewNbYJSsTKduds0iPpbyCIRe5PRLismyuaMyU7WT/VMXGhUF
RTlxPiB5delbhVlTG4y3d3yZgr3XlIjECQHzg/HSSy8F+SeTv4Xym45dMOmVlz1CMr7MIZfxuUIT
NL4TwtwaSBvomd0uTNQG49tcCQEqOV13rr2HKm3CtRsoNu8FET43OTBhXuRJFMKNTw1MlIhsuzEq
eaWRwo1aSWOXthDmXvRjEFynvofFYOg/d0v02OKLk3k2apDiWkyqp2VA9TLOOsoLv9XfO8v6ftcT
V6t2FkxC0GyehHMYcvpkJSAnGOl8bcmMaFb/7hBKkiWWN+gZXbHddE5AEYHHD2EolIVJkeJV9WQ/
LYcxlmJuJMx+d2PVdCDQUCMx4JpepC7mFpFu/tTQD7gCaDcXM2ujRyRess2eDRANyvabBFcAFpfS
MiSjM6svlzeHq/G1y2InJnguDyMZcJ+cdWBHoC+P3qKYcajjm8euTPCDYkIRtl4idHD4OoGe1y0y
2s5kFKkhevLOultd4Iw32b124rg8VLe8SSIGrGHGtofBfuGXAaK1ed4T49tF/K4biUwXtzR08Gqf
UClI47pzFf0+YZEppftxIEWj6pDXqWWfIuKTzKSQhsouDICG5i7dXiS2YXEanVuKbnf3LPw4t9X6
F5SkY3iWvPcAvtCJK3yGv49UXlPinSpdaSBfYogxe6z1ma1+FdcWfHUlmRs8qeK38iV4IoZ19C3u
gMbAJpeT4WhnE2p61QaWafi6VBJFU9kALawXHyRq6iZtG9J2AnE8yC8lLORBxNKhZG16nu/+TTar
AULkcUOXoyLjctZ5REssr7GhI4skmZ2UxMb5rKIP2eQmm/SffVd/xMHZ5EQmCi0tXXvGuREINK58
kQwXIPKSzanljab/VUZNgCT5IrJLJTNkJUFiAFeV8ZJYbtAfbvXhpCuTZodzX9qPcnZsf9CYA2S1
/wmcTWf0t1NVt2q3Fi02z32faK9+2pEfgcG1M0EdNZhG4lwP9veQKJzH7b4w7/gu2yHXqmWQuURQ
P5tT53qKg44os8MqdgP0K5aeY0NyYWeFTiFHgxicxMHkb2D2Rhd8ag6T+9czieKG3yu7bS8az65f
8GJhl6QAE402yvE8zGxY9GOWuhQLQJ8XBMin3EtJeUP0MJip4h4/+W2Y+CMitY6cHIEHBWapfZPV
hkmpOXmLEAicLoIRbEz1LJIXI7ki3bRC7ygoX0yk6HFAcMUalJVGaRMOtJJaf69MNUdPlhdFP5w9
bFMerGCqWpBUdqwh8oVPAmJTM9e+XcXW16MNjq69RGo8UZngfEQ3ar1hNN00niTrTrE1n53kDhFa
fXsScqGmpFTliAMNVdPenccaart+YXhoRP4MKhF91sYtC2a2QoN26Br0rK1+OaNBC8WvKRUqrf4p
iGFTNc1fbrYDuFb4fYXUnPQYQBY0dG9YNWFtknr42ZkG/L3QFoszLBK6Ue028sAhT38ggwzIqFpn
bSjmxyuf3smw1Tv3i9t7Uq93cKzmSv9pXIseBQkVw78H1KnRUoq/Sefl/6btxOhN9PdOSuw0GjGR
TNRfftd2wTj3pHS6sGF8PvH9XOW+bjPPvNxnuR6Emh0TAt1O+kdH1HVLD4yDLvEJPkiQ0lWzmFjP
tnfHyYZsI/TYR7DgSuZPX58wiCHqbOtVbbgwrd/FqyvgwKcqebusvRXnBidVGVp2pZz+TemnI6Ai
r2Wo92pLfMAsgU+hT3LKcSuLImgGj2twaFxQZlhEhtK+0/R7gNiT54EkzM2UbKMY4I044mQnCPBj
CeGx6ojShXFzMgeMbA9Gngx5Bj+qKQvZQQGj/EVidS0DZOEnXZjvvUFeJQb+FFPjM8SWxEkXtzDb
yF2ts4ieRiDyI0RObZtFNz3SXcV151hy7I+o9aGaEXJG2lrpbwVa57R0ykeceLI66cwclEPPXkp8
Fopjfo2ybWf+EcBXK+wdTjEKmiTyGo8KyGEWyES/GX5wGIevOyVJ9Dj50MmnecmGL4v2w6+Da7Hr
/1n82XWv2a8yg+Fa5UcjHZs6+1ogw2X5u4Q0uEIcrMkiYnwAulUoRfivJ6Dhl+GmNM8MNdVau2uI
ZXBcHLxd5mbjLBH6Kfq2TwFVgQvov1MN71fu5LNPQCNwmH2wHgiU09ay6LRrodlhnX+nl2WCszgg
CdRPEVgwZgbWQYS5j8IiNSyQrPdoJzKGZvt6httBIclNsMMbs/HC1Ox67XnQw2c7kMNtVDvCzB6C
mw7+ZLtpWaH0zS8jrr1fKY6+vnl+A1LDWh5IDX2U5cBEf0HFqDDzBaVU9Kkmq0twU31vJ2TI9BJT
QUdd2uVOaIeUqRJ6+k+tnFMa6L3skUno0WV2+ydPWDo7T1UYe50rZHC9ORVS4nhNP40PfXw89JAx
oeb1UA5xbVycqbaZTyeE3DOzONXe3DH6MLkpEsb1RizfsNsdpCeV0tX7ErO8enKx+wMYPm3XbxtV
hiq6ZeWpK4qUWQLeY7ie4rS5ob9nCYej/A1C3anVUVD6xTw77KjaZhJTZgIZf790DO1GXfq54wyA
0kakU2kJVzY6YPPf5jOhToXauQDxH0UZZwVt81wGbipXPmX8NbyhlHb4I+V+2BKuGjPg2W0LNpI2
b5KVMUlNLMNQG2/WguDii8b1kw/Ts1xEfD+uUtxgwSBQVIt05FMbTYOTqTrewfmbuTocObZCTeca
47tuW5F0RWrdklrTl8CO4S+s7iC0VyqpUxeFPxDdnuxj6qghmuknEl6TlA8xB2jMlaeboShRnPTZ
6iUEtLl0bWZco6fj/0lU3RwXT1GRgY4P+0//LRIORpmjbvdNqpoxfE6+dCLyEJz3U3DCE34tMnVT
3JfoTknoXW32ICyS47INGlSdgsDhXCFqcYe/4EmaYYBiYn23sn/SmBknGNecfXqcGN6OgHCs0KJJ
n2QGhzOhu033IRMAN8P+cG69UrLiOk124I2WnsDfhNlTDamCURFlb389IhgzukREXYMhrrzSkEzE
1TN1NlP9mfjs3sY/yY6fGAdpqdKVChtmvpRqRbidy/xVVOYaSmdGbUZ/SCWJ1Wo0/Gt6ab8sB50Q
7FWQnZtnhOPz9HrpEAnTw8YPlsidfVhrqXXP4uprSKsQW/WkWYxqlEW8Acvc+myO7IQVb29K5Rh0
hN9drag1/0fpnZN/g2UXpdwTzwfjJP5+fHjgeQKYTyL12N8JxKcmtNjE+lrW1dfcYav80f+Add/J
gf1InGYINJhXbHNOhZXUrrTeqxrpUNdsqiM68FV06w61EFsjPpRjqx5UwVIvLESOECBxiJ8yr3Cl
Glg0x7M3warpjJJ2ACuic2MoDLI62rvyT/RpFC6thualSGbpSCDI9iQd0Ggpzvv56IXer0BMUtqL
z50RfAXG/I3gaOeGbc6dzE8F/zaeV4xk9F7bHy0PYRyGuo2iBLuVl2bBzfLd82F9ooXnJbYQ59S2
9Hl8e6aD19xqzhK1zgUrSjsCcoySlw8ITdyib62qr7WKDpTni/LQdhd+UzXOsSeYAEoajshs8iph
cpTP6ESxGXMJCxyUOyD+gYmX0YEMkD6Zgsc6B/OAFfCussWXTAFt6zeztI6dEieW2rpuYz/ua1If
i3QwjfZnRqq/VmUFWWwN1XdjomI9rY20PG2HSYXGr5hCoIvxXmd6svM36E942qVjWyjjyGYlsS6+
QrVqGwNO6t60v+MIJhEp+RxpFJcb9mZhJk8+XCuiJ+2jcL8no0q3PYNmdG1DYC8hEC7WCvCMQRq7
esvOINDIXMSrmoUtag+MSj2T64w/FejB133QcmDp8b931Oi5bB0usgu5PYmaDffevVztYInRLj16
I4w1FjwhCzDz8nJhg7yPPaOogReDL8u7HWRToEPkL9kq1kgyVn9+cg6bYFpIfxB4c8Bc1XRs/TDo
Mo8eAsHk+ZVLuSGL/VAKgXynHnu0+Sz2dT7pirkDaCaHmU0EblHUbBC+z0lWl509x/4kb1AJTL0l
vJcCSDxvs0Ij5OgoxCYOA6++wN9yFOtQcpw7O7l8wr07RG6Hcrsfcudl5nMzy4JWPm8gUEPYW8Gr
BBb9BPx1uRrFKPoO0KomUQWJroRLnW2LHJG+eE4ybztdP30poMSwmvUcYvPfi56hIYW1ODNmfjbp
zDCxBZ/5dMXW04c5efaV/9HWr7UaYqv72ARTyheoc6GvC+VIDIX/JLXMYH0rtfrmUya1cbCBf8up
qtBJG+oAfJWzBV4khgQWEePYaLD4K0Wd5nlIEA+LjsMgYW4TwmZkCSA+m90aLz4xNA5N4gvAgp/d
ctub97ZBoOtCHH2IofbhSPWu5p4n+lV4DL1+AbPRUou4/NZkIOfYUirmjDnHttrKpo7XUMkCNjNV
NJBfTv5UDaYfAPZ2j9lw7wDt9VDFB5dS97heMh8Ka9fKFf77Tw62Md468vy/ZvydK3xRTk4O2cw0
wNmB4gITPLPn1nCy1xLkUKS5a4GKB6Iq+6wUVwSfNs+UeUvBXZFz35mXf/aaqwXJY6KjJwdhsaz1
7dwgL0KFGXdE8n3HE2eA665aqkes9brMDwBd3WNUDZ4YzspSqTKpWobCHLbHFF2EwkGPzXauTH/L
XZwCzCZFugZoXT/+VElX5GGVGB1JOUwY4bSVluvEZHa477FyLncAdB4jWbDlWq8KZ1AXzXHfJH7B
HWnmi56cafhgwCoVvj2mgc/XOpa9oEXihlKAeRYoyK5VfXMbeCcmBOlcFhf3WL8h7xE/KxujnkHt
YgG2AbuBJd3JBu/7IZl4RmGf1YJ/CrsMlDtsfpjQdkvVHtKq5PHqimEsp9jSJd8TVvg1Vuj3Mzgo
qkFUoue7Z+hCcKEJUKN9Xv7Ia7PyzoIkrzvZqFL1hX4h0oU5+6+tv6HGHI6y4L3WSrMU+icgASfX
3qAJ5Ek0HX9tt6kYktqJHOUK8BCMZShzBaphoVixyJVyngI1bhVvQnGM64KULTNJ8hHspvJLgnNt
7R2uQYTqIF7Knu7iofysrf8/6Q4385TBDHpkVuwP1hE+dkdk1bGMPMnH5mjWInv8kUA5gbO7tVj7
ebvvgQ92ThKaHUT1Vi+Nbj+pSdnvphcwBGtqLgDnVxm9RAqlVlugREHYhriuHdx12R1ki4rX6QdN
06sCvtkGBVU23yDD1yDIiSqTKs25MtmoCFMvvJa1g/DIjanJq7RyQNNSfGaZYcYSA75zpVCxJ08p
S7vRI6IymPppNVWa1eTYbtPUcDv0TK0Fansvns7O3lMhZ1m+vl5ad+MX9QO735BNx7smu+hrgXpH
+YK8Lz85KGYG/MKQQ//0+kMXFdayfWDk3iMd3OblU/f9UB7TKJA3YPhZ2uOS96GtDxeTVORqmlyA
Da+RhGTCwSYr8XETOj3XMfqmYK6Qm+U1jfnL0x9hYMfopLCoaY+uPe6aBk+SUFI5Kkkm0wBv8wiy
1rtcAq3wLrjePHM/XGy/Zg49kfIfocyNKB9mRyyjfdvlm6d1dfvUlDp/+MfUMvwXD5LPmlgsF1i5
FN+9oq0P/Cbt5aKODFetKKYc/XYB8QYu9vNppmOBCXDa6bYgHCJZu5jzkBiiTmfCfSj5HROg4hjb
ALtsMWsh7Akhl8oV3QTDvVJ5J4PAJsn3OpOO6WlbIfS4k93L2eVVEUE1B2sX7d/o1xlsg49RBYb5
oUm9o5cTFIm87WqIN0BSX5ktycL9DwO+TjZ0yzBIYu2n0Wwe9Spwb5R6dGonysn6KSZhpyLrpAVs
lPtIQDSo/N/HCYwBkAj1bJMPDmiOUZlJfN1DirqifsoT7A5VMwjBlES/EpXsvZQ6xMHDcAK27Bpu
FqJieKLGkAbnwS6hUy6/zj+Z1JgTr/DhuIyUjAux3mZIMx5Jt3slnCkEsaEpJzg+LNeGIA2Njyvy
60MN7YPLqSbqV8infUbYk0rCV7AkEiJoa6UHNwp0XsOQ6hOYtB2O2NfMbDus8M8NqxVISmaRfNOi
1e1mGuuoqnx6erjx/gUbtruCOOXs/ZKLbUSyf0Nt7VchcN74cocY/0VJq0QhlQ1mUy+WGYtYtEAU
Ke1EY1bnkmGG1ONBkyPBVipuATprPA7SMQdLCN2q7p178Fv2z22mJV1fGIotzzYxWPfeD4fOtbX6
HFnl/AFZeHr74M1HdN2HFq9a2H7sN/bmnYjd6qSrOE7nr73SWSJexboK6kT7EReHUJeo93Dduola
VcD5o+VMW8wB5D+IbXaWkrm+j7gj0gi8nXgyeMiaJiL0Lrfqsw+yYDxyre5LFqr4dIixLopt6BdN
0a5hHbm2t+t6ByAhx3tR4QhqUvr7/BGdy70rqJJIjdSTgO8E3O1GcSxvByKinNNSomYSPzNoXcmT
Jk9ublWs3F+248+u+z9t7TZn+EwxUGrFOZ6wOf35bEF4z1Glijj8rA8l9WBSxgt5GPuzOfr3jV30
5RLkZp770Pf2J5oi55Yf5WwyBboM++rYpuVQn9kE9wfAOpz0Q2JnPFb/iqkWaEyM/hK75SCzaCs5
fyQOHeKi6QZQ7p2JAFHMIajyt/DNzPCAPF/7Q9YdCkBqsLMYGA39luYUyAgeEzbpCBKIlRZfNhF5
hcE1DnK5PoLWYsFsxkx4PBLJVcmjTLP7k6nr51DY1KShslqFRn9XA7LWoroEHOLCswnPjT4ogpQH
3K7HdwUA4zPlu/9aVDgqlUrCbapQpe6HpCUdFztM5RGvZ4NE2KZfNQEzHq275bKT1OyFizY/z+pd
d9RJO6a226B/AALSOKH4Botr0WE4BLDWinRlCJuPzxQZM6f1uW93jf5USquEnq/WJr7Gl6jQVG3Z
ICDZvkInYEuqjLks/JH+7C2OlIISxbXLEF4FvTMyG6bv+jAarjW3ZL18QBOjSQQUCC/ZBxhl4uh2
smJmWxVTNIBX1uiaHgAlGhEnnLU2dGvuOBbfkJQU65utQ9PNhHpwosDZlgAlKXRTJ5xDObuOi7tx
E8E7//GskXOIRvoEfT4vGu9HMItoqUu0/ElRwob/URZwc6Oo/n6Xv9PgJLQONxQWbIVWh1IsFvP6
a6eSfn0HS+fd3mYpEY7oUkwbduH75vE9qbvVZrbkaBd+0Z+DQAmz58VmP0VkundamCkiJ/Aj/7d0
0EP5qMDRulGjpSD9NdzvI21G7jdAF+2GPaHfw17Yl7lrjaDBk6aWfV+XLtJRsN/5RlC8tKeMbcwh
ZbFJ3bDQ/f6teuWw6OSL139XDDVbl7AGPuxtZTXE1nwJkq47nBaBbTSRbp/zena+zNJf78q17IZn
HdRK4HB0MVg87ONmAXYQn9J5QGS7PEkL1p1VtWyqmqOe1hY+A5HQ7kO0xbhMemmXSwgmNJK8NS3d
XWTmYUHOEguYmCWaC8rRGZMzmf3Jon+PQnVg9mLgATQXahL5HzpDAvxWBn82H1aNfyxOxBdf+y0f
6930HndFDJhMlgGbcHuznNDn7pGDgz2ndHK5pGU0PidcDwwsOrUC1uNc1IRve6m9NVUI88GCuEty
G/p090/A0qA0y/Otrpx9QKgtwz968pM96Er7biRZwJAjWLCrCaQq5uBEp0Wq1vq1uUbNQbkmSWcU
Iqzvc5XDZ6dG7zGyJN7VHkLY3mOXpdr6G/7yKSyLe/YQ6JpbgfAYgWY6MXN5zjD/fbOhcrbo0Y50
+mCG98ih3//Lql9ID2wOWIVreoXQRRBm3YtfY3Zf1ScCToZ8c00GYNCZi+ask+NOMRecJmXNLcfC
HpzoG7nwKiDGzMdSkC8fs/uuLQRkfZ12FWHTyjEcbiN7ouTjhQ5EnROX1ESvygvOKaEGKBbt5YAG
PvcJxVxfpeE764T84rvwyooOhiXx4SDh8j5qyl/g5YcUvr4Pf2tgzJ841eJq5xDYOLv0UzpcobFx
aD1U6rzaomD3w+z32CuJ2hUvPl9GXCJvqjMzTKRU6UkGZZHO7Qr4YomQw9wBvOraUPyMvYo63ZKp
X2p7v+qxwPSa9YK4C5HpyZ+64lWgcZMNGdiurDVIPUZPoYsfIu6f/0dOeclcpKHb+ViK8NRt3ITo
Z8Y0FhJLKofevP2ZQxk5XVbgM7KAspbeQ9AwZ0uPXJUx5PD70riun2KxaBVjuRtpg1YeA/P2hSzS
ua+ql4I1Z3fO5X6Z4rKl5VSP7OUktNPwYsYkaA4B/sT2dp1nDDxjZ9S9ljwkjfYPnnPP3VLd4+dT
3VOhR8RLX2wNf7BZLK5HI0kIAhQbi+SdU7wQFRs2CIm5+fBAlzhNqrPA8gsuLcr/2YGmFV2+2aW6
gypWOI/FkqfMrKWT/Em8zhEcwN3PDsE4tZ0OobYOwC+THwySff2vHNEKGtJG2f3aCqR+Ay/cCFbS
AiNUu/X3c9Qly/23y9EKrFFFHpn1hvpjQw/IGufbQnWKr8aahFzqulvt4ZkkxukkOUsiOdudcHkc
6pmm2C2bdVF8vj5wUlR5UiUEG3ouvfCgApQs1k9DA7wxwLbXMJHmjttt7/h9o6nbbxQv6DzEQQ7+
A6YremvMMjSXp88IYJX8Q3RENuEsJOXztrH9tXZX1DRUi0dOdNceEzGGM6ezfc7SnSQl111d5WJS
xpX8WjMi2ylb2SgEunEYJSTQZxBg+AcVBkIqH2R2MFp+py1vOC6NmfIHevlpWl00Ah/MF5PglEU7
LKANObfcpEH/tl3K6Y6ooGKJL8B4ujCZ0OOLqoaYhkr2pnISDd9IVTaY/BFAUUZuEX2oKPijSuLM
S8ndQvFem2Imp+EAGy9vuN9xmLEZ8dZ81VzJ6LtAFOkOSQ+V2xD9wGV6eczoN+6bASTBqSZdHN6S
3ccHSv4JZmPJu55t9z5HGSl3X+SvD365lWtpzWRw5ojI6ZhH3SHBS9NC5tjYmv5uj+Po3EYNVmSP
iKrS/bs4BAZw9glrJuDot4kqIOr785qlS5lx7eNli133k5PirghaT/w9oLr/VVgpox7vsaMMebfM
oSQvhFPg2ZRNdszPRA1096DP4r9ikQVfy/abnyCVwLwsmad8QKeYDwT78ihwfIOmKjOjasn1Vv95
9NA+frd3wdHJt5u/fwA9O5mfI5g8JNyUQktzBcRCPP7U/WObOomcU2vkol1YQfvmz2g5lqv1BL3+
+oNWae5Drf9dedqQZfCUK5f04sbWNKV/xDTRQxXm17AoBZ3lne4xcnnF4/+IKHviyNlRY/cRqGD5
WFtbcRtFZMVvAWKb3rconuXuz/4G9njyrTG3CIuVCiK7Bz/DLbC/yJQtqzC9hHjrAgjprMinRIRt
ucuSw5si0BYBgd0sXbm7U5Wy6lKsfvtnjoXwdscrXDp+hXi16vD8qQlNHQS3Ony+1FDE6NVKChuw
78GmhKeq0yMMAP5FWxhZSX6JiEKXlUVKyWFP9K0w3ox9338qw1ZqYt+p/NDDwvqcbMa1mV/e+m6S
Pt0avzViueleD7hxdydK1w4sPwnOrTCDmPawcDVEF3pFNCjb3bUp5tEetU3737D9C1hT1wKsTO10
+OyJN3WvNxx/w5vfrwf5OG2nLaDdLKVWChO7Q8XoiKaEgl5PXBJm8n32w429MrviUgyrdcrtHvbo
F+bQepAaq8SUi4wyVd9Ez3G6DpacCu5iLLJrbHA6SVVtrAkZ29ldRYYXY+f1lOJ7CNHjRqGVpZ9i
gMmCsSPyjn1rwteTZNk+dNhzJPEKByg9L+sNsu1UySaz3iNLzEcsg5sdTtYrlEE8h/jU5ySGzxAt
wcqkHBFgvAOKwWlACBcz6JOrEcKc6rV1+kQLn0UOHGf76860wlHefsWzuowx4C6SPmFNNd1sDc9x
aRXiRdNbSfOd12Qk85Cmgpc4l2Rs8XIuAd1g+O+iBDriPjtSRSbud3193fhOa9oJYNi7r8KGD7uD
5P5S9FcLv+6H5J7G4xrjos5YKrJ/fVC1abMc/R3YB1UHsepJrcDgwg6nFoC6dfHPf+FyPuZZlt7O
57chzi5JcLtUsYCyUbHxVjliNyXh4UYdVqJ98Aq3DpObBtiEkH6V0r1O3WguF/5x26LZbBQKW1Lb
p/tCDi18aCpUdPNk51JI7Ay7ZWSXhnc+W0WwM/B4FmPn7//gFvTJds3ZPbLPrc0d10g0z2RebPC0
waynqZbTkaX3f7dRTpbD/styVTO2aipO3qFsQ9gLTD3wxHzl5exFx7Qhql8x5oS3NT0VW+NMlfNB
hTcZ4OuvXY02Pf0aq2rPjnCK4oRM+Ge22aSt4jwN+G78hXzBKdcKl3PqHaJ1jxX8Tg7nMoxufMWr
GvLJQZGiclHKPxskbwHpexlCZ1vLh9LyPkiBDiXU+eaX13YURkNGdD5YreQzOCrgLGDsQcojsz+o
2R9A8bnRsD9A0FwbCRVYlCixZgN1Gw1AJdiwwS2Vxa6vF2M4rJOKVVqgXy7yqpbcijWVp3Trl7MK
HaEbPVmXRlLmnI3+wVDWpXlILw6GEqfda6bcjv/+iYjUXDTO4kHCDqUGBeECslSUwqYc92NBuXlh
UwC/ZIjNegr5v1hVngcE+B/EMMZeqaWipKFep0UaGkTJb1cLuKwY4X9q6V7kmKpc86QOWv6+6LFp
a4FBORB20DoKUAFdqyZEQeiN0Yu6Z7e65a3MeNGwry4MNH3jlpEFC4StaRQlgm/9L8sDxlGmecu+
lC6Y4iyWiATMZ03d3rvRXfcEXpcFySqWkt2YqRMsOthZT4z2FGCvUhV29VBHjdGJ9fG+lSkCAgh/
/DFa2BssC554nILzeGm3o9sieF22cpV/LdYTyz6f1qlMvAoqFqa46SD6hoRQECA8IJkj/RdnOi6h
GHqMJZaA/okJK8ENxj36O965KueXPUREAPFJYDspQ66R7bb3Zwyd30hfRyv4Ha2VT1rAzOS6fUvo
SKe3zhCVWU8Ub+6so0nxR/4Slo8HEMLU1mEF0hL2SYBaNXYvbedCavIyrk/8UvpgWQlkdTRbaWru
TmPKc7CM5HnPp0nqHDmK2Q7zPoFpfx5e2rqmhywe2TRuHN6PO+tXNfFb3Mf38WKBA5Mp8JQX3WwT
rtNjLh529tdJ4rVJy1/ZEJV+GP1bemNMVPdJg8Btkm5xyobsedbg6/M6TQ6SK67wzUJ9YMtyMXaW
maEHTUsMS9HjSFpp4wFNSQflQUsEUYDOi6t+4XxFt71MTY0hZ9L1tImIb1DKrhGnNYYGwnBkmo+n
N1TxjpK2UYNwuBCKDVm597a3ofjZcDWoM4Usw95J0usuXolQEvM5FZZJiWA49fey0EmUx0Ws8mNb
ewdyIPNOxFGkwSLwRgRBl9Ng1GQpJ7ImUxcklGrht6SBUm+0K5a84Qon1qRC8QJlTTIDAN/ZXRH1
2vAj7FXAVgJMAtU0wPt3JKiTXoroxmAm13R6ca5HBT7xaghlLbUrv5GxHXk2NeF6594VR38RnQjG
gxbNHv81DI8Ne1Q1PIcb0Ay9hJOw0KnKJjtFt02Ba1n3uWOUQd6XvRd2f7k2iUOr+O5OZfeBYH1x
wDEo90UHYWKgQczyr8YfZEnNO7tWtCo4br+BtPkE6yoog9kZ2LfBrBNDcX6uklvvy9W/UW4QZPsb
V6YpTXHyEFbbEqgU+D8WdHkwIrzM1Wi1Qt8xC8ZI5zSWoDu1WtopTYl0ByLaPuTxRHVeb2LXGYkd
Qvh+sZ72nYNZno4q29mfcACEavj98k9KTHOy4zAfVakCtBpqTt3cUrI5akqFU/iyBl5e65OQEU1l
rgDqCfUEIPwjmP0cHb7iwJPifzb2IvDBABI3vL5RNSoPDg+03UZNwKINm5CbG2pBIRq+btoK9ERi
BiW647EUKZ4RffwIVDy4oRejjYdvDrTCTxMTQDUCvsUbeijFlx2BymT5jw4NCirA/io82DVT/aL2
HxCpK+hXbqnL5c+yQCVyNo96ZV4kvMxTy+mImUU5imrXeksvhHJWanxHJKTDZLS4inCGSvyfs1Yk
LL+iAzcBKtY2s72G1Mrd0CuLDyiK8ZLmqbW2MdHVSBpiUc/74r/cr3ZluzhXvc34JSD3qGj43ZoB
Tm8n/H9cuWmRTH3B7pnXvHIWCrAYQ4xcNbNVK+vS8B9K2F12KvwvV8BALvPHdQabWXztTU4lgakw
CIKUsHipJE03ClC2Wlav3fGprXiw0iZWdF/QbFf3Licgkgzi6fAP8zXSbV0C/CkmNGeTmwP/5y/z
pf9BJJaZ+mnBcAJ7+SVpitSsjaXXxdjMvyBe3vjLfLON+s6h3ff3bl06LhjfDMhKEQwuiUQSvQMf
sAqO/P47fEKaS6mcrRv9qiCtOgBDwdv0+CmXsTQ0Q04CZmztv1F844zd4Z1hFhYjCSIR57qy1nPx
Pic/vgBphEN5U9DHMD0508guNT6jF7H98U3QfbkwjQvvS4kDsYNQqxA7gqtv+Yviua3mggMmpvPz
UvZgUanBXDUJTC76MgAm8YAiU6/L3FUWyKWG4njiipZlyM1td5gNh7mxGrB1VvPFJaglpu9uH5Md
FpE4+0vOwA6cXDvBpxAIJD4Goyl29zHT7ywYfHYLEo8GyLLLHLmPbbQHZH2P5OSvXzJfip8NHIN5
jSnY6injEHPprKt200m29mCh0D1nvKZ3CGweV0/k1RTLTRYvR4DaXgVOtqYsWp0hLAZ6BZJNXM7v
Qcw8o0oLpC6FDOSlrjlJ0uuUYz2avVT/gZkcP/9/Ud5vNvOk31s1hGHxN8wvvsvph5UmFrkPT7HP
ByvHrvNzD4MfVZSlCXnFStSu6uRcsW3CXU1n+vUiefZA+tluAieUs7a5oRvdoUIlNDyyeXxTdeVz
tMwZqbjFMHUPc+jey/+/vOfSMeERO+RFaU/v8uyY+Ok+dvBsUE4S4qb5auYGhbS27Z5d3kWIXIzl
Fo62Opmvvrl0yFLSytMIqb1ksyW0rhRU8CKWkD/TfJ2Cqnvj/BJQdsNgH6mZSBDjbiCn0xWr641I
ZbBaPUhMQAPOM3H4lJNV+9sYJcWrV1flDuzU/6m0cfn4e06OAu8bjwKBmlCIScVguy043BbKP+3s
A3zZurNA3uLbX0HvyFcNhLzlIX5L5webSYEKNle0flxd+YvtHh+DPd5CXmltCovTFoK1yr5QV3pQ
A+E4kkOnt2pfwUlx1Qg/FnhRY9DhQ5JJQ/nMgnFyX20QpTv5BSz6k2TvLGmsKyPtuTFtYm5XByj6
L48xPCTaq36GIJOK0F/J8/g1q65b4iER3E5uiDcussyFV8I3f78s0aXDCXG2XGSbdFZ5Q1vczMgR
bsX+YwP6POFpZDKMxQwJpeM9n5qNIQmNiiwoty50Usl0Fwn2az/D+HV2848qyrUg6MK5psqVc29r
u+ddkP/AoiXO1XKQ6vstmRtLC5WjpEu68tfX6r9nWKjVSHSKiZ39IpWWzynlIchIn06C7t19NDFr
L437HoOQVSQGYM4sy/SpgFeGGjtTszHu62njsxMluOz24cc8KIb/jjOpQ0RuSJ6IXBv0j0lXRmy8
NK9rGHESJZGHfeu75eYrnc1yXuziYrKVJGG0atWcKf7NuSCMICPZ3cDu5NWE5P3SKAwWpvgavETa
Hc70I7PiiCssj5mQNgPzczopK0Z7pphUa85VPnPLdwoebqmUFAPBcVYWyCqvcfCgsqNZabv4uNn1
UU10QBoEU8kIcXlP/oyHcyZvMOURR+Pu/8VLpElh4snW+jHkeFEz5Ti8USJ/sPtgNKvN1+6gR0IV
bN8JX56xndhkQt0ih7kWPAglnwCwc5F4JkQsM65MRCgD+BpDBeaFl0jaFAtrVBrOAQsXE9xI3/59
S0zPcGNe3jjYGXUgJex1kPvAh2X7hVmZqozPmMzRscTJZB2brKz+PuaC/U2zV7KAFzfnVFWoTNnn
bROshmLvOZYohGxQ6sHU5mdcUrcRaZGU9Z6Qof+xEE62Ypei8WY/OqmDWlrTqUQOu1ZAEagJWFm0
aHZPIE0rR1b1IXPO6UsgrDYcdb43Yvd1QJqEACKXMJtEI/JVvnDwiRiJLZYytHubwJsuM6f7SPeT
Na/+r0ztGH19EZRW68GB7ePdR/GATkiMxgHkyoDXJ5Tnpw+GF0vDBIgWSmRHU1qJ09x/YfzR+qKC
f3nPNj/USjkB6ohOMNdM2+FKwsnWIl4D7G5tliUhpMZ2885hnf5mIRkdTYIcZ5QrKrwh30BaKW6s
TClMhepPFuE3Ibma/jny4hWXylGNPlNwFq7sshhLWmMHrC240lt50AQoRi7LU2XN+iLeruUqnw0B
nL/8IN2ZLcIi9WJ7dg2eRqteL+pWWu8oODauU6I2yK7NggIutmFerMj9JOM7vUh9O/HuL6LAnXAE
07ic75m/s2SjZ396JgYU+hm+Z935ldGxAkOMjmzBb4aLZUppNokQIxwmZgrPP7PiKiAgR961cF8N
EbuNpJrYj7vwDQCQSn8mDxk5xmuDJdvmd8jyPfbo2hx1GpRb64k4hjjPbUpU7hH78Aaa29DLxgQ3
AUYJrUb1AAH3QlxDze2H6rflQt1gtOyc80UT+PeqnWab0AFfO4byAptDn29dSww1Z28ys/rBPyrw
UsFyh/gPKnQKKjCJlv+BFTP3u+wXBH9YT22XPtZ+kPIVJ94mk3C5cfqY+2ec6TCN02Ij6nX68YyS
vapUCfmfGHTDEsbyMKkleYJ/m6K3C1oXisU6g3FeH8+Orp6h8a4ouDh6t42ywzaYBzfALwyKHi2h
tFwBcwFc2ny9Q/JzSTc1LINyfA7PPcgYvYcxcpJr0Xnm857upPj5pl7D9ZCMup73AHQdAKheq9Q8
kFj0yFU9pOlHrJyGNmmiWjNcXbItgox8UsAMI21rxgraKxvpsp64h8ArK0VuDifMCKB3jzcfhKbK
u5vZCI9Bieb4BYujK4bFGcyO7XDdnuWaYK1MHWaxJmDfieAaI74QeCsUodVsvZqBaS5Jin7mYLL5
3nAVtjKAdMMmqdsEwIcJLJxoYoTCF3iZva5nlsjGHmUPWajYdduTIB2f8Sq+aJlMJxW8PAIWBvsA
rGaAV4gACqYteNe0CmEbuLstKdBHumb9sEsRkcJZUXugHlHZpTpj47FPQuPoe1I+fz65EiRwpm+8
YT78Y/V8nnOzkKtpfmQfIDj+pX0yDucCgPeRwcpRC7HAq8+1+3PA9p7HAnTbTjVN7n4aO3Xn/oE0
FaMHlPdallX7Ya1k94hlrXPEAYkS4ZpSk+xs1JmXp6IFLx2eEHTjdJw/Wn8yGQovxMot1nYH78z9
zgKE2peULsTV1fcv2Ia5pMXIsUkKoQhoxQ/2CBP+Cwpr2fjeKqGqoLoaBBvvnTuC0WR2NTSPnSi7
iRz5+QRq0kuSzw3/7vdC5pacyTyGrEf8j8GtrgK0ai7nJgL8aoo2iT2AndiJO7HWqNqbX/Gt2iLo
tTCMQyxZpmEak/a9mungapklM/Z4Ht+vRZFILUG6MOQb1BPDXNFo0BbTNsPv7t0J+HmBw8nX64zA
SWkBlvEzYnUiM4CxYzfTceHezS/5AmWnlCITtTJT0TNwJaXlBIVQWGVW9vJ/+Yo0tYAK4MTj12rH
+XbHPtlJDHQWklw3KrBSGdHlaDcXf6kawS2gdY8M56UTBP1OK2vPHiwL5qpoJa5kkTybp9/5A+EH
V1sCi0yqCHmksm0+aC90msZh4WwtiyUDap1rVk+Dv81hyg332nncMDnlVh+2nlWKC+jRdXJTFQDd
IJYrgkWZTCifh3Dhy1ftx8pgD5oZMhOztN6C4TTDYAmRARIrm4FfQK43QD8bn0/eo/7l0eJVdCRz
fecFeyfE6dRppPJVJkZIMUMS5gnzLPkK9bP7JPheGUNJh6/I/RoQ75xrMwPfsZC/ix2xjsIkC9da
8+Q87M4gqOzwXO2EB2wvzNUqq/KkNCAOrGnD9ToGfN6itpFaMyjMF+dpGlVO2bZVFDrN48q52Ypu
JNGWjsuO0kINJEju5EH/+4+5EGr2XGBpRecF/mLRkAccgwyCcwvimRwmqFHiArmjOk+/lo/FwvC0
vnVbHYz47YZQ6ynjX7DS3wH2obZHWZU6mpVEOIZVDcXbCL+fxA8rKDBa5ylp1I4w7SMpl+yL4MBk
N+GhqpAdag9PFAs1A+hYhJwbe8jwUUgEf6Osm5W/iKfrjf1SuyOz6j63G8cOdmd2zdtYGcYGOV3i
K/1JH8DfIHXA0/U2f9Cfsy7/jSWn0mAgetuOIsk32mZGPIUmglhgVaOMEVfA/5T4deNkTUb/VF/C
xYbqZpVQOCK/k5crG/+i6dtMUGjHT/0u0BcBFWO9Fs6Cv/7SFOdt73L47eE0QY0xG1YeO3wJcz8X
Zu7ixMkegXn2ycOS+3gPd7sKVGBoz2t1T59DPH+/29GwCDT9KyKkTKCwL89Zfb4YVHvS0kEUaxGb
fzQqd8KPF9EETLRPUREWRqKdEzS8I95O8bcy1PKerGcC+NZR4TIyTEOnnH0BvxKqG8ZySOFyW1uU
hAwHZuVOTlWd9taZDobnJOQOHT2JgWg7C8uuXdohVpE+q9Zz36uc1cUhXHPA42yBD/6R4ocxAqiK
45MeJM2OrkUd0yF84SDKfwjt19rbbh9ankCgib13dyakWsEhSoYkFmtWxve92SU7ZVdDAveJoefl
fUI1JIvFjUqfE69F9Gi/d2QbhMAhkT9TcBFildrldwK10EtFdy5g11jb4Ks1IVEOHFxwrto/pNZ+
e1GPlcaAhIxrVHvFdFglStjfLB+kLidInGrKJ5r33gVRzIn5JIjrnfsjgvzp2qtxKC1QFUBVpyC3
3icRY4WXquKUbSKuWxX+L+ueEH6ksp0QX/QcYBZalqq9297vwioiq8Uu+PZRL0v3eZtLVfVwc49O
JC4nEIvyJ3NV/paO5Tz8lmpcBcVe5pTt1a1WCBk9V2LnvXBP5x5wlufha7XV9UCVE1q07iSR2U2T
/yInDnQ1+jz7gx0BeqSXdGEvELix/I8qS2ijy7chjKYSV1GuIX3JS2PXIPv+o8DmQU1NCrlr+nzQ
myuZfuSX9rlJbur/8KAIKWf1LgSsAwjr37oZ+RihL1bxOaZ4Q7Fq/xjpi5UaAfwXkDE0AX1OXcqv
v+9zHAuX/EY4u/8NU85/EC9TV4OSlWzgb+8cmO43lAFjxWChTdYdcH2rOPiSj0aa3TVfx1BywMDi
4WzRfQDKHTXJVvjUeJZCyv0kiCwIiylAEuZ1AdA3JIom6h3aJEt3rynpATb11nLyLcVX0CAg0G9q
oyVtNusCRwR/+K/OXz+gxpJu2S8Z4Ok4n7u0rUDfiLBSEHwzeIu3O7QYDmCso6DI4f8H4fnljxuy
+1DLdV/uU/6PyajeNmmjQ2dGPy+3XOrYuFxUYuQDxB4n4pK3JRa1cTsRuThyPvKPvjD/xg6ErgTl
DZppR3wNscJvTruHHtYKa2wxq0qvPRl5KNHZd3GeC46FB7vfTmg949GlIqReVATyrtQ1a9LmvFAd
hUg5h/xrnuCwzV92NkN615bjqTo4Wyoq/23qGeJBjdorw3osxF+Q42CRQudnNNb9W+Kl17RDfW5/
OV+b5X9EkgyNA+6iIlzU16ntkRcHgKiW/8kPpaj1roA3luVHE36y46zwcX2M4bvVb5xzPoXUgTSJ
myJDx9Khih7lswvO+mH77DJqt+WjKoqWyPbHK6qhdGFdLtThcT9IvAr3tWf5hwdU9yx5VniOqU0M
kw+8kLI97G6g9hv6zvigm6yuPRRQGzBw5+mr92wQUd9dsQ+A+y6IynbHpakD7n9C6klCZkRqw56c
fyhum3IerlUjvG2HyvY8pG1ZZ607HfTHdJSBqsovMcTZQUeUw41etU35q6cqvG0mAheJmHvqzFkE
wLGje7mz+SP4S8pYt0EDQTt9Nex2WuECpPvpSrUvv5LUxih7oTJTYeyz7sEn8WUClvZ6bJurqBJT
P/2udoitM6j3u9966phr5V+fOezLMBfn3B4KCcJRXTu8Qk+EgYWq0dWe9LhBFZ9ePNqgVVIbufBU
UZiscWZmnhCsmqponepyhoIOTRavLPHKRA6O6LvE+92v5DDU4gQGmFq9Ng9B8+jFoFhwhzYsTxA/
AMPb5mRhCxDw2DEpA8XRYC1oPPZkaUKDu5NxcGSZOwXMxxy0BsVOd/CCNI1OGa32GJOGZDpI/YHN
qdKKGAq/1+yPHQtEslCtqMRx4Nun4U0G3VX5sFnZ2sAtSIM4d730buhuLLd82/EFcQJXCyOUi+K0
LdpPCMTvrYXJXI88zV8SVT8QDT42IfY2kg244Y0XJ/uMdq3P/tW6qDGE+wowevpPmvNDkybaQJN1
/rgDAKo7E1WqUNLDRI/wUXJuEiQPZdyludP0a0DCVBrTCgr+l+I71ZawjBAbcAiSWKHoR5unnPEF
O6/NIN8yTWPk7KzpKWoCcDyYHZBReKXfr5Vx52TwedDo4c6j0ADDk8/wefY7TWq0TV7iXFzOuGXN
Ih4yAuyNJdt8GQfIOqPZWyT6Bn2jAsdHRAjZe4z0fVIYtwgwlk41nHNAzla7G/OxXXHWCyO/rUWZ
1AnGlmO8K/zup3paD+C5P1rMirIeaivmKv2CqIYklKNlMLkOs0FyU1MoOiirfLDPLPaWDyPdesfi
WGkYvnFRe8EdsHYvHQ4Ldxrn2dVshJHNY8mUFubyLmoFcclmJ2d7t3B5ReEpZpE/mjABxBFsZEmU
NV2qoP9Gf/kI80V55fdTLVx+00iEKvnp9VR0AqzPvdEeVQABdfWsM+Ktb+b1GSDYj2g0VbeKU93e
5cr/uhUOo0RhdjfbncjCCjLDPA2l5JBO/q97iXDLrtNLXniaZ13jKhfqutJDMqQW+ZrTFln4bxUQ
DXxiLOclMh2K0dIyFqiKvE+6nvslRDGQ39+lddwGeywmL2II1BQWxGogRO3xLCi1hoMOdVmcAfPh
ArerSXTrqexZKJm3qgXzI8u0KlNMc+U6DLFNBUJMZc9HQmUNQyXtrFnU4qmF4N1nVs3goD7ynXGr
3v07/hTTO8SOSnzykfeaDssF/mn08OPoWfHJ9ZR3kdUMdFTaDjAf8bnioYld8E/qMVIqyoDHAp0E
4Exn9yS+WtwUH/5iPE34ROfjgFFLm/g+IyboWNvBsg+92joh0aApUPqICe5Hwm3GdaKwwfM7Zz8e
gZ12zZPMXeBCLVUOntktEbwuckgecxQxs2eNVo5vVX2GzYMG/vty1GTrq42adpj+qNtyJkASYF4s
YShk6tcfKQI2vPDkl70oUIKQaffnWCOBw1mknXwp6w5Ll3qawFpnMbNQIPmqjIMihzTk0lqlyH74
fT2eVmMyTrJI+VhTBT+7peOdyBQmNNhAxddnQK2yFE+LRsPiwgfjcZO4lhC0l0ejS7pmljStkGz4
2yWByxO5ZBr+ACCJOVSNR+Kg6mFRrTekbKHqXASvybOBHH6LCcrh1ToDE2dq8zdhTEdSIiTFGR1Q
Xn/iEtDp06RriCP0vZTLblxKb2dnXi5/Xx28KCTbEN53o4vLvHM+w0kONaQz7C7beLqB4NuBH8EF
u3CQ8qi1HMmFKr4A+l15kmfyfyYEQg3QTypoNQjVQdh5gEO5c5D7Oscw/sonvPb044e+yr9w1m/B
rp+DbV58aV8yAgF998/g6ZWswhQ0tSs5aU83ecghKm8UhqkEk39C2Vx+jalit1YgAMV766dc9OkT
dyyOSZ7JeAtzUA/j61OWMY6PMvcmGdHe7AvGQ24s+I8plMpIBizWS6HYpt2Oz+Y1WZqHXSeitvkG
sWFjiNGKhQPmeI3JcporLX+Vg7CXxi8rdzyp0uVu4CxoAqOOj191ZSLzSNUYbZJllOtHGttueQzd
3HhBNM5vXqjep8q1j0QNrsjlVybCqovyDQLZ6xIRLwjII2cSh/43rViROqWIHJX4XY7IXaxMLj56
g+qivlojquWovZ0TC63GnzS/uRdYTsrTDXuyUxl9mZVnjQTpWt+1+49krk0MU4zUkXx+PM/Eq+OC
nBVRz+YLYPXt3zzVtMROqE53fJgNb0Tkl2qN75Haw2htZmWTZXAzsKCKdzKSB4an1BttJDVBXGBs
G4FJq1/EbRblU2Ps0YNx0pBKX4m91zXWRbCmduaHHXQmQzXTppt9tprL1CXNlUD04D8gzEUU8pnK
wH4ytolgiiwl4G10uTubfcnmk2u5e3j95oS/D6KE/CFbUZt1LCWLsCPF2EkfGZh7QRHFGjJNQ4HP
MbT9YIV1LuKN554RQWmqA7PQIKsEBFAcCSutScV+wW75Eu3TR8QWb14jcwUSVyXipUzbVabCu7ci
x6sjCWoHpu6YI3KDDT19eKT1NVEW7QxhdHWWuoR363LLTMmNpDzl0FylgBqvesQ7ncJNoyRQxhkW
OvLSOSIrzFSbX0mpIzHrbXF/Ebo3yjgic7NbQLTMvYVuGvqlS6i938VN3Mj1qSjdpgJgvR3gySSm
QeewR0NzXx9drFloHGdE/YWAtCe5VgOofOyhPZ8DDyj8sgK6rGvLl/+o8r/PfKFiTgaItLv791MJ
MrgTEd1Pj+SR1fAwgxWjTfylObQ+aMGX6hWjH0fI1CY8WkiHlVVa7p/Bpo30Kk6o8EMBw9I0oP4a
FXRNqTpStzj6py6MSKnv9Hvj1hr9vrGjOQEZm4SSBREBs4Zh6bnm+VKujqapvffyCf9hf15czWlM
xyRJaQnH9jkUNIZXs2LMDkFtTux3/DohdxN24K8jFa5PpPzTjZt0LsVVI1rA/Xc0Bay42mOjvpHT
sIbJpQRHDtK+IbY8waV2ShkDnB36B2d/STct94pJllkl+FtKwqu5g2hVowd6GP5DmDOsLpP6V/9J
U+3fcr695jJLVCBzKvJ2DfpZM2vC1MDWN0aa2loFfDHu04HdM2kBExkOwy1paoUMHD47txXpmxJo
JWxqfHmX814Va+VBByzmgIGCqaP8V8m5pIRVNvtvgNb9P/eEc1hqVvitMfSinzMISo0e7yCTScMF
r4BGvuUMRCsDpEBn6hw4AQx2jUpCqKDUoAIbujKhqm5oUzMF2J1dN7eORrz5RNUR7/ywuoEyIZJ1
6K2xb180JCa922sHFRJNXYfVurTniD+O2OL3XGiq3njZCHkFknfRX4fg+CSsfFreuL8xyzv7Fdf6
x7CGaiNAH7D9gle2rbMGxHlOJj341a0+yKuZGGKLSd7ipKwJmVxTqvUUdywOLLN+hBxyvFGd5yv/
WfQIpmioK6ko+AXRvmNtrJPjF2OUMLVMnIcwbqUVSZrpR3Cpx4rNsu1N1dM13ynpfblZJ6ZY2q6x
yBhtBWsgliy777ZWd7CHOhxT3qZes2cLyamDffzO+TZFapFoL8Y81BwK8GJS0JEidhrOOACNfkOk
i5O0zwk/2pTXGU79gZLP4Dm90oz9v+JUKgEeJ6J5UoZGT57aM1rHpuBXr2y7NNElKCILKiNCPDHN
do//OH76urd0WjIexA4es5BCd02YqG9vpvT8wjbp/a1fB7Xc0LSUwGGz7yXxLyZEbYNJ+DbZjHb5
cOSKrDsDqFW/9ktznX/St9SnHt2HiS9E/wdif+NSK+0ijYaqpr1wMdxfrEORZgHoNQ9xryBjm6wP
+kihx2rcofGkD/Df1anKxeGxXdep5OHcExtzMckMxJBBKl6u8y/KmuoIqHsW+t420khahFrr1mh2
G6BezSzBs9XXJCzcuBUogCW7qBaRYiVhVRd3OPt7eyN7lxoY7Q0VvobH3mEc6W8iKAqDM4uJqvSF
QsVxbVWNurMqy3NY+KLjKFMGwlomWnbKNE5K/ak+9iHv8Rd+Hc56qs6vnGslpNBk3sN960okQBiY
h4dqIMEoHaW4Bv8RwzuOcHXo5/CWxZHZVgwowpPMcUyIapqOVMP0IMK5nfgWG44o0x4ef+83fu07
bsDt4Kd3zo7iqPRMPMuJPMbtyrZFarfUWzhpDVwzm6z/5AEuu4S33apLTTl9h6vqireM6ixQ2Tyn
djqLtqRbSo0V7mybNrS29MrR1b0p88vZgby9+I+1XGW6jZQ6RQtQwyB813qZuxuMT9TRqGSGqv9x
3qzpNHK5s1A2SvQ3ikH0PJPKrgp4g15DbL9ylYNLXhoPd77DKZ22oLEC1zghQk3RTLQ/0BFf1IkN
e+DRtjqrifVNXFA32f4MLc2chkg7fMSd8/V0TUNQJ/OVaQ4mpEl3/KY7NYWS2YmJMvY+tUWyo+Vh
RJohAf+ZPfzQLYlwIDuzYrq0wvd3GjVCOEN2yAyjfDHzXmwPtHP4g9ljjRLcPYwUzmLgzvqMLD2t
OmP2mDFxNzFvUCxtE+Iq4N1M9QujAWeMM1Jtgg9DWyWd9n7HiRZd1RIKYHc0bo+7Y3IRhcOPPOE0
EB+rssls4F9PjVqNMrt47Da1XC+jDg0nztnw7mlnVJ7KNXOJup3Qj0AV68Qz7rqx5pW+7pxzbqHk
aXRaojx4it76a0dl8zZIQjU8WHDO5dMmbmtoYGXeYecRQ0dC+l+9QiEls11e57h3gsJkGqlZl7wI
f0RFk+rbCQbp/wEZDcAfKMwRn+8MLTnSwreAnJdR8LL5E7ZZYUzl87ieNpXDPTSXfNU+hVSlAdhd
wN+nIXosN6BGcxObUDfgRhr5WsWx/EnD8uX77rtoZxaUy2wYlsvGMVJgpa6VZJMVirnhwUChD8+L
EmpYrDbaBCBFPCNmBR89S9eFmI6BbBYFUdwGKUYxpL6XVpVuqsVfA59P8ZCXaUsisMaWMumal5mv
dpyqFd3xclLya3N7ggJTh9dsbLEHYRyy6eI5b5QccLjXkqa36ZL0LNSp3dM+p0/p3J8YGeNzej/z
10VYSWPZHiINsUFN9kbIoR3Wuj5OItyIxUadeddIA632rqer6dJrqKdgKddcMQchVeY/cp9QZ6kG
frs/esHYYranCeNxgmqtMQ61fnhvcYuH7AGM0HNGzNVdG9p2N3n7+r9mcYHj2KGOb45UwKD25y08
O6xUe9HQXQ3HVVNHII1pq9Bs0DiRQT69ZoHqpo04Ee6rMob6jd2PW3EoYKLEwaA+NFxxURjTyh9u
6wZd7UvTaYQmySbYMu5/Ag8aazL5iOUX7a0tE+a97aC35b3PeqgyV8CsHwCLcCso10iSNqgLSTBl
8TO6vRVqV/5av09/TTAN0ZrP5s8TkFsazR4SvXklA65sIgsAMKQcFzHqo59o861HvW5ElPfBGVEr
cr/TCtC8p4tnYxgKR3/ovGT5O1UKl/AR78ink5zXazlu6Z4MXA0F4IJ8j4MsPkGaP77rqQymKywt
jUkym36CV7s/M506FocQzd9vpe28i/ME0fouTkTjNoUmx2oFtKbezaljqUIaGYvMwM+ISpDaize/
5Mk8qwLgqeZeRMgbi0eXPgXxs9okow9KDPwgqsMml8giKM+oMUoEBRoWlsPyYfflkAvdpJcdhHVw
sriB62KQscbgRJbj9gAtRDhrURRhPDGOZmQWW72khdTIb0Bk6+QQCeemo7wVUekB5cpkIo2VYWf6
Sf+bTz7A6fzihFrj92x8q3Ipjeu4Tje+1P7xXQwY/MvGOQdmCndxKYYxc8gzFbeUVQSCB15/eRBO
xz72nK3ykJ/79tCwHdrYN26JZgrukcLJ9P0hD2zvkwLRjatzwCXVzpHkM9hObs3MPEEAz+78xWkB
VdaxZiSej3sdEsTBvJ68xS0yF1YtGjjnjaUTzQeRMR1XfnKGzO2g7B/vfV+MxDtqg8cSg2aieNmP
FIunaoCUtNJtGV9d+r186Y8ceqJnZvEZ6KU9uHyqgNdahAHsrnuZS3lMH5ewRj7+IgU8JW2DrV0Y
weOdU4MVFDr7SgoLVHRderN+EC/fD9P43uM77luE+fzMzXJ4fHW9b6qhv3GxQrx6l8IWjUTGL8Tr
+caaxRvtJkY7vAfjKv4oMWqwULRg4JX9zuMPuOCeG/S1OfMz8hjR6Lb9mL19wb5PnRz3BCV+t6IN
+CkJ0t1LDudGoeLWJVsnFMwNSBwp52exYJ1basx8O8orZr6HzC8OEnIPXXLQSLm8oosndXjQpE5W
vGMmZs/NNyYxXNtDDtF3RgN6A/99MkR3C1s51HVRu+9e/ewqvld/Y2TKuUPaAKEmDq5nv+3Ige/R
y+gVw/yAawnmSvvHCIETRvXCjlxINvUdwKDM5X6tlLqRY4hNqHT6JzwKFrO8eu19OOYZ+M2gsCxK
pVGvmJcuuAzVsqS6DWuyf4W2JtFTp4m44r1IK36I7BXzsX7FiJpIrLUDBqU9mA5OQapcgODOVgXv
dhEcgDUjD2ppDX28s9mrZ8iT57CnFkNvqSKSxz8p2KIHJ+SzypVCPLfESTllUZFfY4ftpEdkSaAm
kZEOdgUHQVrWPdf0aVGwCQBcWvrN/UgVJRq/vCTNTJuB8fECUrIHUMondSL/Y2b80uuVPKFXO2jd
HtRXOCaHqg7SQhXYvmE6OwqtAPzIbj/10IC0YTpkEMzfkDxE3YbnGxmRXGNAkX8uB4HlwHZ+a4Vf
ZIa2M7JxlvdOwCo1TvfMD2hrOrPS3+uug2pOW7EdDCOAvGdw5Oo48DLfeZpd9E8pzfTXZ0yDtge6
qSlGDE2SeS1GqFmAB+ff+i4OrRnaiHeyiGax07EidTiIPnvxv7dqirf+y33e9PZYq2XkFlG2u2K3
berPF6/0eMhSDro+nCxkEo9hTUdXSUKQTK9fXmRO1izCKIuZuefgZ7R+GVFXdBwvN2oL0WzTSnwD
z5eUZEubMxw/VeJLeoWrpmvbeuKP46Nz/e4FYJ24IWwy/OZBfW+6/KpKnv1fF6d8NWZVV14vxzi/
bFPSndgkD5uZD6H3kEvEnS0na9dOicuJusXGQhHSpy+1H07S9lLeoWb07kc2c7wTBihZEG+Pf0WD
MdORyoaAmbbsVz6jFX9hDBcVT6Ae+YRbhQoVw7k10xdnCpghGh0eDR7wU50dt7UDXWgmotXaTvRb
lVQLrxoErUVh3IkohRRgUAlaMiZmmz4S++iYQ83lniTDs/L1uRhcBPNlK4XtA7Ushcdj7fpcLBoJ
0Nz2Wd5Lj2IuRJOMHLXLksnLkC06e1WVSzYsAf6E5v1AuB4RXlwdvvoyFBIspKYfKVIjGO0wy30t
/ebldKc38u3xsv0yl24XrUJarnHNtAW3PJvoWIjvqB67WWvXIecpMxybbx7qDV6y3IQUj8vEWGEC
A06Mqf7wUvIK2ZikYNqv1yw73HU42izfA6/iE4aXfaKPd4gKM2FuaRDbRDB8OIem+Km90A4/5owS
i2ygGGSUjuPXEdjzQAxqpGzpKXVcXTnDwm3ughmEHzARy7vysJfVHefw3vQuyEqXFOMlaak4gF/p
OU+6/64X8THr3xUyj0VpGZMreNWO8NOC3Rj6jB8xbQQi4DgUgACIKuV0Stq9hLY9XxINujdhmU6S
24EqQvMP0hL72SHromU0tK0jceJ8ET6ZN+MnTdOQsYnIZRl4SAZrVxGGyHzAbcVZ3f0l6VtuWWfP
ynpiYDv7gbhjSB3c3rSW2xI4kTqknqF52zrkgZOjWAx7Ro9xHK2Xm4dLl6UfpeQFdL/abaZDzjEI
poONAyTuwkCic8s8MWNmzKT5QIEzFz2b0dms1gFEJWABes/yI4utUkWThWThfO4qP3ku0WwvKF8w
hWfx8MW+ueuGCtIXV8YOtPvTO9gFi+9EikmXc6gBWgQwyhBgZihZD5jRr46ekg8Pcf1gi/kdDWdD
11etAh1n0Se0lBlPfQryhW6wL5shEvnkdyY1q2DaCWsR1CPOYdtxHZnT3v60J3eFDC21GP31isY8
0xeP0EzMK/+3L8/BZkHef9GwhPOZK7JbsX8Z5vJa4by1Mcu+NCzMEtA7zXmTpOlkUGHfKPzUvrm7
1Oc6bnAcNeSWJQCJyneprwnaaZriW0fLNp+BqSfC8IMWlKEg9LpT7zLmlekLEzW9h0z3GeE7oK31
CRqTkIx9Q/kSXaxZ7iTv7ksrdO7TQ+uASCuPzjU/fG2XukiPCDGLDeq5cPJrdEJwrv4vIbp9iIB+
Xxrmj83Amcc8slaLNHpAQIJcI/jmJbOG8RRDGqJjZw2jcbi9amFA0aUDlz7slOjCVqSZnE+63u8G
oIIJfI8eS1orpYfOh0oxXnlDO32jrGPU5c0cqAsdUKAR+bN03jDWl0gXsIvNWXv2pnIWF5gMtNZF
5l8s8DLd6fz//JoaUEmAuGXa3ISDvGoKanPvGxhOun9t1DINQ3OOi6MWM7B9W1PLTTreK0vu99vU
Su21Gigpe7ecaXCOQR4j1bQWq0tA72hdEJpZVszzKT+7Kg8BZLakCMlvzHLw3qm85GmjDYhMPXDr
/AtEtA6XwZDDLCNRkVwQpv9abSEsigS4it31OxyxyXAXOb6ldJyODeWJm5Hpe8C4WkcxlvqCmrjw
U60bsBEjAaN3GxGdtdAenXWtb8L/Dgj0IfqWk1ya7YejbhDk2XY6ZDD3P3KqVqIK9d1RSnkoKrHl
XFqQC8737lT22cCgGITRZ1d6f9h8LxYbOaa1ppXoX7muUVAmZsTJKKB8j+DtK19jgynmAkSq6r1J
Bk14Jei647VxxQsZryL2n4eHmE8GypwAevGyXTq091E5n1w0dR5xNM7nHLk5JbbdIwlp/8CkZN7X
u0YxoXTtd1N1XjIkAoCRpD1iU7aJus5W9YffL6U4JNE7gp9Kvo6OCcdcwjHMm5bSbHjJfNjUQTFW
E/3h+n8v0kvA+7lbuY/Rm0JxFWEIthe4dC6lkDO2lVcUPDxKnhvFdLGxU3+8ZrlX5YpYDt4Lzw/Y
WxJHJdqrGTg9LAp4cmrRWcyRCwnZ+1cGzMF5B12eCqj6d5k6JA3gnNERozYXXmaUA96nIYYCLKpn
RmPkte0xkQkNr/bZT9IH0iwBcYOa6iF3mZtojBaUfwvrqZh+4CmivpN1URBkgyFsKDDu0XC5smki
FLQhuPDY1EKTpEEhNvRGKgRSViUwpfEk3j+0OSVVjc3Ap7tiruf/aX2bpnLQp1KwFjLc/rv8zLr3
5J/qWSfDMIGMQr+Y3XUrtc+8/4FM7JYZx67nn42HdQmM4mMQeoHDSWYoTbLCPw5gSebT+t38eq/S
WRjrlTiHg42Gk0QuyWG9pgIq/GAhgYa6nUixTHVuxxZOxavsc4wi6eDtnL/5y0mOQM+F7txvIdWI
SBJa/zWukhyHVQZsczYHmzmM2QCEW+gozKlIx/RKf7SGCjFA+QUcwxVhInpS6xgf7k2e1Dm6QLtB
eOCCykZTjE1646lKtbPPUWVe4PUW9RtMqzsVtCd+4wzwNAyANidkTJoUtJFMe63JIoV4GqZjAou0
SuWfxPNyGdbpQqeQZIF8r6yX4G0Vnxk1rsTvxryXfnsjLO5Wo6F075XJlSEDBSlmDjbe1aYQFGmP
fYByRGpEBxuCHDejtbYhXJNbZHeMWuUdseYSE/kLi8psOyUVWJBNa2G4Zk2oDuYNTgY7Rr/CztHH
WjRmM6PLcqcnqnds2oENonJdwc7IfO4I75sjYy+HV3O55reDCBuiCK0Y85uVEIckU11iaGpX5YhX
S39Q+GUcV+bWr9XHk9qnIQ7I551ZuzJHR/33OsNabMuXT2J/HM2oAFCI7S8Ptorgq/44Fo0ZD232
5ZzkV4DXSkyj+hV+p1jvY1ptrDCquw4qE3WaW88aGq8S85+lXQkUAcRmHovaT2zXR9GmA956UDo0
kmEVHeA2+dvgBK+r11Rtmo6UBPWGpcgMybo2XUTeIVJluxQiHbCSIobYBJQVLlTp6V2J9VI14/Zs
ASffzyMy6m7EUAdsSprH6Lh/NDrlXMTIDz3bhNOlrPI3TJkCGE6IIgIWezY95I36GCS5dyruES/X
Zj3dC20ZwTGWWR+MID9WVrvjRb6RnJApoP3QkacASoDfkhH4yEKcA+ZzzvACCT5093OEu+UQ4Lf8
wLv4u+C9ul6Xj/rx6XmFRnlYakJVrMkCw9nslZ35/7VvDwpNaXtLb/BXVP7i8Q9mZBLxhWnrYNTv
YkH+VdCIyiLsT8r3G0QkQ1ALthTSd7FVC4k2DJknIxcqBEg3CGLBI4XFiKe+FE7WizcwUlADh4PL
BcKkA72Jk3FsIaipWnZdwHjcTVIDzCsswnZyumbY0/hJPiHxSFaDK7cSdfRess9fJwZlZlN9ijWw
SiPhMeVsEelvyK88C1SXpwbEP3gFCITF2pBUvoy4dcWqOkIZKLAYldZRRa9cUGNzNtMoAynpfNUw
s1bo77BUPqOYAhSQK0gzfPcB9BlQaZ5wwALmtlMn3wzFqtK8lfoCADmk4NpMaqCNIiM5p9Hgr6Bn
/2LiBlvcA6nN4DUChvlFwVCj+xfMYbD5e60Y/L56scN7wVH/Enl+VmvANjx6WwYUXPzWi5MD8NaV
jEkdxn8Ri2ScVAnlpPmbgqptiueZijIBTnD8aRJ38ZSmQlO8GTprzAgM6rmCnD7fEif3vOpmi/R+
anGXiMh08u6llUc9i/b8Fkm/PxQgWTmcED4CGOFOHiQhWWBbdup7hNaVXkPBOY3Yeq442RocDiYe
Y77KxsGbrIJJbduxCFFbK7FxIPIdebsPlzcTdm71arJ7HtdR7L8jNHNubJSpbHiB1ewSCUSNm2AG
FXRTaBUADZBbLMRxdt2x5TZKvYRamrQsg4FpgqBZYqG0jOBetPatt78zvnmZNFklJU0MoBJdkkK1
9oYKcNNALdfbhMP+rBmxWh/4bXdWOZmOup69GLpxyixkvW6sLHfz3QI0VVs/SknM9aPZV6I5hlUL
8ukDibElvFq4v/Lsd1/wlfhj+TOHfTdyLwOb/EGWUcUDP7hQ7eDls3mLaiEv92pcBpe2bshRHXTK
FCEIC+Z+Y3QK8hhU1pCgc7qAuAvBQ6s0MVP9txaCglElsJCERw1bDkA8tCAPIJT5USgIWas6+j9C
o0rimNMMuAKhisaxoIWnpguJtGjXk7ZSgCo5MiVnTWEaUb7q8ALUC1RuM3gGt/TNY3K0uBnq/LR8
pVoUk218JXX6xDtZFfzWtmWmzBqvUIVt7QkParKU4fsUCcetTye9RuOedWHGBXf/gZmxCGz7Px87
9ojwjkgrZA6BqQae7VmDyw6ZTnSmHH8tIyR+v7z989IOuldpHkcRb7gHh09FpHHt8CEhGjHqbhbC
ddL3o/vGZakKnuTbsVShVe/ysqKG7GrPXHfhbqJhW5zgT0imDKnwbWwXJQAvyUeTkFLLdqTHHe8J
5sOu/A1CAU0GBh9UU4gadVqanZIUtpnTWJ1Bm+90z5vWdXuJHVOv2AZqSO96a+Nlv7//BKsarxIk
u9AetbRmWwTG7MqeB8Ngbh8kYZTR33eIg9/uq6AI+I2NHPZqsV+KmbiRN3g4VCDAVoUbtp+JZutE
YVhZ8TvsDtfPUNgf8n8XIzgX/6mvbp3XEhgYogn5gFNa0sLfl+BMna7xQfldiYCDA6gTwJi1DU5p
lhsZibxKhCqH7x1SZ89uE2BwrozCLcm9ytTS/+ULGsfy0qb5OLzHCs/WPWYB4qSOWYOuanT48Hdr
001ST5hre8GvzLExa/yhLckAPMSMulRF/Y+5xqL83ANGJneT7x/CTKQf1omK7H8DVpIRl29kT22S
vXyW3+5moQZJCt48HdLj5mGPJOwRRdqc389+U7TO8nv11mK7LpqXqsy9gb7AKfBLW1NqoqpuPw3j
2XqjUDwfrkVXsRj/EncI24mFa6+XBjwEejMG7im5PU78a0MptTMRya3zgTxzZBdDcQmfa+q78tdp
YH8LmO/BBaqx+Mk5K8hEIODkUdQeBN+r48qZ/hZmEjsqPfosgBqqWVQhT0Y5ElEhsdtcbi4CFXxP
LYtGahM2F6VGWoVQvAwfCJTTL1OqgeQYVLMsf6qSzcZE/Z62EQqR0JGLWHh7REF/OySqzcWNnQs3
rkZnQVBGRzQ+OIHnepR7Rn85lR/BsYGTSTAMXwmBbQym1jnPvnnlKLijPCMWuBlzs9D4VkLUbpgM
HXWGfdVyEFd6FNC5or8OKUV3PGVkmW+IP36JHVZkqY9Dj9ZgvYQcFgShkiP/awJtQ/bTUEXmHbOZ
I7uA3sywiWhllFE+9Iq1E36Ao7urlPpHW3es17PpTePtNa5m0OpXyiyaycby7w7FB1xgq6hvJSjB
hPrwTDUZ5SLwfu11RlQZV6IQWAlPHBci3PmZrHNEK0vpWGsR4zGKOElNiw0ihrXV3fUmbOXfGJ4g
OTrNX36wmVScUgMDp8sHURFYjRwNsaaSeGdzRzeMS1imyo6vec4UHr/I5Qh5MqqwJih6FmZwab/S
hPMs0ERTeqOJrmjyA4tJWKX85V47Ro+gG8WOhcgg/WH6rCuRC2yFg+NHH5I9UrgE0OieMgeQMDi6
u1FTXNzm1hMrCWMZ2YIDJE19i/zQqJXeKMtxsao9VYn+P0xEDBgynkftsjYky/LEV3CQJIOciZ4D
H7pQyCqOJgZ8VKv5KEdEZ1Nn4jTvqsb5cpLAR/mjAX9dC79/jSjA3RSaJtyoFQ03wpWrTTDJaEd0
FfVJLtRXBDumJBm8ro3Dsfho8ydMWszCV+Tw5TJGHJPHxEfHiUMdwOlXGXqaKFGWM9tgiyAlp8lg
oTqdlSsS+9+0lHfuTa6SdpQ2JeUQdjj+V1paqlWJyjm81NpXkvE/a2nZ4kaK7u/u3vCNjMz1TqeM
bHnXrBekzqUgPl25uIZpuhoYNWSy9+aESm29PJnzvyXS2y4lwYTlKRT9haQI5butgu0J/ERj9qd8
rh/SEIJR08DtA5VpcF7EsX6TjIm/DQTmtUUSqx3Gk76Otnw4SY47fyhUQu6rj8rIfdrZRuDehtxV
hjseTlx6/s+RgmdtYVz2Kg2i6NrwEQ6Mdvs7tyf3D0GAG8o3KjVucg5bFmMPZN3VqzUU4Kl2na4I
C73FRs1qqiJt81lxxymwYAIZypArJ0svuMzMKNXj6fvRTHbKx+2nZK/bq15/ewXmNiMehEoj8Wlb
92TBMK2f1oe287Ud6hdoYD1+yQzNlXGWM3ECW+chEPPUxfRE0eNhYo/rVZAF2yrKmETYCkCM7LWH
nrZS4LFFjuNfJcoku/pYp5dUY6wJ35OaVEd23I3l68tvr6gg/bq368QAVqVbuP3/4szgNgagiB/S
oUM77lXEE0ecuDKGnyTmpjhao7deuX4w1+xsgp2azIf2wnHKxOOLYNgv3WE/Z9JYkw6zh4tQzkn/
YSWY9R8m/env8GY+vE8hPYgNKdcnD2FSzipp5axa1ANR4gnMLBOBoHb8JfTCiwzyytL9w+WwABvt
F4FGcn7E1NpOtd1ESOUbEo6/VGL8Tc7WL5KM2idzu5yCwgV/yLJ8jo1tbhUtIEIzL1Htkj60W/O9
TF7RJIbnJtNEwYz9FnSIai3I/zJ4gggFFy4Y3DMnS3PBDI8lnaGWTO1AW4NkAOHYRV1WmGH9rzxm
ScZMtJPntNDpzIJtPlwQiLdAzw5Y63cXJa7K+fTMQ72c6AsI5+/y7GkPfSTDn8PUTFbq34ns6wwU
Tdn1UySFbh2k0M+ey+jkDnVe/fm+bLyR/3Vom7qBR7aglYOs33uTeSfQpTe1gucH8cRuX+q/QwJz
iqlrnbOx0gG5phXavDV61vaZ81+MjojS5FY9EqJKRAkx/DN6GtSuGvrQ+quOGGEuUJeWW1JHlrue
cn4gVBXZTL+7vhRR/FUy9o4EjD187WokXduxUdn0wpV669Ejmqye4W5+5gE8g0dAY/y1XZDjfjJR
XWHOGw7ju1Mr159/5XmBK7/P+f7bkb9EHBuYzsAXUJ3kqln2+RyrqqCz2nohDEnxBxAe9PWRcU2g
lEPZkVQXFqnufBzbuV4x++22OzaXiVEpkW3W896l9U+061dYBXXHNmnOqjWj6GiJXxvYWiXH8YBP
/JlTovXHLtpfWh3iFR5symdofz4Z2mmLCtIcZb1VnLsHRJhfQB7Ybb7zRY+4zUWeGH1Eq29+aLXG
uZFTjNuJs9G1D1orilKfoRCx/roNLSXC0YyTFtUbnFVZ/dZxZczWZBkdzaPKwU5t/gn2X/eSCGG4
mo4aZRBXPc3q9OMxaqhVyRnxSogHFKvUCPAtM670ykB9ul7B6B/VeRFsVzPTg2LIABrTm+BSabKX
xuk2jKY0yB/DjQELyqYgE7iFT/t8L3cCS17IzMwOfJ6C6AG5zeGcGHsKTC1rqfDcSbmZwYPSsMUG
X3kjIF9sGcZWY/MBF6m5vzGtAFgCT5qOy9KpkxSWV0mW7yj2uP4PAUk3N1bcqdKEGVWNQoWV86cC
y8DzR4rudufL6ALw2XZKQ8luZsARA+CAXQO+yZdKxW8lM8tXcEjYz9lBDKvH4v200AM+IipL/6f5
DJIjVnWdLDvzGi0iYt7QiUi8sXH2P7aEdm8ujX6FdRqIcYcpsZSImGAUu1FzAn6k/sbo9J+FnZsB
mtLWXkxVGB2wkm7XALGu5cjtX+B4Fc+mY9OWm9FRCTKWaWvaa51TUQLLvdeHMQNno50+VmTR41NP
Fv3/i3gdaew5dPy/7hGhM2V0FA15vV0aSpx0JNP/E6mhg6/w9pdfHAS3saMhCiLkBUc7DSFURolK
v5JpqU7ctfJWU1imp8KI7x19btIBTw1XOnBuFsH/nuA37X2t+8VyDXvwj4Ss/kX1kga/UQPrZU12
iY3FAVhlpsEzMf0CVUFSz70hH6EykQ5cW9WTha+XS10CW2v+T2kniHl3L50v8L4XoyTvdl5st2sR
jmMdvZ25SC8aWZxKqVlri1xTbi7V3WtQ5yN4+8m90oT0uC3t9rw8e4F/UpmdGYZ3Wfv6c4jN3qag
+CziRg+PwKF4/oXnFJnH9O5psi6yTMltsVpH2i434aSQ2NMUwCsIgeSnoPMfEP284gIujUKSX6ho
iC/bRYKYfXyyaEDkN7RN+tsE7sY/aa24H39ArHNi6bvphpYUhZL6Smpds1eNbJbDXKXmA3xFv2FP
NQV5FhYHzPGNSwzhqTMLo2gpHxlhAZ2khOwssumop/kIrcIwjV1jAcuRxw0qW8dTgPuaRGcsrC8g
kWFPKQH4hzH6eGmAsPyLez6XM2SDEvHMQZ2v9c2RXRxN9BES54G6YoC4CAjXO/oK9X7sJ2eNfxx/
m3lCVtidJSl19XcBozEAMWzz3wXGJ+b0IvpzAAZ8swTxU+i3kmQhJdOyIg7+22TUKXOVOg32QJ8b
32hnKV61f2XsEqKn6Yq7JaIBQ5dJxbE3iLCgBujoYNH2uQUfmOxzAR4GjEj/K39ycCCp+5f6jwKR
q1Hi9CxlrnbRR7QUBrej4eHkSqTuWDA8aftprUg/1d1O01hGBuNo6brGUi225cV6Vyr2tEu7MMaK
2Al8sqF2zMgF8tmo/x5HMX5IRYdJMBYxlOwCrQTCeu+sHxn5jsmB/bEI+8DL6xNKdtGW+oWbULl2
qDHc33wqXQyG4GPxtCowZZAWmK88AplgPAG9vcJXT6HI1YbTV8wGG4NxEB2h7AlWE9ZsPmZcDbMK
mR8pdrifDsoHmldDcgnIiC3+wht2T2rSwm1I5/+67T1hKrKa3iJ2MyetKl+HiT5pOhEhdQ8zaPcg
7dXysim9TQhDo4lWACxxri85f6IcQZgRGG/OQeMkHF/eCCH2sk3w1FHDgTy+wJ8sYaqQiAPiBw5K
pATQpD3j0HvWAieY/yI59AFMQ+gdizzqzLjIEYTNDa8kCntMfSaUwvmaG3Om+X5NsRrvednPpTDV
bjAqQRYWkCOWhAHAVJ7Yk99whdS5fyRjWeStJv6OVbyeMWcs+p3kgrO2R3wMV37u4xFi6bKjT4iG
6z/rm5c6iS7ZkfOYIRqBLV9VWrj23bYPgKuKC8hof9WPRe80h/4DEupYVPLWCjwTSt21iLVeUkCJ
yvtOBNa/rG9SuqBgKSLZV52YPCMuHWAsHgtfSvyFtoHFE3VxSyaRoXYstBR36kT3A054Dj2QSDrR
r5y0wlVkkeXjF+lo3p65owS2832R9cvDRvsXuXZjCz8c08EuZE2abiFVQdE6tcsEhA7yG+oMhp5i
ZIakE3dYDhSohjdPxCLxnOLl+vOUpadSMf+VU2hIm02O+Ko+K2MDd5PlkSOOJK0kyYo60RvSlVUp
ulB5Jm9wOVIxxQtNiptGV8/KAx/bpAl7x59XZAjeptMzGlMqOBkhuIZYaoImhVxV1gBglBTxprrs
o4fe34KS8YsyYZDZ1wwywHe0BryiSBwE4vPunrR3FzKM8K0HidYCcUBZnfsi4jBMidZeFxWAGxYT
NK/Uz6z75Vsaaab9qMuw8fr3UIpxrHClrQzYXmRZeRMsE0+YXNZ1N7CeAnfcQPhKddkBrH9tuCxj
2GAMBGufCtc9Td1joyaQ1luOlK9xE2+rpBgukfrg309sz+11u24vo4PlNWp0BF3VwWbtKRgXHvKz
oQCQGNSmxmGgKnPU+bflfNU7HqdZdkJgeOWu9ZamGXgHfBT786l88q8K09sIt6/Eew6lEVjZzwlo
Z2zcLMS+p9XrgqZpmMyD6PqhRmPdI2y//OKcP90lN+w1VAFijACc9EHr175FnDu5zzlQYE+59Hpc
M9pZezxA5obG5uVBoTZUWZRLz0Jcv0RjUkBiC40uB9FHgJDzokrh0Q/WAH6+hEgffCTGlZuzu1mZ
m2weRUjBIzGmbMw9dyovZIm+SyUSvrMBh+AxJd9E+jv+hzCTyPhcWtpJS5S9cmJxdAPfuCnlLj9c
d90jf9g55tr3h3vY8eE9kZ7wkLGM+6ynJZuohpbRQInaKtxC7bw1/eGJyEU5nldzv2bAPpE3uV+y
HroqT4NX498IgTO+1EFYmxLBdQnmUlID8mKvYsmI+ld4kUxfZYJUqpSL020EGx0lzZRb+b1g0/l7
mJfqzanJPLfaVhEzon3/Jc7rlhO54l0LMhN3L/YqgHTwRrrzLu/13pf6H8mmyqTtWf1ECHZfLUcZ
p/BO3OvJRlZujB22XpmlPVdLaXGpPi3l3nQpWI3LjkyOa0lhj5oztwVQcuuXwuegAnL++JDSxF9R
3+Q8UbD/KUcYVu1vwJ/5WwMQf+aQm+bFrC9x6thxq4alCh/jTNXr2PpgAMv4UyuR6xtEShACS66m
bD4JimO42rYa48ENsARcmeBDDouFbvj0Vo/6yoRye5CHHWoy+jwK6WVWgld9zzYMtRYoDl8VPYm0
y2xe/18hMB8zhjIkS4B+tkx/2gWq+7kLDzHdQApEuaSu0f9nvNRG1lj+OuapI+4bdhD+XIdhxauO
GRhudI9jU+6r1sVyG1Dv2eBIMM1ESAnS72njEVf9tudMIhONZUZ4Q0YBJNDkaYplWB3WAqF/oJSx
ahSyHb4V0Ieqi/I8gx77q0g0J8TEJFvPsZpEawvFVd37MnQpUiCLR01Z4pYg2KWXWHMoOad0fctw
GAQi9veo7MfUzzRvgdqlOM6DlWXc+jHcea+O15rDSZRTvJ3DSNXkA5ih98WaEl3In8E/gQaUFUUr
12wbDhjGRTdkb2yiozHmOAO4iFJtxIZSNrArB8M+tcR1oPFyXJ7XfUglDEOdjejrWi+Z+7PeTTIP
CwUYK2jUkoIUm6ZRJvmz/pUhKjOs/FC3/cJmqq62oV9uPKviZwM+ixqQwrGCLsFeG9wH5bgWDsZh
3brjhhycAKczNcltnRhR8+MynTysz+FejRpCcB0Ah73I0UD8wItWBo/XlonhHoN2E8ITJYRZySVQ
XIqlAfJ1MGNgJ7taaJAU/U1M15vC2EFuj2d5FTKNWKVeVISiVoC6CS6LyzJlrluPE+4UbOFVX/kC
cAu9ytW7CGTA4vLSCxJgTw7zmB/LY3fz/QbYKa4Cac0vIpDgbW8XA3Y8u0XRB+B0xjxaDHz7GyoD
yf96KGUSOAXBPjqa5oHVz41EHPXHjmo7jqtQypvGMgLHecn/i4Xop7kvAlxC05317c++lBVdKniQ
cz92d6hdEd2aDtM2joSpSvIdDYkB5F4nw+KDRTMXYnXT/5WgWn5cI+hvt670NIL07sVlt1tEejNk
Tb6tCscwTmO3EXTR/qmFoVyYVa4zyIQ3rbG4pAjGa6xO+gJRFuiCG6uT8LbTJ5buVhYty1pgX7TA
xl+mPiyJHPW9ZND//EJOQtElzh6qn/HCTRLu5X7rshlUwX//PfjnLkzVFX996kL64BPGEHglmriF
Q0+QneqXiken5QTawddZnS3oTq6RHzJ395gOZnbIRZ2PjG+wu9vRW34Z6nvluaYEsqlXi5/4tC/r
zS1MQpyGi85zKJSf7Hd4sS1Fjq4ttuuwZIWlLQSiQg0zoI6hV0peUmnmCHHY6onaE8YUF2u149mw
cO9jnHGGBsZ7HPTEOmX1dqi8UR7v6pnYZZRbiVmwzRXPF5itdGOUsSLFDUtYllKp7emi0bsJsiiv
M1roU1+8RbCr2p1/RHmNmQrVKPW15pVAJ5vHMa/SsBHEJjqPEZOZ0cyhfq5z/KfArYIY47Zt4cVW
I+h4Jlgp8LlOUmLzftY53RBvZdtxZ1mjcSIA7QFLxmJnJP9Vwx1+LMHD+XlaCm/g9q1yOB3kQKxH
JMVu6X64n5cr6UfIKy74vZq/rsJSkvAzdreDBJMQnzLy7pt50vUOpJ2N2RTr+FKUT4qvdsi8vq/C
4V8+3mZCv/VZhdAqOdOGCyLC2VAtCyE6epOUNxaNicTUJS9uO17+xRs9+Jj1qZbE9YY2MpdtscoU
zP3lSPKPO9f6U3PC2alDZJvdCGe1RnjYbJ6NOC3DpeWY2aEuUOWBisTPEaglYGhRd+pIYSiTMe4A
DKE2sDG/AzgW/Bm86qYE1nFflGCwR+va9AqIOZmYC2CR3+KaMh1QrZSezpYPsDW+dVAIUXqSTdyl
LQry1T44/kX8vPZh56qITsH6ze+g9a7ynq9GqfEnoRcMAcazYSSQ2VgcF7QrLOch6niiqaPMbsPc
d8Xjbv6+TX51T7gI90f80ckb7q5rZz1fJa6uuTyT34BRKqqYf97783tqTGTW1ZlupvvZQOXtPiSs
5WxK3BEVEHj5nH9xaBtJK+tnvpgGzax9sa9nSkHatIqKB6FqxO2Lw0XSBJ19pOQ1g/dmFqI8ehPV
7sm3Wmrai+vZTSaSEHchFfFY/WRzAwa/6wOwGxZPSLuroB/I+063KkT3nubDQnZXkQ5nHoNp/t1/
r1WrA0ZhOnpffQmvlB7s3sg+AiQEOtUQt+RX6kBklsICMngYnhgcvMTKJ4+qIwTOP8miyWsA+/pJ
iLmWfbtlSxRA+odto5MQjtmnZYAfzPPqKl3uQtmH7uENgvliw72udBAwxMADN2rVMeLVQH7ZcJse
Mro08BUefh/ycEHwVkioFzjlqZv10Cf3ntC4t7iQ5f1c6z80EtskUi9zUbdA/bQljiPTRuFnY40L
nkMqjV/cWE0pvkNz9CgOyxaWDQsGmSTlOlCE1Ufx+OTTLVdh4/XknRv5cAGsZX74YvlbQa1S6gBY
xMJtIzakp+mZhIubKlapq6XDv8j4H7lbxN7LJjF2saDjWivA8/c3fXty9e38R5XGp/4xPdVtUfE5
wnUlr/je3yLynugNU1IrECeDy5o6dhrOE7f/0UxlQZSyIkoIaDy8S99qyMjwpVBeaWEI8FvznvIM
kaLnWQYM50fT37o5hgORC5ePXqcbvXCMCyExb4gsigslou+ZjutEh2xpqhKhU+h4cujPJTDNr14p
Pa76cb8CXb0Ybjf0qCycI499rA4eT+yYtvkbONZzjGvacYfRs6zkevNsWCBQWaEOdJhliUeT1dV/
smU229i6aYmj8HUtuGe0+U5ZaPGZRcQ9mqQiT8kET/p1XP4NxCim41u7VC0d0LVXeMAXFVzK3ePO
T9t1j+RyCRyMVIV5CmBUsFoOMZO40N5+D3/tnL4thkwkueb7h1VXpRMCfUjTeMXMvnkwyiF5JkZS
DvcKm910ZagRK6hC9/YYq5P743/+2Xez+AbECruiT/irCpjQw0s9wWyozcqIeg/O+58gPz9H+Ltg
WX0qCmaw7r9FcO+GH33HKyPuzRaf5jcNhw03OhPTXGFv5mg/LiOjFrc8UjlzkOXVUUhmzGmHeDZR
TnyNxP7i+bOzUvayg+CflmgIvKQujnWxnTaKMGe3cn3okOEO9Bx1nPW4igJBKlwtuqP7opyqpTSF
IMOdEEZe6ff1MVmKaFF1xB2RFbiOP44ocDDW2VwNFaTJDviIhWGOJHpZZv7uHM32kYAzM1aEN4Xc
PSzf7cejB5FdnQtFMyQa7625wPY5srrt/aBt2X+OLg8bKT8x+L3jsN+aNaQKZezwxaldQHrHewOp
oM1SuMc7pmw+lfcEEdS9zQYEKKxXNWYN8fhimGQesuTYKxaTbbeyVO9hbTNN0EL1R8SMo8QI+4jH
USaNHa8hYcQMxbtF4T6yDo4epYYDAne8I6SUrg8igDwP800xQQSSVAHB5rw9n+ZihG0pAEa8XK4H
C+66aoGBKWCQvJ/wWeqwQVgtB4BoB3yY9VoMSRHDleyi3ou4vLO7Oq+Cb5fWSLkhuO/At0FRfoBK
obQ/aoW9jXSXqAiM5olIYIqtL5bhougA5lmavLRjNC3swFusSZoSxMjm0XZcO89zXv4+1AsJZg7N
+Jlmo6De+zqGPfwaQqOW2WI1rbGyCYa061i+EZ2m1W45Z9xRyp3B+UokLaeoRGNPP0dsAMafV4jr
1voOQdH7YIk7Zx19VvOwBTE4/wnxPt6qZ1DSeWMCxFDSDCwhrdhxb8V4YISH+ov6vdpJ8QMqQPCM
k99Ork1JWfaLUP5TdTFeyy+rvEZ6B96tV6658CTSsBBrcBL4GAFchiIfejqOox8ZmUZ9KzOQVXNw
Tu7DiINNY88G82c73WBg1OOYe4wTyoa4JMN38W5bz2vTmQ71+yMGJ1wWdIKJae3NkcigVL7yFokk
z/rFctY9iFR/P2z/5v/M2BTm2kZRXRHVsQc4cc5CmQsaTqzE1FTWtLdg1EuuF/bbrq8Wq0qZOcEY
7ggKI+iPKC/mPTaRrvEXBV7ZhkYfRSRBizUxd2i6+1B5CS77P1cdxnJtbqh5UWFxFdS6+QEDdF48
dWWOR3U84puKZHYjTfbx7xyV+rWubp9ZeWngg5FvvEgHeLT/nk9IMJ3+3q4I1gKQcKE9IK5wmsAS
qDBLn8IAvIpJdhTyL7QVeIBoLyEaIkq33f/zkGdYVOQ4wOA7ocOjOk1kNDhe7GnJrziHX26jclTr
trbMKqcjvnDLEdU2rZa9EXXSIUqqMGRYHMUGNhggXoEQjr9+cQlavx4XxYYrdmkRfaxWQb5Fd1w+
Xv6o02D+XF95GTk+QeCZiOj9KSH0tuIEzHig5rR89eC5tMETdnhlbp/t9gujNQvcybJaBDEXX79f
zTL5Z1DYV4LGaZtbJWUz3Zkeju3+u0zkhVQCrv4FArjz9xdev8qWli/UgIdPd4q3DXTaaV6nWaaU
VDchvfHzsCMh5+kbJmkehBZbQ3IBw14fMu/wK8hdcnHwhq3sKmdHKYI3lgJbIcT5+3G73Ek9hJ4k
5s4OEErBM11FGY8ztbJ13OylNeL1GNTm/ZDaEsQHeCwPM8zIMiDkwpzQzr0xs/LPii+8vj/uX5/p
HghY5iGK4ira+W35CO78NZc2p9KCGoSXWvKqk5ECMoRKYWgOtiQRUMhuqaMSOO2/sqPuYGz9l5I5
b3xWz+FRTHdYySVx4blE68Fh7AqaOUCGASwQ+lp1uRYy4Gw6vgssJ4CK9Pc1PSukgETluW5z/5Sr
SptmZddAVjlTOWSx72uydBz2maf6RXeFQnOl6QHtTJalM8mhSj5ZZ6TY022cCtcZ0vrhDmhOzNWD
KWF9NvEgN3TQxiPWTzzWYxtnbnNU+nwxANvmQtTyw5QqbFHYRE2YHmWJizrzpvtPSzGm9l9yZHJ3
TDQ6dtjOjeFvV9dOXLpI8tcRPiXek9LxDnaEM+j/vys4qymFW8QUxZomZF917/1k78bj/UQjrb49
7PAJA6zOYCDfLYC1eHvH9z3Q8IJd1vEUnsx841bVmU0anOuhusifkp2HDlHgPxDEBNY9IeW0ZMJS
4CdNW//z1+Zip8ai3Bd9ZjGaKAhfa3gQMXxsu6E2oFeDYEyOXvEIcwhe2LOjwboh/rSUhTYX/7vN
0gUle9GWqwcB7PhqIazTZR2viujaUyCu89I9Y0/B5rPmzDmmU/GiHEEbwqGhUM6M/XlvTrSrErhV
Lj4ISJhhsJANcWn0HlCo8KV3xB5iJKdHUDwKlt0mThs+XnvMtb+Khrvtm/kiDOB5TB5h/izl7oDP
KdsRFviaZUvaMsIUtnCJnTNr6KvikHs0aICCHzDBKEI6jBGQwVt78WFlGhWd6mXqMDqn5g9dd343
6rGmJrL70YjmaKwKTNagO7rRPha3IJKgjISBaHGUuqpP24A4tS8Ys6TxBXYbmrWb/F2rTH+xPa2f
MSdxKkKXtBT1uR4vy0XsgWgYFuaF+aL/dPcErpWlJz1buEKAmshX9iifruRwFJP5dE4kJ3G3+Pto
UgXCEVxlbzdTsLBkYbIcTF4K+37IcvYhUdlgv6pdM/FKf2PkYG8oRhd8hA5w9extc3TF+sJjBrGS
38cHrG1kb+ndHa5uXmD4zLTHEpXBksR6qWJhAEZ7PoFtmv42iL4GsANEhbfl+wChb6AHVWU/PwHe
AG/jwg1+sBQdLSO/qtHDQ9bQye/BiooGQDNIGXq7sYclDjnW+tc/tuT3pDwrsKgPev6f/W7Sxhrc
FdjDG5ilnb/MVxR3VkhBjPJH8O9gJ+CLEO0eRIApKk5ItP/tCagnQlVLF78jyQQOOlMdz04fU2sv
4e661DJ50aUEuQHpke9iKb5kdE5gIRN2F0yINwpQKa0JGYLaG8H8BeMEc8eTPRuc5ak2l2cR56yZ
2ED8q4M4M6VkGcvJm90pW0mg1g8qs9YMR97PmsvtsQrvAQOmVdpj2mFhGgsXSSzDYHqMm8W2SSLN
p4HiooH+hDh7GUdzwxHNdpsYonw8eKvosXiCw8gOtvlhocJajxgTwNJ9cziygbJKGMaBVxVnBOIp
j34VeaJKiVVnlPwHUahj7WC2iNQSqhCp2L0VXUlt+qF0ORAg9d2AnC2b68xK86Qf8n5+xYu+Q3rJ
qMtzmeEx6/USZarSOFW9Gv8NwFcjK7PJe5jORcDTiMkEism+TaM3gs91qSPa6j2bBSUmEXyZkjfM
WgfRw2SFnF6B4aYX9KuzgR/wqi/tN6fxm1vLGArpAKn09K93TKoEi10+Kyiz1k9xjGjrIZrzbdiQ
H9T6wMCMKOdVmcgWOn1a0TJzjh3+yiC+yg3SfZHcYlKD7J59YnJ7I01urK+YTLfeadLB9TkgLivU
emik7LYjll1vZHV1RWJBiRlzuP5JtzTYzMQc/ZSgh64f4KlwGmvhOjFRefD2OgnIQ9SSRsUQZYBr
kX/AcnORtInMSKe0VUfvX8/4BWMOj0xHfFuUrc986S2uVkUMCffL/rKwLPB6epDnwGV4E46om4gN
mFb1m8Iie1BQ18WmU02gPaZtiSkge2PgMknBe0T2oeA3wLsgBzTqd1sN6Da28saSBv871j2xWpXA
omBoNjM8YDCHTAFedaObs6a0/1bNcge1jHZG+0svtx7RPrh2J4L8ouLgFryk9JFWxtSfJ/At3Qiz
q1z5nAcNHIO64pmyliOr8kayPIu5IP72fDZq483UahFUYqgT0P6fNe94TlxaJROieYpkwR26Kb5Z
+sI7zsEUK4ZVAfaOYDoKCZeswyLbWdS4OLcuLrrJj3mPZ7Tg2LPquIxo0DoBamOd/73WEuT8KCh3
2EZx6QZ8vq+Y0JXZxLcvFmLPo7ibz8McSIXS18hX2KV4dDiilk9flTjywLBRMMIW8+fn6Lh4uNrq
5UoMPpSfao27epnnj/BLLq63B/DyDHGOjo50R4w4h+bU4hQmAoZ06V611wVdBtZMHTg3M2mw4e1X
SG3b5xD/BdcXG3yV5tPR7ppqCqeYFQ+PKmuZ/rdxtXa/+zaEmgH2/2G9KeKEYrF+5Svg79EtxuxC
k4cRFiZS3bsK3KU9Q9egy2P7v9A7vKhPnZVcABFgPcrnwM99KsVL22xxDpIrwMVB5tNoYvNxUYVI
yDZ7eRFuKMfJca6oJkwLkQI7Fxpl+qTfOsqGqx+iT5TWFSzTr5O0X5t3bxYslDOx8t+x4Idt27Eu
SFCi2nz8Ctpvj9y7SYkB/QEGL8KKGHd7Q5Ou/L3B46CP03/rT7twzcuQSFPec+1l+65oDeMveXcX
xdeXqVDyxS6UOi3oT3fHXS4ewOYHSlXFfCfqRXZhtOA2amITFIqbcJdNDqDlfarlNMqzVe7NMoJk
vpQjF/Hod8SnEo4smXMiS7xyk8zdolHvznXXGtP9grYIcj0ZhW69shbodaTvUHNBLCpiXnrdwOhE
sdPRgAzO8VlsZGeP/u3KcSu0pErn0l8yLVb1wPJP1+rjYKacJ429oALlCRsQlk2RZZYsgDI4Lvx2
Lb39/SHDbJlrGyhGo8FNl3NuZI7JbxgXqtJklNzd/imnuqAXbsCsobAXYsHhY/zBEB39eg0UypQW
3S4Qb0CwqvnfFyiDXu+Wo+uh9qtcHTZi92d9xdXLZzKvVMSuEmvwgBN5geG/vH/7Xf+EsCQi1zTi
CglHg+Ntnh2B4FKa/5uoY5F+NIWfss36VjAqePIlCBiwccDwII3PdA8nPlovCK2BPxErE53IFhHB
6pkK1KYdeFs8uRrcR2L7G+mfAA7Mddte7we6LbL7ajXYKoU6jSRuN76X1odRO/bB6ZMqanV04JMM
DSesdGGeKr3fScCgBm0pV6PzHtrEEBtNncjIFmlxqp2cNg6nshWakKPKIhcPu3Yp6qx0Jx6fPKbs
4mx5CmN235SYd89ZCt61vkebDqUrXxP5bEgBG56IKKBW4qJK1UKSdbXZJAzjYRfXGfSOsjanEb4B
EbRncT7XCN1gwid4HCna8gf4+W92239F8VMG+XLGoEHzFOpi97SgqqQvQJm/bXoMvN9oiaMd6oQ6
IVmfU1k3FGJupbX+FsmtgvS4vV0I1q6pNao7GTADyKMjIj+FNzPKyPSO2FMIl39rKdxqXDqcBVFa
CUXFehpGMXuhlqdh2hfskXKJpbM6kHghGU+p+SlsPsX2AqiBCxCWxlyMbicFdSUtdr1ULSJozv9N
k9+YBF+/UovwJUkNGxtFtxmGmg/ZBxHa65C/tEDO1yTMikNIQS8PjmT17E4duF7+JL98n7gAFQYY
eBc5UrIbV72E/yXljQfnUBDSM3Ye7ghYGyzueV2Zbp2ASxi3+AE5oDExEPAXuCJh7HydEtwPg73P
aI4Wnu/sH9LjLQ3KdF3MWimnph0jRVjKdB/FhdeIC2sHAC/YfEdyFr6rACLpwESlMbKCf7T5yRw3
7wg/xNWj9w+Q7lUqsR3F9XUnXOHTivmqBmjMAIFdpWuAY51zhw76QhC5AE2O1i0AzbdFUYjMuuch
ZnyklWJBorcD6flmDVqdfNEFn1Oeg6QsrGt8XrdEU//hpPEwaVddfj4H84n1wIWVfhncwhP4t3ew
FQaCv4maZ9uD1G0NMCiFMBX/uilIeRDQp8Imk53ll7JstATdh2f2YtwkDqcAZyuoCjChWITTxdcG
iACs8mqI4XN38SwKAoR0cGNM6fqhUMJ9GaAGi2SZi8JB9NN4L+Vq3txHW/IeeIDMjg4DrySvAXqz
G7OGYjtjCD0H+NzrdURMgnW4ISNkHdXBxKC6PKZyMOdtw9+uPVjOBsQAjck4hDwCbae9Tcs0fwgv
ldePtXrIsJnTafrjccdHjUd2LUkvgGREqHLZDo+iOgmWAt/uOc3jFAoU3iNJdY83jX6EhrjcTc5A
KqdptoxWM0RfTpPEG0eSqNyulRmsw5uCrD6el3feZpRpU3XhcnNNA1XesxRE+SDhxZGILxIg+MQS
vfwl9r6Haeo+amkc+e88vsVw5fS05FJ3yMMkmCyKVWChHwd8YS6Q2TarIzbLpundf5w0Jm2LisRX
hdc4Z9KDB5N1EDhJ0HpRL8H1XxRv3IaIE03namQ7RXyJ6txpI4vN9I+2xwN55RBtNFHlsa9cfguR
GkO3FBP0d835fWGnhfTPG0DC/gP95WrIneLTmbqXB3+zL8lBi6Jk9gTj7WZOu5F0KBR6bs3X3O0n
ECJCDc2L4hs1vgH5BbbUnUyMOK/MH3TyXlMxpvZoAnH9uMFUBTRer06yvolBxatZ902rhNNkNPbJ
z4cZq1GO9WJEVNsaV3l5JnuNFHQELEDL3sEJzeMJ00XJTo0RWbBnJii/VaPrSyKjMNrDY4FNQGJl
ZQ5RWa0Eg4O7p7LkMUFWGPXtU1BtC9h95uhHOSUOJ/qMhdhGbkrdSeU/LL4cuad7hTrdd2+w3XQo
5RQlgRd9NulJLa1cLCQJ5B5MSetHaDdUrQ1pE9nqGQ4xz08mMYK+f/hWaIvJvCus2HnHNhOE2dF+
0dzLjaa4XWlbvXGC67IcZY/BGghXtIe3kkJCT9W9SbdzGbfp6cPqC+WUhVealEVFwX41nE03I2ep
+NGVtxwfkYIosXzymHRR5BhP52WF4aqpFJxW1bkAXtIk//8766FLgnnmAHVGE41nGAEfGxVm/pTd
MDBR/69zcHcGlxlAn1a+juuoNIECfAy2aRgVgB9yqR+dBj+iEqSXTFxjVu4ChsfB7L2kQnbQP0LB
9j+PuGC9QqQkxvGR+UolqHwj8GuUrNlJemfogsCC4j6fkSK9hKxbEBaW520NiI53uQyPMnIVDakm
aextp10STL1CVlmZ2BmAwOQcxBmjVCt8dtEpjj2hxIT12Nn4v31WTYrUqybLiUbxIc9MxK1TcnUQ
R2CkTRr6wYKbR2c7IS+7lUtcHK2UOpDr/L0Cz2NeuTn5n3sbWjE0xschnTUPTghTNMrV6YPAfBU1
TUDxwDY12h2qIbVelroOijPKvSrHuo2F6vLlnGD1uDuDlJSc+u7GvJf11USjaa9gWTgfH7cBM2sB
bKHFdILQzwaUvJ133Q0BiSmzGUmahijaZLldDjK+fUaaHJFtJUBEt7A8hDkGwF1rKpFgkHdYO1tJ
FY+PFU3cEeQK6cz4REQJs7zZNo0U7dzMLQ0znbJmEfYfK2lSBo0rZnGjeoDdEBhj9mJijhCtJo87
Zi9LnrvxhLrKCoX/jsLpAi8dxwqSb2qkhz/I8+pVf0vS6ka7iEaWu/lJRQtQj4jIDDnei1pYyEqu
H/ul7X1UwQwXKcybxtlQQRqAm+AYqPz2te+psfv3vBEQooY1WjQ7k4PGp1DJBFd8L4wI6ibLn7YK
4ZuEzbfWMYE8+F9mUjqsGdjKfLx5LIbpsf/nfYZypXO5zaKRuGLpkd0XA1GoVVo81dGu2BvrALqa
NEcJxmeLNgIaVy0jNx/rHCDkHGe3hhy9ZVUcNy33WaMxYPJsH7dscLgb5AentAyf9WnjmF+55r68
oZyrkR+bvqjML+3imQqX18FbIxLU4PdH1FT/Aca50TdJr8gJ/7kFcqWMX8eFGbBCtODAeztMD5Xa
mdFHYrf6JBXgGVJwZjfyIV84p1L7YKb4/+rIIAgcOSH9yZgGrbnAHsWKJYi8Fti+67hMwuv1upvS
1M+CcdtxEqoGLY9BR+F4i877wratPUk1zJrlaUczFrxQ4QA86pysKhf8gHufk8PbHzJHyDVYfLKJ
jmvweYWehThsh0inWSDTwwZyFuaLN8ktkNBeRbOMRcHJQ5+pRz3QqyavofKu0Pxj9ctNUQyVKqi+
uF838xJb4lp7JXE3TLV+sm/c7xxzrCMVjpwiTCfp5l0uSjO9MMy0TqMfD33GGvnNZ0EhIML/u1Qo
b3Qz8k216v6aNOYb80lEncKGqrrcpCzoYsU8G6443PadnYdqqZ6OQ160tyLhPWrzTdAp+1qpRGjw
BqPjmCt+IagO+vKhH+onTROwE2y1Ifw2R/RhP+CfEgAky14J9TPqxBb18EeyFPplN8BMzKxchGpR
qn6JA81tlsb+ki0dEmD82qVXGHRw1M+hLFLTTAjYqFZqLhgOPU+sF+onxA2KVmARORPjxJinsKYD
wNOkmoZcFxZpBUjOs85TD6sO2E2zNQ39Lb8fr760Pw/T8D4tgcj5DkA4aLHSvnRNyQ+JnIIxSrtV
p6TOtyTIz1eI7LueZLzygCjtXVVG9PPab+4rWa0sZJ2fh4TaPp4YpCUfzLenOG+dK+7sXDDAOTfj
42zVBiei3RLt7OL0Xoykcudq09qcjjwpefFkj9jIrsqReHATmS97lv+nAMMQWWE12hqoSVJNBQTt
oSsaXdQC0I1PJmrftB7B8yzQ6VZC1XXMYXUiTRNR04M7lSjbdG3V00wgZt0VuiNALldQ8k0ps/XM
9sFx30QsXPJUnbTJ4mCrT2zlOz63HTcUABWVSyPTXYC5/sB03+tchoUWi0N3wTjIxHBYQ5gaxMlI
RtSzaGMypHGgIIqSaSnUSvo/rXtzjf2Ejldmxlh95A4S/PcOpzO0/01i7u24UsKmbRrQva2Dwo6s
cxQvl9HNvoWHzoj3Y7NLMKSaUzjbTlFfal4PImM58Yxhm6HqtHVimTA8GFWrRToSyNFbT7h2Dlwk
WP+JKgIkm4oT8x1l27WXXl+isaZ+4ZbfSa+YVRebTBmJ0QNRUkz5FZvCzdwH8+MyJF18NwrhtMUG
E/S8/PLOj3HwL5xOBr0MjgS3RggVplw99oWbumvkRuZdffU2b9CNiBisAtsdHxFTQoWoGqvMBfzo
q9IaRNrQcRMxuvZY/p5ja+eWVHii9cowAgIq+93tAaZOFcltUvB04cRbfwaJN03eX136bKcC6qYw
D64XgLgRh+vlAPv7FkpljTde1ya80B5nglAIgcVIoLbjaNFPSHCzuaGDv4dyMA9QIGxTJlRHZuhn
ID3KoUMMw2AGyekJLtcZZIaZnGMXCNT/5OZzlaC4SsD/cOW3eksDNinT3sZ/+e5/WN4GqWpkDW/K
7O2ejuc+P4oV6lS1tP/qg0nShZVhjszjHO89SiKuPEdutTvFv4rhBOZE+bSFEFaaQpIPld6SSYg4
YKO93Pj8d8jjR3PvWrQE4IOjltMpkGaU0+eTlMolxEuyfhNu76AyG6UMQNPaEfeyvxSEpZ8qMgbO
5af5l1njz+jd6mYHQvFhNhAtpm5aBK/GDGh1fKJyH0jWF4OlFR1+cUk/HCDKuZMnPigYFnUfDSr+
O6nj8PDsv76U7zkMB0Vcc9PMVguTWeDlvdUwK3vAjPNR3kXpytZcV7w8h8QJT07mOK+s8n26ILVm
NEb6NrzVjE8hPAoIPzGletqGqq+hwSjwn+ZnMh2ZJTYU+8HAj0+gxx6K3QxzDHfcJ9TAhY7F7HpY
zJr7dpk1fp8nVzit6mFIM57FY60jtveEvOvZkhpfOpHO6GNy3gbSiysVobwgEtZkF1DKbA/RJD7k
om0JlIg1A2Kjn8cgssQAYP+0FwL8FtqaJioMMJ+FbzbXM9xOR5FAkIY3sgmvwqWQamQhCbdH06La
HjpY0u64bdM8ueHAwRuawedolZgEl3GU2qfSPbjnaXEP5T78Xgh8yTDnHQVm424pS0q7CYzBT2u+
cA9credfKi3z3DdYGb+wtUMBaMrFGkO6G/FSnncePUFCiJW3J/c15T+cJg/5peGOIqEC7C7oXb3m
nGa7TNW9G0Nrok/4HOR6vptRTYhjgdTaIMNXKGUsCl2pEA5i3FHsPwVoBbCCbCgVjTW3RjBT4LFH
nG1D07UMGYFuazNyprEpe3qVULKMsCbUCJu8of9MffMf88VUfuHGn260wWLLdmi9tAHSGzgIh3og
SDtjGiHgUnlAwDY9Ih2pn3zguqKwKqilbKuN+hmXpDpZKxUyw7b72JH+z4/sS7qTW03Yj8qy+Yup
9IT6w7UxJSCMk9+zG7z9qC6V0FvUtPhAh81Am2rTZGnmTK2FZVNpQH+4d9rEge+0WZW9fvbhA0B3
RtqW1KZzIUP7r2RXKiymqCyyeh4jetKmMfrAyqcrdCcPdwS5IZzEVUO4RQmkrTwNPLAWCfXeEn8O
oxgOWt7wYg5zxN2wf4INIiJ+laSFyUSgcDo9mE6RrFfhFNehZ5Iv9Y9TktTmZbpBNHr5FifuM04V
r14fx+UmO4HQs0eWc+P9UjuQVvW3rUS9xOL5OF9MGRhak10rdOXl01w3Yz//HLyoGYOJCE59wEM4
fhnuMK/VR55tH7I3Hno+RTpgQEFeo5Bmnt0/AkUdCNa5BGOuH9JqI5U9kascvI+kOhZZVTbZZTdZ
8/EBagIr+wMTuFP/CyuOoa9Io2PVmDPUmMZybLiMmFMPn0xkkEQLhKNry2sFPiID+BhZmF+4zcXy
rCrpvqCgf0K+8d3pY3V+xC+0AGA0SAM68EQvpp4YFNLYf5DK8cpfvmCHdXs9RKY5j5CxrKOy27Ym
FmN+G9q5z2HRqivuAovGBKVqGu294XZSjhUjsO+CofHLjvjIJgNXhkZXJycEaontvtkW5ClKMyJv
9c4LUpuEdSV9oMsLEUMZ3PccsTKHJIu7gPAzMHOB/7sn7Z9pG9qJs4gPw8ToWo0FmV2YFw4YeUs9
hXeaJeBUei7A73HwWAuglHpna7XVqOLwWMyGHZ9sGjL/wxg9FwNlee/vjsxP3hosZ0wsyfTYM/tU
y0ze/CPv4RU8QmhmbnHLm3Y1NFL+XRb3rH1xW3U+fSJER3DKe4I9/b894qxANSRZ2ET7gCG4APTf
ZHHmNzeap38VEa1QlK7leSthoPGLzfrP0FM+C1UHjSHFlM8uvOFlI//aTYfAq28Wj//avVui76Rd
eIo0VAub7RlLDCiz6kUyBfsimD6X4pYwvmp9AvMjwcoc+YdyTA2iWIHUAniDAWXtHYu29+I0O3t9
fMvLhAT19MX40B7osasLuFRJOcHh4v1mh5xIp5v12FUVD//xe+so6Z0UwgT2vTJq+MyjmMizU8sT
1cruD1Eh1ksbXDdJ7GYbRw+OKZ5GFdIiQxqC8O1LuSOzbg+uRELAoqjuvI8Ny7if7ND7S2QQ8t7h
ffWxKcH6vvFq2Tmu11iYewC07wf8pPDX7V3BY1Te695LNeJ2yZa7aesE4ep8Dw4LYXyBu/0Apmwh
folAjOPZM2Sh87JKSPyv+CWxqKkpQGLcPMcgNlbSwNWFr2y7uNdTApYi90vltzhAH9gNbBCN9aYo
v4aBR4iKqYp+xUAXQH6XOisBiTKYxYWN9ZpOa7Ak5LPCIDiIuv8xiZ/bOSzo92K+ihipt37H03UW
YJCL6kxR3XReU62PH//+Fd68bWzL+qi1IQSm+sGHk16vkkDWd+QJBDVp0muAJx23LMtd2FYnbYDo
R3dTIVoKYYTUiqJpmvfJhqczLFDekamozg/6MilTEVeZj+oXjf25P972xgxPEJ2K/isB68WHRxHv
s2PV5dArOHTeE/m4HU7gAF8HuBdSj5XM4ruIEV4Lb0hfrndIi1VMRzbaJbGrK2R2eldurwzmakyk
FirdWnG7ZGWB1p4U8Qh0MP4aSFfsyk/DjWUesJiYSGH/skEUTQNxF+1PV+VpSWDvbGskzGyCi1ei
0Csh/5gOCZXsi/6FAWs1tlOTehhG3EWVdgDeqKWpp1s7FRcUbdys5ZjMEYJurUYd9S5YFqDypl7m
q5BIKoEqsUC5cvPid87WqS8CZdluHXdl/44s9Ew9Td5PwKhmirfUggRjQmBlePIW0YSU4mbsg2+3
VYMfV0ZjiNEf9i2g1W7X+cRIwmh3HCN4/1pvADDbwPj+Ipvs+isTxXrfHLyeqOR9w9yNnJTHbb7Q
/OFxVz8RDolQb4DbFoUl2wd0V4wx+SFn179YP4XeP09X5smfbVKwvGGD/EqwT2oxhaa50l4xSNd0
2FwYZ7mBvYhdJZFtYD0c9Eijt4371Ri+RA1eCN3BEjfnwkZK459uBUqSBW91ntVzqNiS9Igu6acB
6mJS6MFnhiNGhEbEPhdTcmcWbXq64MOh9P/SjdJ1nFM7nEdNH0V6X9hgino+JHLfTsQCSpXBhDUK
BkWfJ7UTlGMrpLSnB9pmtn7qVdO5Nw+YduchW8RLdAU1DaDito/6/GjdU3HYJLp/wPghMlLj9iTE
sB9Ff7T+VHvLimoAiFe0DZHDUttZq1CCiab4XADzTsHtJJ/yBqQ6gZEv0/NmT7yBbxvsA/EhHuyX
WheO7ENdoFC7vyaXnvtckfOvCakETGhaGc/QBMoAG5jOe8f262kcoLnEvxmlI9lNlRKAABe/vaef
HjM72ozhfI+J7u58rl2gF+LEUgOiTuY2bZk2jnxB5gCDactSarW2Ow3M63HiSeycwJtZIkK/CVb3
CQvDV8TmU8zTvrpW0rmMQiJcZ6eMJLvyL02ms8b+5tCD+tatJUs4i3OH3JbBh2brdAOsLiaXBdX1
vUy1m0kEsxCPz3vk+kModYmsgvh0+PweffBEY5dyGmz52Wu0gGnYLLai8t7TEZ7X4pODCQ4Uh6CF
SHbOAEi5CsxRgAazJI6fX6HqtXaWfcCyE4+985dqswfM3gcsK04MQM1N1VHZZZ+bisMWy4+51TOh
Y/cXwmmINy5jSAXE33V+uMYDn5SV+aFYRQA5q5hxTfFPnJPc6bhtGv3nkYJ+kY19KAHW8849AZAk
lUVKC4EM2uZB1lL3Fjl0YivpnwNhT4e3HdvygxUofBznM+q0O3ugbP//TmhMFZ+nX/+jCJlHV1dk
mOiKlnmo+Dy6sY4FPxKNsd6BZupwU3yLVaD2KWOgLrAcRq2r9gKzU1BYSyUSR4CtwwzmfxT2+957
Y/87BluEX8zv8IrPiR47EsJWYIWqz8CHBs615z7TLEA0GmGhu0mJ3+mCMLfkilXVRxRY9CmAgb6I
raWOQRlR2mm2iAsXc6D7wQOKozPTpiHg+6rMs7ws89QvPCmIp1GB0cnDLfOMiA+1r6NCGeLIRij3
WHjFIQ2O57Di5eQtgUnHwzAm5/K8+UMyQk1BOR5mFX8zZxAsR0xZKoYck3qD/vNhznm5ujuh3Yt7
Gms+bDpaWRfg/bY5/OwtUB8ZwZOXlPs8LQSYTIOXv48F61H7gOE3BoJGPssaydtf+fTyPNWocN7E
tIYejqpoJIKs33m1ZkyLBzfcreF+R41VEAy8IdGZ3pYXfIM+XXV6aRCQKj3Z5R28bJT55vv3dU2B
JSR9lRDR/7b2+ptn/FW+2TphJLM2ebNzHEQyA7MG1rZcAip8s+OfZ75kpkbr7thlCB5eLxFijPx5
BTMiu24W+Y81GEwJiTq9txrTJBwwExIaRyswG/wcAz9aQHc6+p2my79Re2g72IbUW0kdltfrAi/X
XMyjC5WDmpYNylkriXBtJFjFHgWN4LLYaNKCBvmbG9EmrlcbVBakZetX0mHoblq2hJTz9Yxy1cT8
wtXPEoLDE94WbmQrrASXt1kLpPeLuXYHvLPB8dqWMEjIJHJvQTBRVfWwzZza7XDnS63FLqjCbVcG
tu6TVvXwT23CWZngIs6/ZcDRiUG7LRrG0SHDWxTNlnrvmuU/V19IZHSJ8Y2gkZIgVR5jJG7AzLJg
oKUUi1sEKLhArqgUAUw1iJGnoJs3uLe/1t4egVrDPzUvsC3CzPPgOCtcvgCbkS/YDA7VZU1w1pqB
kuj69k6nnjG34+CxUlozhGGgfWBlPKZ8Qp8nEtln3W+wmoyOpNJWtvQRfS77JojEZA3/sNxfycil
cVtH3ACqGtHsJPXlIxNFc74yH0T7cYdFIuysxOOVzBt4KQsSvAcg3LOUUXI5MviAjZ4cpzZKV83I
YCx4iKNJ/uGluTDREzgh6xSXKO71aTOk9k6Vd9cApWma3FZ/0yF8IyrfFcpzpNmBGyeAFr+7wZez
bFn5YI1K4mP2beNlLQI7XaHYExcBosrTZVrIqkakGEQ4uCfkbfjNuETkrUqVCtuYneyC4HSYqvN9
D/zhcRYdfKe78LwdEerp/Yw517jzAip4QRWKJLpnbKJK/xKj3qJtwVfJMAk5VKZedg87dHbjhN4k
jucDWq+OhFsDe4d4diRJlfkZvPKtGcCs5njl4wyrrwPezoBMRAFnDCKGAGP3FIHOc7Joi3WUe8JZ
gVZfA8jvMEXJk2JfUQqvgRw+CA36JTc0Q9oXhSBhmJKyUVYOZjgKf1HdkgvqWTDoDw82aHKFMk+k
jtgUznnNn4H5bOnMv9jZnNdNurf09j7cLjXWE2j6dRmdkt1WQ+QBBq8AWpRrxvCF8g5P/Rbwr0Ah
bJadeBiB0dkAD+qmUge6EPWZy8lNfUfgnTIEJAZdCGeWg66ZKgpfPTPqkx2zyN3rgShfqxZooZbQ
4DOczK0aDSBdklWMAKJQG435+wtI578kQVyoCY43tAYO5m2sH/0FPcvLTddjU2shFLg0B0Fl2Hsb
6NPwLoy74V/y5eUYEf7TR8vVXaO3uUn/L4Piiy5+JlDsUnGvNzmgS8N8IstakUeVXhBHRwjl8Wte
glxcXk9ZGlj89KeXeSreXG007MFm8AXZ+J1Xn4NPpfTrZr3yT1rra77Cc8Ca4UBx8gWIOtSQzVUR
OIDL0ofMHJDb37HR5z48sAMRKkdfzTLB3fVQINNIhtFtHX3WcyjhEajoqkUwXj2Y2CCQ5p60tgOF
ujglywDb/GcCREvpHvHKcUQuD6rNJFZyZDpFkh/vou/2xtkKpzfF7SvvpfBylpNf5C01pDIFHMzc
ZEhTpdUhQZoAiQoQNRY/w1FYlRjwRbZj+vOLUjEzRtu9BHnkNcA5vcXoJa9PzpY1vMRV/eOcw7AA
vrm09B09yjBZeJSS6l9dxjvIPmaYTfK5Aa0eyHEvilZeiZe7o/iJ9hNnw3uJ3+gjOgK8IZe0h9Qi
0l9kLG6+CKFk0/QyzWr6uTHobjQTtZjgYWZhacgDBmgstzhrxmHSn8ZGbwiw5bzPlBO271JxFvHF
7qjqDMYjyuU2H69TBu/gy8HwMc5pNf26d5yLfEYr1zCt/7be6VKoNYxzbS0kn88GQFElqfykFtOU
qW0T6FfNTJ86ctK+Fn8XCqdT+duusvWwQm+0tixWuOrrk3Pty827OUjROzHlDKO8ZzKSDHEIR9u8
uaHsOJ5ZS5D+ycnLkMp/m9xcvJlHNy47mXhO1YqlRM4KpeQpCuByGaDbgO2N9WjQ43AXixOb7D+o
pROIUTlIfW8b5uFkdAuj3+/1PxtZ4CQxBwPcbDnXJqTG/U5zNO8+v3P7YdZCd9qjBJvQN4F8RjaL
d8DAkwPueH1wlp4uDjPmfVrrzWbpJTqFz5OpCKSOUivuSDEBQkUUH+yCSZDWcO5sWL6M9n2t7R8R
LN2k0zNc+cib4k3ovs5PzSAR0UKqMooy7IgNd2O2DRmOSNcslUhyQ6k7Ekytojwgke99cQCrlnmF
+4RDZmhnNZAB7ucYtljoGsy9G+tx9HE/aUnPjN2stlJu4tvT91Zh61h7DHCUyx7IRrhBQm7rXaYr
442l1lV3rgD+5wMmVEv5oK0uDnNRdUiaWW+WPN5nE9mWE0GNgfZsAUT4PIQGSJr1UosBCZT/oBTT
Zvma2ZyzM7HZ6jUZ9Awkoh2m6clACAOnvha430xdnTqDFsne+jO8eAQJcskHV5+dXuU5HQpsrc0y
1w0prwy/JwAwp4aJ419U9kkSE8/+Akp0Aj72TlAA/wtwRouJInYxviQqEQgncEIwbcwQf61dnpXl
nTzqwODC8TlH96lR11z0LgFy5fhuQgBXD66kWnXi2+BujfOcX2AGJAgYLntRYKkOO9ZCWoIfh77c
9TFAkG+8bP1Izkb7Cc4eENzEcaEKRpw3yb5NedoE/wZVaaF6o3voXTQoIA8Ve3nkRzl5l4TqzMvX
MncrVLAK/NoCAtbw6HUcv0xWBY2FA5+hSQQq3GGbScHSgkeKNkWta+LJPbntuYxA5nxckNnr6x36
qx43KbTqE+sa6N8+gB50bbxrOghZGIJCGZD6VY3mhK5G9tAVr70Fqh7NeQ+tGKWOvTo3nLGhKAMn
jK7xMOYbNIGXPlWs8CLGg0jkdiTP+xZIlkdS4LCA1eGfL7t3K+mbrFdGCPfcIlQQqQ/wMU6BX4c/
nIRQ8a2IraaXcoRRtw1fB/xyV7OQur80z+VIAI0+lKvaGpKMM7QTuErlSZd1sQb+go41CKNN+R5C
HAk+lTQqycoF97NCB7GwePNwRX9PvBd/UIWSL5qnvSbpFb8lMugHw0jS5JwbOyPkqLSSPavgCboP
2495hH2hNMWVADBZA7Ms5sgP1/JgVVkzDFP0m6Dvug/wBg0aJjWBbchinfTpv9zZ1YOjR1IamiT7
BITdRJpstGO9tYRokiofJEcOseNr/W+XzO3V0bJRmC2qOIt6RCFsR0pKpMv+uxTUJR3q0LsyouAE
TQM/cYf+DbbaNzqYZl+VquNBCYl4H3UdDISawJbHy6TsVurxS5MZdgIBUNwg7Yiw6SfZz3XpbViK
eGNhMLO7eaJdW7cTOmkqBan6GMlCe+CeF+yX01tffBjHAYEZBukJ7kmsJMj2YrmlJqYzYGWrd9id
qwEuUhTbxuJ2+0G7Rrcktk6AJO3IlWdquLHcHHAyz4/IAuoanVLEDP/wHX1QaNG/tcH30mS+wao1
AL/J+ZQ7XmCHC8lgYfSx71tkgMv5URxXO2g1RiJYR0Kk77fh3RofEWVDsMq2lRlh1Vqex6aHuapD
6oz7VPUUuB7ZnloU6R+4q5cxMatGNQOy42z1Kvj5I2F85MGXZVl+NKJOvILN1EYEPOGN2OS1u38f
3cz7vQXBpdTm6Zvmub2erEmHP/6LXBIaGIWHdBAbD650RwJUg4GbO2gX/VhzZEk1oXJbzW56xFme
SKoBDz8qmsg2k5fmLl3IdoG4qeUhmk7p+ejcu+v2oOZwI/d7DkpUFqcn0+3CGQ1Iil8aS9hS9TV8
lIhno0mNVohwyp8UvuVf1BRhrJXhpgBf3mtoOQeF07U5wViyT4FlBgg6LHCe+Lz43i5CxQQSd8Ee
V96Apldph+8W5uTkLVuiA1I1352FS5/ONGvPo7w64IIVXanLpHJwAGB17a++4db3rLdQbes87G2d
O1TYqJU5pX0fipx3zlVV4s5ZthUPAVRWdiBeuYJgPr4/Tvj4VKUM0RsUPpXYRgllUN1Ni/POCFfh
dTLuXaANA470rS86mmJ6O8NsW37DBYNc+h9ZfQfy8MyrnMQ5abbzRFaDzs9hvQyo3WDctSxkWeKZ
I0P6SsGw0xuBXd2Z+DSVGwghG+r8fe2zijT9B4gugRiWykh4MWrPgIOBVwdYHsTFPs3I7AYuIAO4
0+bukmg4lOj+rzev/nkX53maWD8lP36YOAyvmHm0phBvf1MD0MiXvL16USTyTRI4DJnVHIYV5LgA
P7jfUNsVAD5gLHcb8HDIkMStdxrgToM858gRWSynTKDWIayAlAgSqCkbP2SQScgyyh++IEFet2em
QAgZzWitT5WFFmlXWTTzZMCMtPS5n0+P9SshTlc8fQ5T1WODzftJDyPotUjyUdCJJFuezYdcOzK1
TTEtLLkKJ2qzvKe9rGRh/W9PcOa2X2hsjApUjHxN4n4qCCz3e2uRkFWtOQFzTR+q4iaDScQ+d84Y
nPH9yOqi1/3KNqbxUW7qXxOGld3rfGRPMrvip4tIjokumVUXBvu9AsQT95rIF9KtIS5XkFB0fecD
eWt5Z2n8wnCGYOSpjqNFgyXjQamEHDyFpa9lK3EtZrXA0wBC3Ee+Srx1Kw6hdxMfAeEJMgV1jSDj
fNkiYQj22udDnYyIp7QUalkNdPzp8gdUfma6Tx2/KPZbhTt/2PPmsSvUmopOALsUjy1IFbPCnERI
Sy1ULX9YxxcjbOnX6OZpimBcolCFDUivweYztAxR7EbxYuuyL85hA1xbgiwIdy55oUAyx7LCFY7s
W0w3a4T0W23GwZ8YxGE+1+58G+vrBrJuaypLMoib8DuhBVmeYGjU/nH6xMyZQ8VBFkTo+AvfdIBv
UkCK4oKLQ96jjsyXk9sMX/n1Rr3H99oHPgjjM036uo1SlKJK60A6eDZm8JAuip5Zl6rMzowlX/Up
6SmtB1gMCoi5+bLQY9yzYBj2fGB+/NFdV2Q03FqyBOsO9/9YgoF496+Km5D1F4ThOXwxTSwUciik
b4nGuTkAuzuDJZUe1F4ejn446NA3OytGE8dCGwpBLBE6GWtHvsWfnabCtXIn4PBs7olto+PTVh0D
raYDkfqnkzgdnRyEQ9cMH0Od8ZWQk767E9iHmUbhw53Ac5emSEAKk4VzKgV1WYQpOo6k5P87n0NH
CpkfTkQmh0vjw5Yt+806EcUwevbBQ+uO8puikV9XWO2Oh1kP1I1TAmyKeNdOb/Zv7Ug+/LbgK4Iz
KNyMYgXfb2ipy6+T7Lp23FL9eqPOmBHAD0aiLT4m/4XhyAlro4wh3HJFoqXkxTjEDp3w6HPMHQpQ
GoK9rK3mh6P/spg4PVXTAUNjC7QzNfaG7cF5j7x8Mx/ieCxZfZ0osv68UZyFUT3hPxHVzzI94cYR
amvkyZeoCYjmYtxGHqEukkXOOwx6q0UMQiwFR82xa7zL1V+/Eim+fZz/WXLl/PEH9fVhdYnGUiDm
32eqIBCFD4tMlF6j4KUaq9LaLulFu8qD4FER0hYWAM+4RQtqakbW49tIDVCNzvARqz5oqTIJJPYj
TcdxOJjZ5BYrn/XQY5WodJSwsKNUNbJf5yRafwCiKzJMIvdqbDe5ituzLfXHAmcNywjs1agpFTQu
Yno3PQW6uf/2BUETYpY7r4Ibc2tO3DuIb9f+Ziteb8T/MKoDXZ+ewy+lkwp07rcuEh7e6RJvEEB6
mTQ2n5D2leUMiUv+KMQsl2bshWqi+VsFzMv+/vgZt+Z5I5F0y2rki5Ha20ebedTAqZKjTjamnllh
bDghRsWYlnelgpqMnqjMnoUANu+RrvtdUu31RfwqL2dBQhWVzbd56/iUj78NzhQB8ooH+12TjtQL
aRxd9bN0rK8+Um70GkxkTY5afRVY4u+RuTQKVUNUCpv1QcZhZWijji2smd+nm3HK4+7aYhPEaE7I
xbG22f8qd4gVhbKcnnFNHQ3U+IMng/8nPlVWsEV7L66kiFI4ZmS490Io7Xt5oSaUR7EjBOaKeirV
6neU7x2yYDUA0bHvzqE0Y4X6IEm4Rb4acPwb78DHEWzOnpOrSoT4JEX3oFSGVJ+f0m1wxtekP/AP
oHTbW1D81eqNzKtufboJ+xbQ16V136C85HWqwqZhMHnW12853L2pRX0UdAOI8AHtuV9NagPJYPPn
F7dwxmIdO+RIYwLq3B6SrtSKBim7ZE7cUa24c8r0M1Ozhlc1pMlVZMR/mK8hIO+88MMwTsToptZ9
IU8vmV5vb1LjXCq1PgFBP7ASK6ZcfJ22HWSjPpNNQ98o7tyf+GcjZoTkAqxqGQ1oiOv2/7hvaUEJ
+PhfrLBJHnqUVR9joUtj1p3Ug6KdMfXb80eTCPeD59efq2SyKX5jLJkusDnUdgIILyKDYsSMhJTd
2Sy/0VINAAwH6/dORnVFoUjEF6FMOq1QJR0NFDGL6fsImSc4nwT4lxOax+ab+8Cn5uMgSbT4Q/iw
WppcgrgVO1JKCLVeHK5uvpZ7wvI/Lq9tX967DjE2AS+928ur4eaXDcfNGcGsMWcxqz8FXXFfnYg5
WzsDdlKhU/V2IyotXYNXrhRPcrhGVK7DK4eAPhgljxRcoBixy5wSbJVOgjgUUN06kJJf2SsKZTSe
snF8Mbl4gjPAinvz9iJnxutP/Go1IApVQv4fOGEBNiyT4I4deDmF3CraD5d/acYPQzEq9S6Oes2V
RdG4dB3HSta+bbQs80hmsyk85mY4HzYWoW+VnJVQ+Z+JUOzeSnJUAXGlzFIO/XeaVz6yVGbd3mLE
EKCDEH6P3icD1Gu4DhJW53vpf432oWgr47ZRqYb5Ap0WVacO4die78VGrN+JCb27h0rSZVQYYbgD
og4EP9iBpL4fr7NsKB8e2jw9lP/iNIMf7u2lQYMqYvSA2AESnsvwJa3mPWLC/4htGqYrIxYzIklo
ET7uUuSoRKcplrJobAQdRCupHQ6Iz+I2YUbugW0I0nZHxnoia48pS0AhaNCMMdXLwHmA4AcRJt0y
KlBxE2zb12JunhxGyT/PWZ8VwWmYUhovGBenE8MOn4oSH6KZhrhylP/IFig8nlvLfvNcAd1IJcpO
8qsOrKuaECNWuO3gLZLkawZynRfsafboq9d4UUTAYIm0gvBSyhIVKJxbEiDHG+ryqkljTxYTf+Mz
Bdo1hkrjs622jX7Nn/lAWCmn7JkDLTvj0n01MlCS13YvAPj7zDyVkOLBBo4kwwwfak9L9bcmaPeX
mE/mjw2vh+GcNK9O0w+wXXnyjq00G/letmZ8r9f1+LKOuXPFA9wWU63DM9sTETGao7W03ZNw+dyX
N+DWYWOQJanU/DC+CP5u9HAiUhACncGh3bPp9xOYbrpa09d7M08ZmeCRB0izOLMYzDnWhNcflFPK
PyyBc74zPrF5WQa/Fx5p8YdcgqGBVXAePsPpLwf+216eEJR5Jwya8y8yapV/Mtg7s/+xRPSzLIoY
Kt0sURpmVdzIYfDXCZXyfHhsNBuXkro2tgxCsIb1IJP34no19ujjbFR0wNxzc1N+QdIak8JqY6wb
Yd+k/t+RVFEujUvZ7etYGTwzBK0Ysa+FgJZgni+tkJ4DEPHfE3czkxrxArf+YlDvTF3aa0WmnBXn
X1Dd+60e3tdyDjuk1su9QIHcTllpIoS9Qg96TzSHceDC8HS7JrVwq8/00rG2xMCE4AIviDvPo+Y9
x1gMLNBiinCAErDO4sqD2Mi1R9xVFBiPu23OSOFdba2DmDdYoP+jpupDesIR1m31+7R4EFc8720k
pe+W3dsNuChJDQljcp3EFyTJYlOc/dIy5GVNdyspNhlVhILw5uRLWGHy6J+DbUwjDRsVYc/Okn+i
Pi9Q53w/01G58HlFYYDct4UuyACwXf9VfsNC3Gm6pNog8wfLLOdg4RTcD6SX+ZJMx/Le8EPVwYOC
/5TexXXEgJ3+ENq1Owv0+K0kcQZj55tqlOGa7rDyZMObJdcW4w1gaFMWeaCPrrtJkm77i/n65WPn
2KQKIn+LDhQMI7JP16GncHqe4auoMSg0YmjoxapH/8/dEZBeQwzRmkNKBeaBTG0NC3Inmr4epWIL
FLZT03K+TTNurwWiU4t52XZFduHPZwZU5EvLQuag12ybsvSb7xElu1Gof+e6HCOye+W71FTeJvCv
7M5IYSyNGY+13ocqEwJtk3PIANs/uexDxktQGCQYxehlIDbPzw/aV3hxp3CJb4lMWh62R0xMCaSM
8wcFsM58YrbyuRsqXMNgvbnPsUeyYJ5sUa+0Eb+co28yp26OtRX4p8OSzLU8mHZvBdO0Vbmh3lo2
09yw/Lyll4z93DUokH6dbCcnz87Ypn7G7xzpA+QGFkV/1YmZFQ49p6/ms7JUX5KsAo8XYnHM69bw
W5gPnnRzq3didCS9ru1xf/di92q9DVtKXsEJwKf8mYRdV2kHGQP9WluZMFsHrGy/0WXsZkdrmtIi
PVqZbeLQpmb9Ozll+BbY4FaZmYD+OjqT82Xb66LNJzU7qUAToSijSxDukke/0e7uyjkt66fwk3Va
OZ+T4dgowZXyhBMLCsmY2uRtLNu/2oJSjro/PMyLcocYgYkeBRG5fRugEMGtp7aIvfQBBu6MBEF5
odZ4jl0ghac6/dy+E1zjWBzq53SqERTaVpSkAn4KCNQ4H4d5X8fk89KKT5zUQo1W+rWSxiLIyJH9
kvIY/5+Z2jrZ+xZHiigW7Z+6Hr6L63UzRB5uqurD6/NY9E3aixN+gedsRJ/+4q4Y2zSZI2YcWoVH
krVCFtD5v48FsdGCenZjcXwh9LT/h/zy1Sz1f7F+jKcQXU+BKcpSbF0Gxs69IlV2Rdly7SQw+kpP
RSPcWWqdj/V5Vvu0FPu+PQf5mH+/kjb63Ts2q6oHtrdwkIti1rJrHUF5k1XEd11CY235/AORuQmT
KFrEk+EGrse5GDhjyJhjX7k0Dgwde5ADGEHoAuR6M+3p/qO1acbv+R4StgtbLy2LQZRhgCUTDkQx
EB5JBJ3SLMcPljzs8ghyKqYS5HuX8tK5N9MaUnVj386S3twAOC2reMfvqSBWfqdIOiefjwRclKCi
QDFReIyG++ssgwhWMvBcjlCkGPNE5UgJPb/dzeX+sFtl7atPt4H0dGugb/rS/P7JEplRhe/F3Xu8
/DnSly9KB7CrdUbKeayjrjaUIsSxjYY+a0arhfn5IVUEYcTWdJkOJ3mZSZ/QleASRVpPq7mQ6G9Z
GbPOK3wwkDOrLhI1/CQqoA1oEz8HgWsYPUPwayGotIppfrvqAGC82OcXjkDtw4x72/m+2V+urWCi
ILeiu3PRaoLfKOKVYPvP98P098Qipz2Nsp4bTBhDKOCUehWrAwu1DW0h3EF6Fao4ykK2lo9rnuFs
yDg88Gu9Ut9STgsBsB/avJ52k0Ab3tQGblOOB4JKYZP6yvp9uCbXPhCrQRTtQzR3TGE8DhvNoEq9
eG11ywQo8IxS1OictqbTHBILno69hdofO/ucWiZgy7nrzznLdYXB9TYk9JE994H2lP5u/HBTPnsL
tDp6vHu2uRs76N3yZzLV6i1s9vOEMCicti/+5sMgiDwx0sLt6uipjLLeyYIIU1uznbjy+LUeWXON
Van3OEklCtW74Kk9HKzCrDG+IxDvTtX6mwJeftAV4/8R3PHdLKtUt9JlNGle13Oj7GzcLGuIE7SZ
/FTTDnYL3J+l6QGVNRZ124DsIOMj7uY5NMetMqRVSuXavXYsV5CsP3NQKulkQ/dzayuj2wNDa95e
mFQEt1qwVacaXKjuosCULW+OQr2Kiw3OMRZgVppoPfm5fj6+YYdMhjZjD2FR9t6cCUCorEsssUcF
KVbGEmi8g0Jh3q7FHoOVZkXez+FESoLs8YdmHh2G3SZ6iEx/O+8wru90nvid9X+Q5uo6UuWEdOog
S50PURJmNNa9q3SzrTegxs5nrO2XaovIsZdQoQ12rP8cc4ZfYuCJXLaWX0eBVXKMdnoCJUdl7BzZ
o/b5qe5bg8xOhwN5cSG7OSuA9svda3F1lM7OPVp5Axbtm8dHgM61mvBZHzUJ3GLVwmbF+UCz7Gmy
tfu+SXmouVOChHqgWJBvhOgG/9FZc4LI6+Ph/XI3fIeVYEXC6YzFiENoVJaaKTlAhroQbFEB6O9E
FTwFcyCunWZlell1jcYIyW2b5cyAT55Hfvhc/QuIe/A706eqtg1nGzIJfNDQ6HI3f/nG3r/BOFPX
tTKXEcmsBg5Yoz3B3PmoTWHyeFsuNwmmwKE+XCMqVwmiXAagfmY2BsOP74l0Y8K/zAssW3Zfrqsl
H6QQGCUx8s2ceTCjpQ7PPikbaqLE5+sYfEEBENIfXbhc29ZokRmK79Q7dsuZF9tblqaqsBFLvTFB
WNbtXqHEzjopAWUi1J5irlJm+7JRc5ZQdmUmEuhG68ICGtYhKn0XcDv2Th8kDwY/XW+/vRWD6gaT
Vela1k/Dhd2jrs6taf2Jgk2tYgJFg8w5vB6QUz7iPSdSBx05/K2Pt7CUTuTSoxJq+HResNrhuyYJ
TMwUgKXl1xvqolpazp3wataOJHaWChsA7EoymZC4G9yKciCv4GOMFAjRW7+4Em9oqlXbX53YCDrs
SLZJ2bPKhJEZuc3Ctjd2cvV7Zo18j0j4rNXf0bvsIxzMbPaSRavRTWK8YwHU/rsLMM7QsFbdjYQH
8SQb9LwA0JBKBQBJ1eANv7hcMMs8okxMKRi/C65dJ45r1l85aJxV0TXTGTRi4nQAMq5zT45EEnxm
swvZdiZdSThJiww9CmIAiVaaxclp+5GKykoBF+BGmv6HWgkG2XerEEBi03MFipkgFSC5ZHwbgRUM
0wCCNu5GzqTaJwu0RT1NRynC7787pE7tR1HMrjsOjoLcaHAQN7YZ93nSUJIgptL+XWxCF7PkgWvO
Vkd/M2sTMArYIx/4jfR7XheSwluZHEcGsYjHVouG6qAL6umksnkhNj8osioZS3Fk8mRQs2rfEiJS
DPZzrBanqr6Jn4765wXfiInYPzrTqbPxVAGAHQTQwFyWGXu7JrOY5XXKe+vXZTNXhHtwLQKFLJfS
vhO6L0W7US8l3O+xWKWka5AFr4TTtldBeZTWmK3nWGqNR7AXyMvle3obh1WDHHK3u247ZzULPO5Y
XefhAhpIHcbwyMcaUO1wuHU6x78N6aP17+/B52q6xyjHsKkt/9vpEgVjCi1QX/6Gfh3/D4fYHHnU
9J0Xs/dGlDBWF3voJcPCXsOcLABAqPTvReK5yC8Wx4eo7fBa0kJebbHOBTyKU71xS/vC6dZupz0U
k74z53LIpZ4GIN9lzismPy3cipMFSSbXFRq23cpVlXnT6oEutO+6R4+zx0TuJ29+gVhGb1Tlcwlz
YO/53Cyem53s0AKKhXvri66eVWY5dvTeSqaJfEfhGCGrZVhq8fiKNSvXFRYQkuoJ4Ldu6JljZ7Tr
Ul9vUSo/4eO9yfYUtg5CmYAfPvYbK31h8Y+N1bvA4CfHx5tnGX7Vn27fPp2eeZzExnr81fykxNg8
3hrHBHbljjyfR/w97+wLWtXfEv4XFx4VtIdWDxL8jKrDDQdReJHJcmylV0tGZ9T2Xe0Ue1HJCnxz
GyXqNjxL3ZXemY1bykeQ6VhxVyAgonWjC1rIkcU5c/DMkIcHpN/AV2DtoHAlfihd8icVEtzlg/fR
R3olTh4wT9xo6Ck8CaA2HOZ0MCdz8NZ+kuxbGI3v8hKZxs1bFER9/kf2D8/eouHsyhII6kVBIJWI
9r2LK3WwfpJe58cX2E7P0A2Ssg9mOGB7EQDoa/xFJVPGSA7AcUCpTklFxi4YmSGqnEx7ccExP5+G
LCE7BQf3BuFR7S4M1L6IofctldRWZk+3ae6snydSKNHfzIQgoYdwllyBBrjTcoTqLCQ+pc/d57uS
286+7nbCkg9AfAynDuat+A5VyP868HvvWQBonH1bqRJcmxBPES9s2Qs9Nx+SbTtb2srNWHyim6JN
3iyiMmqrxGQ5e2FIXKvQh+tB/BxK8InFlJ6OA4/CIgHRCh2wgHn784Wy7dWobQRB2rfbOqcEVsOS
GL391D5Vk76IW38+/qxptuw4LYZFlT0Vs8rmaU7b/56CUOKaPQTzIeOkpFOg8DYLsDnC2O4RVOpe
GoHKCNithbJNZ9qLkk07Wm74zsXQHot8q545uDw+00+0RWS1q+5d2U44rOP+3UG6qj0Fzt5s1ti0
+J3RKm6VqarUN1m+y8thgPt7T1cLqQcZCN5wwZ3QNAIprJTi86gGmLdrFQwxdQbq4N1osLViscPD
A5g1ry6urLKuG5oXNz8NDAw8qqAhfOqXGIBxe9mGfUx/vKq9+LTvK9V8/dwYIuwgCmL4ap74JSq8
iXnOn0mtml38BJ+UVFGGVRYJByFC5+45VZpSRH0rTTvvZOS52hTMwRbW5KcyyYaBp2HeAH6EBczp
Th8qTXWlXT9nY8DZethxHdxVgL+CLVBRScGpovH6rqivnJnrWVtxdHVDuSEkNNCQshVcvwt2BvjV
oc39ym5c14uFBU8tKYNBQubbTmtz/v6iNJYiXAE3YVGwtfbSsdNThj9jNQrgzcYOR5bSnoUhhxBq
Aq0d0IFbDVT+GKBkqlR/HHdyVytxNRLPt+QDtfEPmmxtZiWRJtcM3JfXg38pOHS+gp2ZQVxmx0Mf
feXvXPiVXR9/4Ns8ophMVIAgZI/8HMYyfQ1EZrNhscGkQGPh1Ko7xh/lu3Be29DRGC17tZZHDiYB
6xpROY8zPN83FDAM7eFRdRx+bgadR3Y6urcrhL/TcsX2IsVp8SSJq8s8fVw0gT1uLQqUtGz/F9PC
6IrkghV8hnvRUl4EUnEt6RbvnhamJceoHL3ZyghRmOFCLX6TYZ2ZafXL2vNWnTgWWrUWBAd8Ob4P
0n9ZiE+xpin/xH84mDseknccaWG2WJNSU9KaSXENDKVM3A3ruaCAPEl6FlvhPOy/mniXvasFGmlp
OgT1eH+KSazlKO6a1gKwZetIIb7Vf7CtBEQjgM1bYmVXtF3wuHdE9cwehdLNgwWGGqmqYyunD2Xv
sYAqUlrXmLBskxNiPzp7FOWzKSPhXJZy4Uhg5LHnujqA9Tv94KC/YtABjGQskA51hPFUcbG4KbJx
+udUu20Uj22r7INzunoKG4odjuPHtFFdvJofWEnpIhnc5aOU2lUM1FDz0Fi2WdOvEI3e0tJ1F1zU
eVoqEw+6xElWgWtesRbjYChYD8QeSEbXpOI2sivE1n4teoG4MBjqXsrPOlWHjrlZ8GeXfKiKPtfZ
5x1KuJ3fnfatORUPjVqmLJhHJ5rzdd1JToMmchhpA7yaRy/094w2jXXYgm6QrtjkFxsP0HH70/vW
sLpPbImWimBSKN3akoh+YRVOmW7JGFLW/JRFgpeeHWy0i71BM09+ohdGjo0XxeKF/VwqCGMJI3Cs
z3P4uZNYR+1aHGfi4rvNaZ12gWNgJhPp1fcTtxDhC+db9/MWMmROLF/s3Nm1a8klerVArH8bAX7A
RDteMzo4AglG+k46i2LEtp4pphm4fHK1nHn0ixwKJXSeoLYHJ1zzTB5hzXad7L39LnkNkENztXQ2
jmoKE6grdnCCZw/w0nJmaQheCR0Ae58OThq7114+ikRE73jMl81wLLK+nRMSGb/XUTsAsJfsyGg5
hBjM4ewyJ6yeYF/GjLVmanTQyDR7eK3jWFM/OP1rE/ftTnjplW2oLTjnZHvWQQfYr0SJoT/A8cgz
7dIj4b8b6RoqmuQtWAN2BNK7jVkyo9694a5V2F2xJEQAxUmNLOdmJF03KJsF5Hpg1p8wG1AO7qNn
m+9u5LSYZuhX5R6Hliksysw8vX62IrK+OuM77HKijrVcOrk6zmDt46dKce6RhToT+SXbjGSF7aoc
iZfmxJNE73VP+lT2xAniwulBktx7eMY98AbF21AZBrp8hUueysoAl3QjOMDidaiaFVM36CgoQQmG
JgbT4EokNkV2UarYhB8h8VpFdFcZH6JQXq5LT4AuodQlLEG1x2lOogiEJucFHR0KIsbYD4Nf3BGG
7GACuHc/3l3WmxpGdQ799uTsvq6s+5qkVBIUXO+ZqTMIujz9VysahynVuxbmhBc7gIIkru3y9YDu
inXK+kE9uSz9KGq06my+943sgat+iEfhHD2UmSB3R1MrLFhOiSR2MjORoENe8uCM84oUopgKhhil
V8RwOYfLpsveVcsNEfrkmENhzVAJ3OU69qZ4feDIxl6xiRjVjlIim9MjLnjLfcGkAx6Qd4i2qHw0
XW6FDXimYTy60s/NLEx1ghx48exnK/qUtGFzPmcRI1ZpC1CHVpuC0a3uZY7ar/RTyf4Cs0o5mrgP
oUpbRxY3wN2VOVclxeEskk6VFpJgj0/ccZF0EY+0KwBYFW7flDL5//r7CYkodH8v3Sl8JHDPT6Bb
6z/VI2GEYw53Sq39r+3ZkaK53Xr0zOcoHW16bZ/YMzHCmWmgWO3eib06yWY7j/uYNHvyFu5iNaH8
+fyw2x9Ntx18+cZPftPFCe8ntga1iJf/4NsQnVHTE903gcvz6lSnJTOScb0ujmUtRWxSPCqixDpu
8YefxFwuItthyu18oLB1dABecmsr/WyWj6jlfMI+ida86yUtOIK2eH3f4/wDhRVBZC0ZPRKFseRO
gX4BSbTPBbHf5EEb1xavhIDx+Zx02XHkIvdVWTx56nSo74V/3Ws81t7nhnHlZ9YKO5jhHOd8oCB4
Idh/DbUJQ3K/qEPOmWtJRhz1mX13CmwlKDPGrZDYZ5r0U5QUSaDXPj5rKkk8TUjzd81yibrkmhQN
/nZ6SvjnrKFjUKTsMLyalWmZb2DLtA3QUZCmlUkwvtHjpNywftsoUrmyCJhTH74g+PO7+saVYdAX
M5zk/3cKymS1rsGYT8sibFZJ5SAVaxgAHZFPcsPkyllHxaCW5bC+imXqaoUqHI4pQj/A0eftYziq
zSmp3t8UNwLcSzNJ+K5clFsUrpavBNzwXOcUYWt+u66DlV0x/yUkiW8sZuD2P1Twfb43IAqC9x4L
Kjv+tj3pdlFDXo3+4kpx5+wlZgVpbf4mzzUDDtXCQVQm/axhN5JFBMGbb6Q4uvQ1JL+SMGzwTJfg
3uz+tbGZpZVUoLE+NdkXpszCunTqSjggosPRDioX6I5M8MXzKmJEkug1cWOMes04DYN96Kpg+VDg
hvoEDToJsl0R4K4xUzYQIdRrIrUwBVGIyFJfUkcwxjkjUtAaSHidm4NI8rrD83gUAN3Zt99q4h8E
k4l1RYjfOxau+KmfGiDSaiNyVk+op0aRQ0fU/6iunMbRRXS11tjdxxw/EVZjAkApJMUM8f7mckzn
yAra8Kte6fstt25ZXAM/YdJm72iFzxdM3mOey/4y47w2OEWgFE0XO1yRqIcWEyx+KRqxD7etis/c
B73ktxa4MJD+nhtZqDJvGqUdEWHTqvHd+sOSlDXMRGdy/bX6dA9DpxsZ1Ux4XTENgWW1iqWiu/2u
a5Hoy4ID9y8sVKkun4EUjMh59z+ODJfcpzfnOamogsI3dw8g1grIHI62MA1kW3DCwNp7iF/O5cRm
jW1O3gGZhT4g6HCzQDwwYB2NpWWB9j4uHxR8lagJsklebLguIb6VYkD8Qa+tEoZmWr10hL80/ytQ
n6QhIjQs0KE2WOU3uL/yCRjTbxvDVeWC/uVyivUEUWFm3f1437FQUq7sRkd3LVjkn1TD+RlFfYcB
KFk0aUf0NUCFaNqr8P/zP4eCnJTGRDLW1fzyU9h34ewkRChq+hJdgk72f+vFJkfUF9hTmvoMi5xE
tYeWlegYe3QEA/RgCXamGfxG2wqhneOEq5xE+qSQCkDaO+PwFteK/6WJnzOadjSAz0RyhTIpJq3N
0434aYCstboR8ZLFw72g115S/W35DquC55z491QRFegCjn6NSym2SuCbn8UM/+7Ru3LbJmVHZG/n
97qrS1ebene3vOIiqIFmHNNFNVyUn1x+5e7mMjrAYVywpkksrhL+9heRu1DZ/a6YxVidS/nCfj1F
ymRjWxDHYIv3yxYgc7ZawTyZTAT744rt4aC/mQhpR7Lb0ynulA27wmRPLTs+6nJ8NyopbsvEfmVB
tq4jC5fuvgkyXyJ9U4C5k/QSDnPhn/Kd/zvp0BpuoZ+j8vEWkqOvHH4cJHTVUoTn5U6+3abYneNW
VteFa8kO+rXro0NJDv1atWgpR17W5JozgnbapmAeabZ68pWNwkba+Beu2Tjp9tI4co+mm8FHqnkB
SZsEIlpIbyj8v4UNiQReWPOUkAlDkDSYN8hN4VoHbNlJZ0BBXoJHEIpMOhIKHTsdiBIkAf9bbUrx
/ika61BQuYJzezR2HZVovRmtXzirBFpZ/eJWqLRVhVC029dxugQq6/BIDn5k78dr73pmuo9x8qjF
gI7zKelKMadoI4D7gMFiDMxcYnre/mBet6KAS0ogKsGkvS0xUriX/cDDCko2y2pst36Du6Wla3hp
70XMajGBevKdzTgCyp9SvoKecAeCUYXuw0Cg1Vc68s8R13XPnjidRFMIm9nd1vZXHGdPpt5Ny7S6
ajzZHDN4uyVDOWoli3n5PDb54eg4GmrZN9J2dYRF2lgfnymJA4R5zxQEuLOIzL21EgD3PqwSSbL0
HTcMJzK+n5as2zdrGtoUdslaG1T9PrQYJP+Yzxhl2bUvuVWzZp8dcn98Cbe6nhgiJII/R3oKTofT
n4PL1gSBdy+JTZywH5kkLVZsLZPHVWbV26rRENxK2+/ThpjcVP9RoqBLi2JMn8ifxwU6Huv25JEC
JhG4fNkPpGJaykEvCSB3+La49iZJYjflSh+SujWnyInuXf0fOtYJDbvMSza5z3FhQh2cu9w/7SCd
jYQ6X9eTAQ6m15nJ/bmCC3mfyKi5Vg7a+gTG9bya59c8Rk/xVP0D4XJUgp376LdC3YLP3ozbMcRG
0+qAmRD47RFE5hi1Xh5jMFXAC/8Q+rO3WY//4M3f6dTHJhNJYXi2bvDDomjQesLNoK4uQ1Yp5ogO
oYhLzckVqjqgYlEETOOtZrKg4180H1CLk0ToXZ2oaMKH0VcyH2HjOv76L5hN9em8R5yhigRCv3pV
vKeFGay6zT5xXwCtcghro+tQuDOsyaMlsJYx0qADgGjIBFw71qzZQNjx9OKeH52CLDwr2J/+cPaS
GhGzAM3w1eYLK23fBzC85ZG95NWR5hEgd15qKi5aB9FrTOrCG3pcjOgTzbMaLOghIxhk6bhg/SDu
A9goxxcoItxZMCjaC6k5eup0Tuaynalesxwhq8X10SohWbdaJZ+JP5CThl2D3OhVoqvHI0zc5aof
CtYLKQ8MZib0A/2W8HqkdS2wHooDyTpWJpIsH4cd23YsCDKaoptbiJJP6p9RyYIegKr+CKVyu9g7
KQ/sMGp5qm6BcOqBfUQVkSfbcg5IWa4puSZCMQHR8Q1pqUerEfjYT7rXlJax6jiCfzxR1hJ4f0I/
A4EGoYT4V9tdWmkmOYoIUQyRHYiQt+oYFKJZkxl9fKXC84pfBwECoDCiSmwMaDW/zpkgj0vUMtoL
i53I8GLLaMoyBOZEfoP/smA4fHbagT34ZEUqMHFF0XpRL0kjrKmff6Pm397GqcudRQ1B7vBkHCnX
mDJGq+GN1NGUEAhdQlFI08ziES9bzu0yofW6CSOB0h6YOUbyFEYQi2TeXqybtAA+OpGDYgHIR1Wb
MDODd+g3qZ2sSQCsYsvNRPFIfMgjZ0zvXFgH5XJGIYD635qHntM0ar4ObRJcReSL9ly9ljeaM3f+
cyoDmGtHifYTSnH6ryehmyHiE+I1v32KIGKZcUL5hMfkuVU9Z86lTIVWJZrg4eQfU5vKgY5hBJ4m
6G36Lcns3Ci0j4qkjal6ApqnvJJxN+hpZpZte7Nbw/o+2ZEb8rSm1glw4Q082VX+jwAqzKGpTw2O
mgZjnHimKYtFFLyfhwwOUHgPjo5uyA+P/Zux5w4jrCl/C1NM4j+sJuWHr8K6hIFs7izl/taYKtoy
ts1fcBFG3M9YsQQf5MlVUB7w9b75hNUV72IACDmUdPzBaQAGN6mOtLUDimUdhmX8RMG3HbGJHLf0
1xT7aIqtnApstqLaGKwYXcugD6Sx033mWML/29OUn9rac6fOueT9rNc6SCxWMZilvY72Ub6wlH8K
gaOdVXAOkPCgsU+4EZC17mRwLxiXdjOhH7idIuQVpTfNiC0Qt2CcOg2PlAGMJWgc8fljMkAPwJPl
jGTBLfcpUs4aSeJZNDrKYOPRNJdgFdZNLdEHfpylG0Ejz1g+8CG6jwHZRQYd5bXa1ySDiDPgahFz
KaZGSo8ni5bOdrZbkPu7kpql0MqrS7IbgET/Y9wDG60GmlvoqEASNS2HjAQvlJZfaEWFoZsbrdzB
++XLWof9crlH/fDro3H2m0W1brLu86Mdf4sqUWuK4jjmMWN8RwBDlG+T69DRdp5brk+WU2yCH9wv
yYy6C1qIYZMmcEpbs0Zjs+fcYDsekKdo0y2duYPfIRDa6vT/97DBI4WE63/HCYNVOMU02upKqvRx
uBqqtgkxtYr/yz4rR8IOblTKxoxFvWBjOoyA8NGE3PsRd37MzUOVbrADVGGPo9xrX3JrBdFJIE9V
lrf6f85do0opZAkyLiJq28GHxMicVW4Whm/zTDTK9mSzwTAgxjBuR/JOY5024YbG5tytjbyj3sR/
E2gamXxzrooAN49qteFotVFJ89jTj7Vwp8QhssSqM8KK3ZHw8Rg/er7DawOpyh2IDIIjx2ShRd1P
UaPVhyJ+KUVCNf4mxSb4FDzYhmDY6ptQyZq4EGwNgLFS8L0/spRrcDPhC0IZlxV35U6baWu5pm7/
LavLP+HYDHA8mQoy8dQ5p7F/d/AOKnBSLUt5g+lQeQXij0ciAGffm1UWQ2t+PN2WQKC72FvamS06
tThHFWAq2fz2PA1uEtE+r/l2hvE92oBxSXDhRnvE6Z3CoM5+rOnC3yp86G/Ys9x0wgpwVA5dULfb
J7G4bFIT8aiD242RFH2V7vlgGYwCwwWGM0xM8ooLiqKgy5sU2aRpTN0AGh8OMIQl62kCWcNVh2vF
bEGsCvg9pf9l9Sv1dp+y5GuMjg5eiOfthsD8ikzqbugsk9poz2AG/busC9BGtYmzOnWorv+0Y0ws
XEeGq0f0i7Gt5AZkdOAMo1o6dHhta/mlHjQqe0ssOm2by6v6hc7QKOjSrfqIJeOelJ/RDpoUKnyS
bABSc3HLklDhxk3ryGTCv7FQaIJHkkFHDb8sfoHr7jo8MNVeVboAoiOHWf9lNdML5Ix5V9HWAivD
OUZdfiYEZM8xn+ycQRu32l6/foqRSEvwJkINFe0HwfxzvwK/0SXp0js90XNBqUhIQB8qFiQJUpD0
b80u815BDhHGVHZSFoIxBNJqyeX7VSONrDWnq0y9K6Exx4vKsBhkfUR5PNmm06diI6uLE7sygIq7
O5tZrwxSWOgOsWQ1K2EBNsNIH70OGC1hmmZ4wX1/cRxneOfxF9lBJYp7IxNiNsMls9nOgERkVv9J
xLIwdJGPng2QSxNFIz3ru41LTeXuOekkU7FemGQz4gwp+wElkzxt9pJqNRFXnzOKQ2KXN1clGQ4K
jY7Rj3Cop3ne/BT/dAYHF9XLiQIcywm/H30HSZVSXFT5DJiZLpzpPrxzLkjh2dLZt8oa2xDcH6gP
wo2Bom63Kj3X2M3hPAfX+RFA+RUqwJk//iN3doG+aI/6Nz3Hhga8d8t9wwpiWcWnHLdKiNNGWEmL
rX7uRlmIDoY5i2ID2j1RqIrFBhc89a9PqeUMp6ZENoysjK/Z+vEJlvAKK/Tf+k9uLs29PKabvoZD
duJKPORQDJZrqByq+jelc8+ufnfcfI+nBtRLkJ5gIGcCQMABSYEeMpvaFfVy26LDVa1C62zflNSc
q/2jCBALoIYBEdhXLPqLYLHJd5t9Db3wfIgAcjnQ4FcH066ESmlT+iZtjTuRclxgZ78z+POC1znz
Bfepz63ibFc1lGzVdti1fBfjf+nyWkT+UnCJR22Pz9YaiKMv2SPZ8hf7TVOvFpLXHBNg4yzFMGlc
2Ppj4G/a1KJ1StelPluPSESfN6PB26zc7gBul4ga1tw7M8T8En7+aA1uSW4H76m5H8/22d/7KjnD
5UJgGNiECdIG2ga1bHU6YFF4ZDW9k0aShQKNeMJHhdA07hAhI7g1ZQtJwYx6herTpyMmCtPw3Dc2
WWNQpI+K5IY/mrSwBKgq0rgZoHDl//Xrr9DaGQAH+qgJXimIZHWWxcLV8w0Ojv2KV6J3r/si88V6
vZtahZFr+gkgDF46EA37lnMBI6Qo9dVr8ynEfW7rGYHT/Zn53dCF1hGgKiZqcI66P440yMd6kEi2
nAqHU7aQHdgrMGy47xp8Q79VE/Z3c2cbBJ5a7iTaf6aFE/HnBlo93z7mrucDyN2qtkIyYzhG3AKG
qmhogYcQFnogj6wX3jXQLSqirbRGd7ydtSg5qHIJHebySGyoPTWMWOyyJd9sW4RNBRvmrpYe+phQ
U9s0EtJCz8GYR/5obdRswVvTzob+Zma4/nSKMwo6uMcSMABeoHswoZfj4um0A5U8Lt4ZjYorwUof
qy0fg+DwbERTYp5jbpI7JjyApqPlNaKtWV5dlt1xfnM3LvVYWn5zHlZHs/bVh+i/SP8nMoCrTqGU
El6sal5ayAmRJwMyn4VuqiabeK/chEz3f5+r8ZeN89eqlDt6Og4qhTj45jALGZVSmUFe9xBZaPI1
I6clkvUojFkbG++KeuyM5hijt326TRQGpeJHcYQuHN04b3c4qLp80p8ZEiWaeouku8BAsSJMgEwr
oKK0n9KagRtdEXgS4TMcDoSt9UyGQqJ8hm38Zb2vikg4px+Zm8r9+Z1kE4Kc608tFMWajrCVknz9
7NX5qmNmAtuKtEXO2ReT0VUiJ83D3Ulc01a1qEi0mx0aVGSaTMRjaIVsQ38P/5VmzYWwUMN5BevJ
7K/v755vMn8XQ3qXqNLcGssDepe6bcCQ5x6dMgAoPB+to/CxB7NOFpjaLYq2rLmJuKxP2ZPTtItF
XHdGXOT8dIw550zqKrS+pOiN/fEkHi1pXoLLSE5Oy0cr8fb7YhmcTlsBSx2W226T+kzEaxPLSdz4
ta67J5TCbglyLmAoYX0lGK4VQizboUeyTJS7JryEfMIwrQaabsBZhakLNzwPF/pH0tlNM2bxDIFr
oc45i4GERBY9zpgVzqT5eosGMIXihJb0/NEwcYWSRgnjAKAJ2a9sjuKGb4FAizo2tGyEFdCrcUXt
10ODTW7BfsZ/LIGGvdDjwYuzqjWkC7zrn1jNmwWoAlHCW4eHFTpsbHN/uJPXxVPbKH2RUAFyC0Mo
XYPoYc45Y4Z0tlGh/CAVnfHdNWE4VS5PPf3GyeA/yrBpvSBsC0rpiGDdQEFHBnOmcbb9QdNJTX8S
VBZQxVpbLjq9jwn5ba6bp4vJB8vuuZC8D8c6HjH7fEG3XyyQMSg87xdwJyODhbYbvxaTV8Xg6udf
Jb3BxV2wrI3CzbyKiIsOyiJxCS4ioAjoAKD23k99vOW2/IJPzZg/pLFjmyMvzlJGuNDUAWkCSf+0
yzhHcTDa0nsaKmpYTywX8DaiRLCBBcttVNchQZJCBOLzgMMTWpf2TzhE/z9+DlvGy5zspA2M4pH4
YxH10gnIb8RPhM2yjO5usSHe30GQXgN+hqXuwsQPQEtwwpXY59eQ6apOjDgQSMrOwc2AiAyycQBz
Tc1ItJAUXxJN+tM3VjKpsqu2DGMz0tsapSqIWE+f+B5/xK1kfO+x+oafYOiHXGqcYTF0DH4959uo
gJjJ11aRwHHrX+ly1ARBz5L1KpSQRMnRkzHwDhEnNR4AdPVJ2XBj70To0/CEARYUN2Zofpybk79+
YORjpvMJABnyT6VVnJ1vWkX0zsiD/o6dKyfMIgN4PrKL++uEIP6R8b1Q5D6UV//pdTBeKX/Vdxw4
pgEzbEysrP6gdd/7rhkwIlTQVgeEd2p1rSg+bdoJ1Bet6UEcb4dO1TiJsxqE9sNUyxKyUzJCUBlC
ub7zKth5iOaBM7d6S3CuxpJyLwnURiTNXHB52mDNUrBtRT4EAFrvIa0tZgvC4iOz4+oavzJP35Wg
IQQp/bl9yoHLe7W0W4k87oxKHCP8OpAmzphq+0adrad82lgcb7pU0pJumhy85R2jgxSl4C2oAyEs
McLLX1KCWtqprabaekeVTqKXyRA0hSFuqoFF6yeYzIl26ZVxIe203Pbb0icRz8qnAzES5zPg+Cu1
qtxfPa6g9+wOfAdwgxwZ8ARpxyJR82TqSjtWsJufx/+nVNvYTfyFfW3hl1pEwwI3nXfwRwY+xyEy
wPC1B/aPWsQNvgZ1ySLh6skkJGkAJvCnnnvLWZFyVY9n998NSeb2UH/NRRNqaZOMOcqzAfIxvsZ7
9/MwBrG732GWUr7+JghaSQwX42C1Od1LmmWw/vsQixmyVQSDrU36w+ex5ILjJsZrBEvaDkXpfcW4
ArBzDzTTlRgEfx8qv8axLlhnvBbnuZiAmj5grDwD96hU2WtHL2NiGKIGl6LpdHrWMFRUl2SGVPry
L7EGUuBz36YDpBe71gsf1qufKxlhJ0o5jxdDYZrnHbPqU/kerkECYuydXTHT/95oPe8wRxxrrBrk
LQ+xv75qOByBQ65fQ26bWnTgt8tjKQu8SH0PBcHgsZmS72Mrx8bzWl8LLANrlgD5TqhaR370D96P
rHRBHXItuRTL+OD1g4ONgcTjrsSEvT6xsgu9nK0SxlklAkbUg510u4NXFDqnsQW7N2PyFmpvMsBi
sJvo2ga/Abrl3Y4/8el3xHhpCHKcxF1h1Q2EmreoP8hywq56unOomgXBcLvxKCWsUdmHTJc9mLEY
GYchrwv/doon1IDqtWlO+HGwwd5qgxhtfPkwY6YWvGsu8mADm2ozFVoHMu3nQWsjfIIAXGAS9jH+
uZ348avikl5QfuqRK9RhPRwtF8xEfw9FYrtKH04CitOk3bCvqZP1+fgnaBBVIyi7fAKH+fxPGAdF
U2/PtnNuQ3o83q0+EjTrMwJHzfpqoEYko7wwI/MgOJJqL/5RXTx7ZN5/0KzziAk0S9UJrLuGjTDI
ZTCgbKPVld+tJWjiES6HLwqFX5yisttMvvVnRVc3YdsCs+U0KwkyNh8LsiD5J3AeBJbaveNZ75hV
UUayAC65I08GodU72VO5N3tu7eoMGmunCo4X8Csad7aNl+zzvafUQ7QvRpZs1+MQNkYgGlnZuzEv
pi0L3asCMaZppEuL8WpW/VR60NiUhqmkbAFtDZHkIFl3pmO0XJ5rb+p7SuPuzCvuEP38yhqXorhc
oiWLEkrD/G8f0gsK/zPUGYijLEAXAnGORFka0vIavjkU42GKG57f3dkSIK2Hb9+EqOAjz8gXyPxf
3cQLVHul9QsNmD4ogH7B2RqTsYGipcGngVJK9grFaMshgqZKwmZJo+sxWDoMvm84ROWnGmZ6Zre6
UD2fgzrMIOqzhXs0GC6hSVs9hIs377Jyr+ApocizfAsGSam6qfFRMwFrt+OgCw8nC5+jx4R1BO7R
Vvu3GWy52ckexrFuleto72BCKLZjfv0E6gLsFWe2XfcfF78wQCsO/PuaAnW5UtRFbYm56nt4qkOY
fXVyvJ9vHVWJAHwIX87m91d7RKxh3BQsJPypjy2TTs4diGwH/IwUbQnbUC6lwfZ3V7+UuEiB/JX9
vhVuEIT3tFOIQXUf2U0DeJmXfL5NkUxs66tPKi2i7bPlrnux23yYhvsfOQ4t4u2nXu3R9GEFjcEK
r+paWs5Iw7c9PwhiA8HT8deoYGK99vCAN45Bimx5+xEI8a3N+44yCDuosnqZK0a5FOQpiUsU16Hh
7cm055FQa3G0sYIrN0my992+xYunvDbZc/9zIIHVJ3ugz4TdvQITS9hSlM6H52vNldXE84dHxngA
21ZsnF7e4eoscW5KPryZuJvZ17i+2Unaw91woFc3lhxfxvK6pRVxRp38Laq6+LDw10IFx6xB4oy1
RXfeYxLefEmZhcwprZVqsFmqkyTmYJ7TVvED7p7Jfmc4rpxqMGCeCsE6tUW5caRBLTnJ4xDwF1qc
SDLxSiMINQAYhZ+QidqJhxAp93JTBTlmkmW0yWj0gbGnMvW8qHjocpdk4JSSZ+ziBBTSmAvTWnBJ
/JefLJQlyloi477SMsaW6t5PwKJMt+QCmagsOKQS+sG9KLmLI7j4VVjEHZFc67eFSHErqbSPG4Sz
ivVYjfnG5e2csZuUzvpRsIcZbyBv1J+tozNw6aSZ9tLWgN77Q/Inys4jf8Qn5pJZw0jOOdITA6aV
Ps3SF4o0kWvjpwFXXq8cLRQh5tebZwb/Yuu+bv0k0odKy2jIzauEzRdvHQcVVj/rynzsHStwMHQW
HHowO8GI4h2wUPyNUv8WLipx8qnO+Sf/PH8CBQHRhh8KoHyOyqWqvRJGYPrpFvNWvHU4NM0IMpMW
czzVn6BP7Hu8LpRQ/EZ+on5DWpxOe23vonthQO8fxfjr1jGDQHHFcNtFHZesyJlDIuJanE9Nyspx
vCwdzfF9soPEBvS0fNmBCuStynaR5azl73Pk4C7g7yh7tuENvbwApVuuKxJjpvYEppe2LEye8poy
oOVtALKr62AXH3mfqeRgNVX2NLXfl7WIq8vRtGWHJQuFTrit6CJn7vcX+HUmn6eriYscjP418E0G
wjAEXJS3F0Cpb3M66ogMJwZYQsaCf7uN4CabdEI0QtFVPRfVIo0O6nqPtvNqZqh5ol/QJw/4C6vX
m36elN97gTR5GrCzAa/CkzpEiUCuVc5MtjrzpB1r1eszqmeRAgkh38FgQr51JyiUnYYGlugbw0Tu
dW0jcTtWqrxyvHjNz01iq7d+Ba5n2ZTRQrqnvZawzCrzWrjMZOhaPJ2RO94mhto3F9/+cql48PjI
XlPr1gDBCkXTLdL+gtD6dS/uOU8JA/0KIepL6CRLHCW0FQv6o7UVSqDsRXLouwNPphefDFZt45jE
l5U5paxBh0oP/JOgftAcDd1ZdaJgG+dV4sjf7s58KMnHUJGAbNPZG3MbZbrNck4+n5sza0CwTEXa
STP8nRdj/faux/9kYGSOC0kJxnqFB2bq4GXX1CkJTP4FiKEDt+S0NfX6w3PGgISPeujlV6KYIUXe
eUMu3C8RX6m2IJqx7gSnZzq1blGvQxGxd3dH7NzpfO7mJC0VAFsjQryAe8w3mpH/2wprje611ry8
lCwpODj4RerWpV0rhLmJPCeq21Emfh06Psi7rhwS5A3soxl1D18jSodhblw9a+mDIhvK4LYPclmC
hfbk722lefXS9Bs0vaqcVHlFPfXWJSYiUAgeZPHOIuHQ2o3lFeE0/gNSRNgL+vbApOy+C/7ANYUn
rN06MedlzjYGTg3SfdnSSPhGhc/YA8WLL9+NXE75jKBLTes28R8/qVsl0a+NyTlyrLoeRZtvxsAn
85EWYA8+ZJMhKBaIkbWOPA7yBGK6l+DcpFGKpCWW5pOqoBRkKNvdnDR0ZPRGTLy48UjH+va38RI7
SQjGo/a+S6HczgI5xxUG6N6QO0kvePz3+FnFS4417ywBYynLHU1ynFL16gPZhidoJSjs/pCOaxzS
nxldtBuTBcr38EtSMII7JGgBQhh5pnMJD35DkcLpNx3KueocWbvRq2QMabnU+1ro+Iud8EahP/py
T9V6GhZ2bZyexY0jW99YPiNeps/mhsH+wwDsjyjRwSBpfOz0oCG6C7/HScJWex98UwMKOmwwaNm5
6VscHuV2B2EC0EvwnwNf3DcNBkI3cItSJsaGB5cj58N39HgyT/URhWTCs8nZJtGaNguv72dRnMtw
IUGDFupeHY0EBS8obsVAxCNWcr9Zb/xO5rmJZQQfDUrrRoHrn10QgeUVM0OPqXCOAcGOwiOaCWHM
7/ps4jPYlipte5mjnY8cNMlKthtB7Eb/ABCNC6HivJwdpiGeGeSWmPKgkBYJvHrYzugAJRMNM/on
jn/2Cd0ajMcriWJMjTsQdjJ+A8vjKQQ/uqYh41+EInR3OCCo5xp64gQBBtZcknLD+ZMxPKTomMgg
H508qcfNbOD2bn9myMfgVLNOvxiwGIg72ZEp8h+q8Ma3TmOSoUFJ1Auw1c+1nD5+cehSQQPZzLeJ
yzZY6mlpOeEF733uzkIPNNr2Zx3O4oRxKZ8RTr+sIs83awwlg2yxlOwIeGOxYvALDaNOIS4V7Jko
g+UH0ba1yA+aYeWCrXABpWBIbIv4WOvoFFlAsvIGikvddF1viY91/G9xYhZrFy3OuXHJuK9mS4Gd
S8ScHfjrhJNqy3uE5I7iSA1I8QvYdV1hAEy2JChVjNXAFkrQ62gYmiBI78r/4vYLW+lnOew104KO
5DtrM4OiANSwsDnUhJcnAvl66YU3ei6wsmwcyv4S/IwbTmP2OEvPwcvX7gMhPgM30/Q26zDT0qgG
HxhkjUFJyuwgFZA+c8kRjnnvdGSn4JUwdkJ85uSZbymAgchegFMykcOBM6DpYjCPayPlkc3eToAT
xMemjo15tlsoFp2faqzad1K83eWW3FR0UcEqav4US0A9chAhRvzjPA8uRyS7NIVlxP8sol9/AkTZ
cB8YHDGugu9CyTwPBsnsk9djbgUVHdGanbliHV3LAGu6dShrS8mlg0GuCxO62G5LV0Do9oWZdRr9
GwcJ3+TnM1olDSP7OuHLy8Xn39dihI8m8LU5jGyeoaXyjswiol7me4a11JSSX8rFI96Z0p17SmTJ
PqyyGcEIam4T8MRhR8mT21jY05MaUS5xlQIg5ZndfS2tuYbmFKja4csaUy98eppTs5J1X8kh0PYa
bj2ZE7Pmt7uTSmaj3Y7Awy7a9u/hCdhP7cUbgpQZ3qGEOP++9h3fk6eiNYNBelh3DCtZbCkocUK1
On9oNZlXjb5dFAO86g9i6VSAYUhsh5zF49iJtqd0H5HRxlmFBMb3kfeajRtizFWx79qBZCLCzFNC
StGn2skJ0OEszr4HFfsXDpI/qgzMeyUVH1ajUfZSIq+RoGDdkeYXGWx0lajUXfFuTvaLuP3ONfYo
RBY6a0WltVRUgCxq0NuXM/Zny4PpP6xUbwxl9WBtKQEH1U/ctOUBPUwF7Alb6n1mjdPQYz4Muvzd
T2r+MIh1o1FRbUb5wp0NSwaa4WEMcQsTYAXq605HM09a5X1UAmveuuV9+Z5o10+0bcmmeHMg5aHA
2FXtIfjkZjDY/y6Hl+fhw9GgtBFGifxqMUopGrzQjX2cPzkJhRUcpRFqHCgJ6/9Cl5qg1L3Aa82m
h7kgBAmS0jBc8YNJVOrnxSbQ5yD+MXGOlD+CqSUgYyEKeiF2/wTmMOggQvBzWEAoim/Hf7Ope4X8
74AlRqp9yIuhp7nxW1cFWYemyt45d1ow8lBZwnfHuAEJ7ueN0F3fbzM9LUUeOQXYMYRBGlbQ+Q7U
JuUYUJCqOKDOQlTnwqBDk81adtDTpZmGQgMzk/ZXzzbuT9a7TZMzZTUFj2uZ3E3ljJKB54YFYe/Q
MYhZ6+N32MLFTQqF3u1mEVJXipGTdwUA6g58NdygvBs3n2KR+zmg16FZUv/lr5VA1q3FiSPgabLt
atls+o+UhIUK5zGiGVB240f/syKv+szYCJGCD1CNHXob1/OrjWngtOFpWZbi/GIuRSeOxWZaVfpJ
IUTu8tvbYU5nehXn3gjpZQy4tBbdszuLj8b90vgrhkLp4xh9HYNbKuWY6pjTytB5CV32Sb9rehqs
3kYtkvEJgJl9WU3SyF1ifZ4fRCbNyB4yRKybCcR9qiCqB7W2I6mvC7XO0dWV0o8Ug4L/FAZIcAM8
MCxheMBdUubn4sBBks6HksjbucEod3gfU0Kx+MBHis7Ccvp50eMbipfWw4Llk5kzuxVmUEeljA2p
QMokOrz8g+lnu/8LQFo4jXeA1l58V2N3jy9N7Np/Eyo/CV5qOKMN/idQB4Vu2nGLr/Qf6AaowZDK
p/7ljlHbw0OhBR/Ld9gcpaSPnt+JQNgnx2hjvPbTOuKRcMIAqf4jyuAqiqGtBTMbhrWTp2rOmiTu
306m9lMUTNU7sQivkQrbPJ2lmd8x7U7jvZb79ffJfMGdOG89vXQ9+9CRoxqPAzsh5VXH68imCOYC
iuJRum4/lSReSDlnyJ2FM6dtLslDgTVIJJaqFO8nQSL/vFlgy2jZidYboDxmthFXSIMfwnDdf1OD
Jg/KrEBlVS2PhgJSCMx0ajQgedlrk81pm5XMKucyus7EkiZl+2YBHFwW3Dl/Ao2WCTVZ3kRF3u4t
Qs2ce9K5Z5Cl6Y+jDsH4CxPZoTqON4E+7yVIqYRCnI231oodYEFrvp3qSnP7YaOVPX4cKnhICnwu
loZUwCsqxMOnIpJteGLrsIK3BsJn90+6aVElWxgAxFEUNxd/y7OT+GTQxiWLz2t0rlLcMX0MnIL2
Oy8N6JFQeTiPWZwbP3MpJXc+VFnd5hBmGD/NVaz0YDfOUThWuRYudmPdj3MQTpy+B0lq6Ot9J+6i
uGwb5LzBbx1WpcDn3Zt1bD74Th9kQaPFB8NTAMy2uk57HZzBE1ATsu+EjroGrWZalVDJH/vyryWI
ZVJbQZGT1EcFBwITXYgZIvS/WK0ZlepUOKUDUNOb6YkrhPCGU4GLNRDVypTd8Bqwj0t8JotJb6cO
+dp4X+/hAB1Ro728N4DzqG0NEnTKsQJStbZCnwa9W4+8kCDZr0h8N2gtsDk+G/fglvBJLGgnnZAJ
Rfhr8xrEHPXFSVNt81kTlPkG0pjsw9R7k/YU6BUM94guSItjd1v69YbrcNdgCvP+YEJCdOQoLbks
A6DpOJGix+BzIDLrJ2YR6yVHtaReLkbam65ZZROMEPc/cE/iZDt9CxqBLLCWhxYPiE3RGq8ufuyL
NQq1so6IBy0rukRSzDFoZ2PgWokbAW7gyOp2lm0I8uIG0rif/V6sHiwqpE5nMUm7mKsHp8E64nu3
+TNBh7SZY+077Mgikq6r8clHjbA4YdGG5lwI8CxPiacJ1iopuovJTrHojXvzohrVn+3YEd4Hn5Q8
iVuCZgB/5OPvRC4u5b0dUDLLaEEjc75fX9Ce9WiQYhByk2xkmKc3AMRUa9LTU0QbzNVcX5rl8g+x
gLR6s5zHlpG/XYHllNeYlpfW7MoZHUYdM3M7RU5ECKIpYf/qeBMjBrXqlUAUafqO9KdVVAc2aJ/s
ikl3Oafa1n85A2i+aKHyMIrMq1ocyp09+TNcBJ63G53E4IL/azXoSjZi5M6ddnWZnkm1zFxTk6l+
1FApOb+bO/pal2rmf10qGBvUey2rV19wVLcKTgA9n3nSNIyWExvxlAA2Sm10uUCNCYeeNT7PstDQ
SeXQSF2LAHvMrDp6KKH80kpecT28FEstB+0ezfI1Veb+T6lHDLjAqGA1Epbk071AudiEgNnWqF5C
rqdwx/+sfpATceBqS6nuXrbvyD+jTiLZJWJ6M4G9rMsV4+tU0R6R+fz/OF2LG6JZ8VP0PS9SBSEo
n/e42fGhwNX5pfvkJiwwkDFAWz3k43W+veRtmH+Ms/hQdOhuMopF3XIe9TeQL46K8Lf2RDlQMw2T
K8gHKZPdJX+oVWmhdZbY7Od9TfSiCuBe79UtEH8S2V+YqV7aVF487sEf5+cTO4RAU/m8jxaqi61w
GyhE2fx1d4o3Okb7Zh/K1SDVYnZmOYaHHTpH/LqopXgi38oS1DfgghE6sWaa+71uEt/VTI36kWGE
sYtauQs3K1ZSZJVg0dkubXLbyS7LiBtq9/PYRA4yrZuAWsWBA/sKjXdUMpj7PqVJedgNaUNX2VUR
VVwkpDwPBqhVk8Eg15H9Jxkz00+eaALxhwVYjmX89uuPIxaPpmfTyd/c0kpAuI7iAcjfrlrTrBfa
N9wi0+P+dGeswwG067YCJj/fu1KKR9+drLCg94U0YAUtfSR73fx2J0GsFjowVljyJv8+BaSkSEsB
BIw49CrAIlLn8K+T1bDCPDz1mSvxgEVGDZ3t+YRgfBKtj80dPRi1kIyTC6SJ0hA+8nkcAhfqEW7b
DQPpH/bwpV8LXQFN0vD2tItbOJQIO4iGA6nj1BV2tUZOHZ9CBMYAZ3f0J/9ftaZdwq4wmhFHRaIn
Ssp7KduUaJxc8JIpYCKgcwSzVX8yVGZ8aXnuarC8WiwQNhGduem3PEHtjg9FVAec4sCrYNT/guVz
sTtY6HauMszJ3sH+E0BVf3uD47abaxsHZiRlGXrUh8Zev5EaseJwLiU/GW677nVQeQkevcQY/wOh
99ajGNMfUq+iQ0PZ4HF008CJ2R5y20QjTpD1Npv3pYSGGNKuZZh+nzLWFUWu44u9ldeNtPS6VoV7
/AIa0kKESBqKUnSgbjznCRnWha1S1f2MolQsaGNjAnT/S0EL4Rr9YKlwrc871TGw/6zJb6O9LPf/
Nmq5KMTJ4VlAzpFYAdaRqd9qXLDhBKLio6xIuRd9vrKUabM7i4cR8b264riUmoPbKym0/9SZoPv8
WeIsqC3PF7IuZvBAXWo453LkSkveysOxDE7Cl4FAtsHweJtR1i8O407E5tnQREM7ozTCkdUxGO5R
l0eC6QOLddoMu+BNN16idqe8yi1DkmsFr/oFpmzfGE0tyVHtj3MtKGj13FPMV0USpF8R3jPxbkkC
gHeVaYtCfaVrR3Jr/5wxakT6KDMaesjN26cuTYWESAIzky9soMiHdg21c+H8hCCbbcGULtsxTcNC
FO387fQKu+tUzZZfyaRMd8nUJQbGGCGCxZs4XoU931gXcUnszjJqMUwziaablBl9WtpWfdhv0nsC
LiszNvpevDqYkWF6wbvSo4G0xJCT6RAmcU80m+SxIYojhgzfsbdAPQusxrXH1fMkSgzzAp1YocQz
APGnBX41kJ4rvajMAzoTVYpPnQguUtA1M7RlNdLm+qGV9hnciOXaCmCuQuE2P3uTQIvyK6L4e7Ya
snd6FAgpYZQOAdc3rLBEow1l7rMmG8JTwI1ehBxHdDllG/9+QifwtuwSoALUTSHsMmIjpZ9Tj5C+
/qb9u+Qo1XCDgTI0I8lHd6lThKdDByiJXUHQw47JIUGyhZewW6w+K5caf9olKi6QTt+mHHBzOK6o
hajITutE/2VdEJ2qOq0vCSz1lVhg+1FAf2wUpzGimuPuGhQIdMzCMTi1bgKDG2ttYIf1hg5yc/I0
d1vmupi+7/aIpdYgAwJbGfvC1qF2ZkpG0EbGff57xOaRoZYdmo4ugzDrLQYb3Dd86H6kLNNxhE2B
GDxM/k0PeQS05oraaN5jdlpx7kXKnAyhQluFFUnpmarU1pbIDA7h7m3+Fdt5xBsJq5uxRqOQPwhu
PzNnj/3ZJPK1OyOae1kAskIxclHMaa2YJ/r62GpFCDemVvHQPZC0Y+UngTD4cPw8GQjf9Y4HEo6S
F2kIlde1hT7f4qjHvThMBXGtNdvGDdNS1wKO8R2SRQZ/GOfh4ZPK6WGrGDWLNyGANG9CZdPX0gMf
kbNcECE296q1FCX/gU0PZXcT1RHZHTESkKgBXYHUOu2uIhAA/sty0Zhr+sHC+fNJGRBBzCPNQvfj
zETlznf3nGdWhEmad8Wp10giKXWFEe8+Xc+3JqlQxd1adh3GTqpNwtTBnGh2N9xI3NmsgvEz+WNO
8QK4h7aoCtEXfiD5GBk6naf1/nT9cpWDDvuL6+UY5szTnxNAxhYslrQe8h3vh+Om5GULFVpZFu66
u07/46KPXE/z5DqLlTE5LJJdxdNHiOLTC8lH/re5KwKsaLMiac9xPnV9gDuOU8eAaO5A8m/jBGyj
2xJpaIIDY05WzkxAZE1STeP+EKV05p39WZyxFdmR6QV72UZZkfjdSxDE//wAPZ0Fh3pMp8Z/69gM
sByyLYI0EJM9cM1EMGzQjdihHtbRbtVF9CDZfNWHEpqJXYg9IImnE4S1tvX/shU0HJcaVlg/H1OA
slMuf/GrRJeJ9+F2497IQxW6BjCYY9C3+9b84yp8bEWU8EG+iEHCIrRNrwdBU9KXhylZ1bhyglj/
nEFQU/FhirQe+wbz1u74y1e5oGnleleep0s5cP687mH4MGNeEaqrkACCpc7LSro5vde4haEPmmjA
tKzaNrbso8tnw6M2OTtQz1OkcqbpqQAiDk9YZMSYvW5QqRlDZj9IrRuDxID+aklIPtnNjAxuY/QW
xNiZq7TczVkPNjjLCrvQs2MeFDYtoAvAzumbYjO1yM1gSXrMAbotxEnmH404KaivbCqCjQaJW1y5
DtKTNcK7DMJuOUwO0hLjuo/3zXzRPlQxZsBLcQa4QfCCZr9CL/z0eB+qCxQpl8bpdZcm+e/vlI2v
8OHd1yxtdRKk5COqyr3kJGaiDx5pBetXzPhrRijHkPP0R2+MiU9z0kalxTAmb5pa9R1pWYD9acoD
hSa6WGuMq1Q6OYwpHePiNQblcdlUoIlTmt3dByCLeNhw7HlJemOHHJ9pnuzq0/K+HykYR892m6L6
qcg5Ym1u1QLnT8d/3eWJKVawm+tAe4B3AVh2r0e8/fgPKvnQ1jYPwNgRNDm21YLNPUaTfDEE/xWf
CeDx0ooI+EzWMmV/j9far6nVkKjeW/4rCt0J3ZVhAkiYmPl23a2GPQZARzi+PiXvHvlOv3Zsi16j
s50Ccp/b9qGh987syq3nlvtTABYiqkq0fRZoHPSxG/GAis/VCn4wtjjZgcvzfkhP02qRsF06r9Ca
YUB6AtVMc7riys5lHTxRZICyeWg7m7ES003MxDCsLjmelY34hLtWHZin4ft6KiMSOp5Z4l6b0Ftp
95JamWw8VXx83tZV8qhwNNbFLOamc8aXWjDgDF9ignRvCZ2FLSMqUQk3rNVnMCUDYmG2bToCC+BX
cwVZUTMfaPg9+qdZ2sn2Dz+ffXpYAnnvYpbOf6mPDWmC2Ea2q662KbHdDir+elCuIdIaD+Lw1nbV
y6ChQIaOiGCZNSYVwStkuydtPRGViZS3zeraAabpUHj0K99kNfB1Ie4h/hhSZvk54CR6EFO68sjE
Iytyk9EURTu+DH05PS9FFbpehzbYL69Hgo6BNCD9ZiSZGRDiyxh8HoNoTPjT6ijoMevG8pPa17BS
gHKMPe5YKPG2C0un/g8ReOwpnL7ths5i+IYrMCxTrbglYrfP50gZzrsRxjrGirzWlgWNPX50UuVt
jMmayJ7pFGVZIeIJJs2kCyOL1DU3+wzuW8OOspknEvyCF2rOh2Wl7jUnOyzqmNmLN7VBHp/Rr4dH
WWRMO9SUFcqT71Tz5AT4MxWrxGxZSpmvrBujRe44tUrq5jF29c+ekn2ClQZIlLrKfH21BPMEchO5
uh+cP8YKz2bDpiWx1MiWNqnySBgSvMxLRzDq9SdZSVJW3PyNSHXg7+DM/cMvgbgVWmQSlRTgbkmd
l4GZHe72JWEqaYZNJN+4YlnvGepRxQli0fKN6Osh6GylTI5NjNVAOV/lNOtUweqP83pt6yrMzgNg
VoWwc401yLlz2Wd11Ps5F6Ketq196TiZ0YRyUjzR0xfaHp5CnoH4GTgI1vWOGLThtJhzS2OvTCqE
ycTIbU9MidO1tZ/HUUqhCQAWJdGyQef9FdZCTZK81UXVbOxVH2dT+bsV6f9NRuUadCOtp6YgwLy3
2a7133nI778aj1Ka3LmKsEpklz4/HI6l+VKU/pjH7eQFYeA2l7bEeD5isbKZ34vXPzJEgrLJOMGJ
ajp9UHyIw0ih1juQPyS0CHzYpNm0IleK15VDYexpu+hHhP2vB+FImEuhT3bLI0CaQN1fyC0+LD4/
0PBu5c/UJUGucanlWrpzlB5ZBuvdGSkLbUtpBumFJndE3u04sDwGnlnlE9c+D8H7YmiaaFPyN4zo
zX10dbBs1S0Px7UbSpQUqDI7lKNnasJ7X3hElmC0DQhq9zqxXOPMlolv44l7PZ+IaSlvl3L3rxH+
AsAtYZ7FgJIHKia4+im/Gdf6495FJetpEnCu3/Jr9Vm9GzvTlbsE5juSQZsKJk1NG+veCyAgZDMS
srKEEjAl1lJw2g92k+3ZN18v+aN1b5lz8RxAYAS0npQxIXCQ8sSP5FnPcqMqKvtI6t+7bUMM3Smw
sgdCGSspsD7JBVhgE/33esaRFn6dSEOwhiaj99PAiBlevcfRyBcL5pNX0t7aHT7RbrVtxZjGZyO/
kML/0E+MR930P/hMMUy11tP6xijgbKxG2KXwflyhG7IoQUwCg9eFoqM2IWqPigro4YBF95eT1smR
+u2F9lmzrUewsi3AWkNmh97LNGsRwqsUQ+r7iBvQU9Stf47xTmSiEaeuPNVg+/vpLiQU/fnCr+8v
Vz+oGYBkWyscUBA60nvt++NC+hQO8n3oA91TVm72RjjcWOtnpDx4rhW4Bqt+j78aiBwh7SgsW4Hi
1Zsp/ynP4wb2BaP2pp6Tu9IcAgwNODsG55GNHe29G7RDCr8J6PqsU2+WvSJLkH6SmvOBu85PKKwP
zJYWtgqMAo/bUPCaMJnuNfRaFnoiO2ZSWn5Qr4l5NKfphn+0qUjcJ1YSmWOu5k5yeFVHi6C2OD7X
ixm6FA66etk3VXSbWs+iTYKCr2pGkgZMrB6kslgkRIfsAyh1abDs4RId1KOfd47K/gAmV5JQds1l
mFK4Grf4kAyA3rTc8QoGLwrjON7VrNEFmicksD/4Ezzs0lkzqkwmabQcAl8DmWbc4B5iXRmoroI8
OEUX39KUuh/lP86MNLw2x/NhgejeDG4AoYQnNyd+CXWstyJ2lGVy2TPKKZooJvd/OuxvmLPbpP+Y
zyw6XhwsGbW5G8pIPbWD5bRX0/ji6/oo9F02YI4s8ElEHaUahh/aa6M4q7kqXEajhsvj5rk20soW
tubkkhBrMtjIQV5dcwr9MGavEOaieVzeGwc28Vnttmr2oxorU0IzVe5/fTMhUrouxCUlvZi5jT5d
yIEdJoKk/TLTARgsIewCY11t9vVX/S1HbdU5cPkeCJzB713KaifiCcIJgk4+TUVnxbVZMtVugHf3
gOe4MJv++ZtZk6p98m+vp+kpUBdER19FP/Wfco/ArfaQn5KtUpNx/cDsB3ueY2PX4pPQHziK0sSa
D4SGSlN782L0I7X5YoEQkfGIqCgKImtelZEYn0bA/5+knMLhzab02Mqe6AoK/VQKyOJP1CbGAxjq
+PxumnLJtT0n0Z2gJ6hpINftjpFioZO8lh1tzKtFwLhYTYXrp185+ocCApXNWSotrxxjQo8YcGa7
LMIoR1/oMez/LSAsrquD2eFOIsA6gn/9/uewes0WQpRHyfSdYYaKVl76fgNharzA9jfD2bgcm9u0
cnvgKfzUekMK9KUPV9At4Tc7itct59LZl7vcdZhkXd+yUjU2LdhRnyKJ8VyBSRT+XdozU4FME7zw
2q+r9FXZ7vdbrsAOdfwtcW2KInG+DVFonb/1ELXfuh+/iAa3FUjbJH4XIVW1DaQn5MMfAQEswoAo
d3KR2QhX5rJmzP9T7AWziG1n0Uju1P3MgzRlMCT8VBfWqSTTzE3Q19Liiklo27O4gSuBXX+8qCeY
s9GHI5RmWU2Www4hYxPcPGHQ1UBr6r+OZdPiCidmlcAeJIARVTofa2KALVakqYd6j/dkLeprVOy9
WLPvAsal4exB1rv2hYYYHP8o/gzTH41Ub1p3dMJckqaJ3hOsnEpZJyO6ypbxH0zZq8y/Awg64zQa
xI70LCZbg5EXzXtHU2B6Ovo1ZuHbRrpRMI1iCUWjIdfo0WCp5lAf2hsPxrlq6OBPk7IryON2GVDJ
h0rj72w3mPLY01GwU+2t7ssLMG0urL0kHcTRFFfSB55iqARtMPerUAFYTVpYjjcTEHWogflEG3pl
JKI/0XE49HXYf6fd7ZKbI+kwDgs6UjxkiJ0VJp90ZyljGFTcQ/xkGneIh7BfRWxzUlrYAKAGfxFo
KdFt3249tgj3q8lwI9XxjPLmictNh+Zfi1wq2IOuJ1LKojU1TTwc8FfxMViUIagibUqvE7whOy31
+kftpHUcbjd6VNAxWVAlPhHNYFYiG2JbxOyaNlDYN7vgCXGEDdIEWBLB11u3qPfDCyrIqqYmc6Ng
dknbDbivvdFFYLu5oj09ejSGxMhJyOwsOOAesniUB2OZd6of0ENyeA0s+Ac7Pu2HxaG/T+uymW2u
lUhmuPoDdM1ZWRtUmfyIntgSQUipcioDFvza9jKdqLFpxVhxqPIiYNWQse+43/xRzPIVllQvkUE4
9a0jiS0/xNEy1FBu/r8iFyXIsnGTIFgWBA8vy6iwtrePgz3hZzcI5/Mhmivc0D9Yk9UXN0KKcIuK
0iMgQeScMzXaOhxaLd+yr05zMHh/jFpgXUzlJ+TeKmy+u4mocQ7m3x2sl5RVnC4VRnXIA6+YZ7ws
wG9/54tWZ1ZUxeW0basarJR5P+B9NrSJH5Jm+NELKbvFwOoGgvLcoHln7dcdnQTjZ2qSzXHZmnhM
04CKOk7O9HuAY3ySCYbcogZ5D4+8fXvoYbQ46QFcFtasRG+GOp5ChDq40+l641OWQDOe2PmdUkrN
JNSp6pk8A4xy4ULSSUqFDeHay967OP2BxTBKemwpNPGJWWOdmh+Tj/sFp53t/sV7rHaP55NcIP6C
D3WEe+K2UVoL8aj8Mte1X/IW6t2T0rk8TzK18GVOoFj+Py7JnHitOyDn2qb+8bYeE59xuaTlLnNp
FeVlF0fPfEjisePsjcqG8luIoljcy2JdI2rfrqxE6ImeYXQUBQPCH6JaQk1Zr5xXm6pB+uXR5ghx
O743DgGxDL+Fcrlc6Kfc8chSS0Qbq1BTHk/V8mfoVHVca/rdmwSJI1GrxwFgzlUx/VEIMhTGirBQ
PVRS0PyZ5Yhfv2/RT3dEI2aHgPeh4Osss6OfyTBR0n2ABOQYy6f2ay2k2+N6PUaZGPliJznyAl+v
SfQikdhvF2ymjmKne0i9K5hfJpfpYECV3d53I/tyksAvFYheK1V9GVoaJXPEjzMMSqT/KnDxJU2n
KTcfaO3MCw7dcm7puMrxFm0kBaJzgKGdr4yxBPNoUAmMYmBVw5gBGO1GPS+1tynBJhcZK6uvElUi
KYTK3qSdaWqcgVe2AgThvGbrH55Xp6TuhDKt6SYBtniU03iSSHocRzK5Ai5UoqFgTsVvN/VbmCPK
v3IQOMYRpt/K9tu4005lqUIvrz9Rr0E9WOOirIQwSljxV7S0l9d+MBgPWgYUdQmM6xEetMUzu9Si
woDb5mzGofvI5icXk6Umvdq2i3//hU/r2TXALtmaMbaPDW9dAUECMMtX5OSycQ6w1lfXoqPHR3OC
0pucci0gGpA8YCu7Xsip70XAR1QzB17YJ/QlYf7QZWWNy1BjT11SVWCR5rS8QQVu3GmF4stvITxn
BqLhN0r9VP81ZEreAwo8qN2rHF4+6qnb3bXvydvOZBPLoBmn9/jx3x1oWJCCoD/KfhqVoji1hQUq
YIB1r9XM+9g64gI+dpCmLwui5TtJjUhx04l5CmqDlkgMWNINXe5VcMwdz7NMgjT53FdLQDDWyno+
+eYDwWQE76ZzIuXuSnvTP5p6/XVaoh/+7vDwcnUjmSCy6/5PxohblSOkrzh/gVJwk447Jol7Mehy
OtPYpqY+oPOllAUdMVicGVwH1aDyP7UaBRMAtRwjVQB/4MTvmQCFwhG1oDlynfxggmZ4EWvhzTQI
X7DquDzQsBcuyFsV37u/g7ovXoaGEybEUsFxB8YV5M91lnsQWgUgwvsTmDIj7QzsQwJxv4MPJNgX
nDqeGsIF+OdnptOY4KrHBxNj3R/tHpeqvJuVAUHKNG9Nrzis1cljffieTetUr4iH3P+6SyFckBGh
qr8pkKfF+mgk5VFIg4Afe1dn14E1MQ/M1NYqSoOcnuP10BpA9iOQXsYfkDrtIKc6vkEaozkplx7r
iKvjxyPV41obP+KBIXCEncU2PfFm6GbnYQO8EvS7bVSwPOdxgltUIvPnrBxSMVeCFM6CzmOBz+Xr
xnuv7oGbkXGftLdj5ygYEjyvZucpzjakcG/LniPzY2ArfThS7osIGnUxcJzVfQsolShb73DpCcpg
bmPVwXPqFeSg/KrydI7myZqkzYVwxPmyZj7RPbmcPORGPTAB4MoWXzMFEuXoEJT4O689PcnQXgm7
uu2pIPYT2ibKfS/0JvuO98UR7lSg8uGPk8abHNMG5jdugEI6VWtFm9I7JUOZMFSOaZ0uoo8y0CPZ
B+NStfhAGLbZb2CUamJd3Dg2/fe0fUNxoFd+jcbOvsDkV6tiNJAkVucvJJPcg5Sbx5AGH0e+/eZC
eKyVsmRLzhVDHP46VNHDGqO6lsCSmwrro8lvMy6FHNN74Yrf3g1AHUYnl7gNOW1lKUM9H71Vsk5C
B8Rsywl777KTBMKR5y87IKPEpJJGTYJkWXIPZ2QBN8djRCC/1Avt0CGl2guG+P0piaqVOCi5+ro4
wZ1P/STKsyXwe3k0vpWs1giIWm/GDh5Fx0fZUMsdLjgM3IT6wNmVNLN9qsy91+ExnW+YEP/1a/p6
mGK8jX77wygglWDkmFXX4pD04J1+AEj9w5UOaIMveKn4cfoF7svZ+/Jz75XCTiZzewI7MKsngW+q
YVmKzav9NlvTJgyemPPvVJjCoZKHoVtlD39V005i1i/UOBs9paUjm3IBA9qmc5tm1PXGAyWfIGAu
xSIM3PKQtalIlyfADzWvOywwwCAkDYgWW3imYPKBU2U2N5/vnSGgX1z8uFDu35ObE7NoSo0to5KF
AUSmYAuucgjXS/GEZFpTlH7TwobDy6y9Yq7dco4fBwX8Q/dEotMNjHUnbl6zEIruWSnnMDboZZNx
FV9GXbh1ED+1F4kg3UE4NwoJEYkfDW1pOIIsocs348cqWfPZMId1PIJLixTxZOM9FBKZo9YNDakA
518p/uVLeHiOuGvg8oQ7SN0zO+/BJFik07hAHnSbVsqmh+503e0eF+qSIwmMXRxs3QBOb8mfGQZ2
KVolEwy7ty4j9pzYAFvKKqOQKHpJDmR9uTLNSZcsBk875cyVvbNGTRYGt0NuPeXPP9uT+NdJwa2A
fiuI9J5xOpXWSWGjbpP5ReDw+cJp/+g1OEMG5jwLtg9nQ1lHf/krXVnrX1gYdSPAk5VBbPRr4iop
IXe9l6STeBUjGxF2ULLFf9pn/LB/uuC/kNvGgGOj8IdUCnoGnCVdBzJMov/HiXsOIU8RGvGcR2R1
e70lC08ZZodNJ5x3n/pMSuRI3VN/TGa2tGPHxNFAEGrdgX0faDruJZ5U1atxLmYDMISgvjAW1RW+
4Am5Ckua7t38L46jbj99jGXe7yAZUZ/DN3rFWZ7a/IrFlq/UeCfwjVq8DxQguOBpBRmJi9NZT7UW
q7Q42ycp7/AJsuWBJyLZUPDmVH9V6jjwLhPA+enzAVJLcpyFskZOiVsRZrXoe/0PgSMghHsOoCY3
n0n19Kso315RPrlcyEZYzwuAkV2sCQ41zqTE9Fumi4X4WtqxEMDoF9sMcRrBwcfLVvOI2ne2ytT4
V5d81hWTZjR3agMzKGOjWfgLageKyZno7ZYOtCyIw93iPpb1PumsPu1eMfOKIFlG+nAV/x91TGrv
WeAxRcCU/Umk4gVjsY7MZIM6ugfo9FlfwVjpDN0d8nLtBGpBXlitNUx0H8M0nP8mauVLVqxsnchk
H39OWzg4vsUZE092PZKleP8oliiMLkMJFlCQ8wfuadGcZQxqKqVecgvWEVXV6skflGC4COy1D+oN
QGV/K3jImI3RuhLfzUlE/UoEqa54VRmeyYZEtLgexog3w9DnXqE+wg89kllGfdHxcF2R/euwKTmu
Lj1/Fgc+GKX+KM4Ev+09sATvLiAlJg3lA8QEeFWAOblMMfBviIrZe5ST2Np0dkDbI8lCyeWYd8Y+
sXLXLawqjsrUqn8BeNFABIrzvVudbMODmM9LlRB9vO7PBv/vqdVEnmx/D5cfc/uC7eR9IskdLM1v
tjqeMpEtwdawbOwG/0RikBKq7/Hkzfs0g3q7jz/KgbHOjHq0RpT5khlIu63gMQJG5+okHTjK3KI1
6ebZl6aEwpe+O5O+9uYAkPdpdha8Z8kpLhw9MFcpxVU5sEJpZ1ovYwXCSZQPUyT+AYS0o90ZpSs0
KS65ejlW3MNc3nIPN6AEniHglrKeuW5H4nstaD3aGdIwYgJNoVqopLgKtJiH+CTi1MuldRWyYfqR
3ntG/ziNdfDbjRSSRdzLQrmW7e1Arjt6gNahhdekueP4/V2tDWYLhHawu3QiJxfMDRsD/O/4bx6O
95nUEMQCR97GcfIJ6Y3eJjDZehYSsZ8btoXYGZZX+Tzh6hzjVoEp8ElAa//2czM8GosO3lq8+/1R
tcIAJYtG6aRfYDSR1zibWx/4a9oUGdRE1rmnjYgv2516eQhFjnxwxlcHrElMhcYrNXaNOGF1TYZG
BOwf5xwTc435p6LBkFQPclw4UJoyJjwoAnD0GZBnQcUhmlUh6ZOkdKfm+kIX7+kq6IFxVbQRuLKU
s5k0K36SqTop2vXTx0km34+3N9Nj0qLGlWT684vhmwqcsL9E3xNPuIliiCR7+1EbOv763SuJ0tsI
fY0Z23IZqdx8reHzlLBAV/zJ35ZEI6GyopK0+8rKNVvCbJPcfY+Jhly2TwZPMZCqZdGrwE/QQ4Gd
XW0P3pOI3kG+OPI0tEKZVCUjHOxZeIzh4l63oMVXIhQ1X8kVvxKBvgRyfRo0cFgOH0wjcZBj3+dJ
t3KDtDV/eCWeMCVrSR7/EKKKTbIwG+rNV3rQjKMLjVtMUYk2++Vm3g4+/EL1CkCEfD3hzsAuiDCl
t5TptyAqybvTFED/NN/awO1n1q0XHy5LgCBtRC65Y3+YxmfCzQngQ51Oj3zGju68D6vPKn1Q65Bd
5S5Wndo8zGfxNAFa0nlTnCCcaGo3sLa9VBc03j47zXbVCnRgPNiAg7hqNdrQrPN5zvrUPHK09dqA
Cy00rqJl9UopIeXup/DJgKFsuotO3x6mr1aNHk0/0Z2PKP5rpu/085BXl5hynkqGbdAG8YJoRTI8
JIyabRlGtL+b0vrik96Vym2HwFoewGa5SQmEp0BO+seabBSygdML8ATZ1d3B5bN5kaL6cukKnDlM
PRdLf4spr3NR6CSBF3pxUBBnhXOP0svhZXct9jh05BuYlLRHB1DvYF1dzY2gKj4KzJYm9J70yuFJ
S+mNOrNqnDN1wl1rRrhABTwbLlC5gw32BysqhTh0t6zRUdxuAYkzypG+oOOL2Tvj58eM1uHbmciA
xCz8V/jad+5WbGsUp8xN189/CukbUDDF0dnYkStyYPGDHzBvYc2nyE1rs+sKm9vsmzb3WtzYCHU+
aJAT2DPkD9U7ILL8wDLmfSSHbPZH8KDrWrYqPLvR9/xdn6Lj9eG0DCRVwHQmuLCmhplPdo3P2P8/
CY2fV/fj8ie/Zj5+bOf6wG/Tg6kZu6/eGXjj5FKcOgjr5mNiYYZeCbQz2az9Tv2p17OukLX59QxD
vmp5QBSuHP4TbFGeNcFj2B712Sj8vYmgptVfPssQBEJkPlP+XwEhs5NOWNfCZE9wgLW4M5pPnctR
YkNpQ0hnvJ+jswUb1dCjbL5EgmvZsOR0wAVgb1ll3ermfM6VACA4pmzwO4abUINF+s/osQHgUuSe
elPM1Gixticn5mu5QNoTJsPfCePoK4g2JsU1Bua4Fo0ViDIq5Vp3sKTYHAaRKsuwHb9cTzQWchYY
G7fY0p+yYfFlr5ynRXjbctmOCq+YH2Ka69VH4o3xhxbwoM8ajkaehdrQu72S9sET0ixwBpAp1ytd
sTU360Nf8+gSt0P0MmLk9c25Xn3PpRhsM3d0o5GWvlmcA3GuZSigS6NfzL49UcerwL/F8aqAcwj+
dweJEb8tBTJkxAtBlslnGXybesTbaod6/y4qQLed1dBxTLkTyGGNRXmNRDs5BwD4q/hAH41Yj1+I
JNufOmhCmUPL6ctKwwolNXM+/o53/5+AE1lHT5ZgCra3qKRlobX5xOe1m4NCXYMGKb1aYB+9H79Y
maRDoAGAJ9Llsiv8BESzJNjEUG0odGBrlxTvXEHlKOBA8OV/biUH64/VjIEIWhAYM+0GWGhTmd0Z
+TuEd2ddRxXG9jXkI7A7+XQuAPwnOrUelwcFl05KdcrU1QDeOlHZBwnpI3GXtijHxUyM+8UXzpnA
IxFOoVjlqvqnovUomPNbZrERgAT2mzLS+09TdNamBQ9F2iMpGtKxfO/unPjF1BSo5ZzZ+7xu78bT
0u1AQ3tYifODI+T8HasYJ7hutHHOZcBtOSGYZqPRAg9NPH8DrRcEfKrPOjnW1Oek9pu2KBZ7520Y
P8vGN+rgTTkrFE8eRWRNxCFgb2Ta3o9j3Q3Myc9mFbRNO56KL8U1Zyb+UHv2Cbzm7dghVWiyNuU1
zTmTs+Q6xpHgUk2zrvXEUfit7WF5EqotRH4oI4pZeI9RUcKvBRagjS6iLjs6eVqgUkiGqE8YqsRB
xkjCaOEd/ZHPTaRGSaGyvPAXCDVF+UYgtdEZAZxtfslPuiDU2gYwe2hzT1FAw4SOdQVdG/SHz4kK
Pp/lFSr+tjk1nRchK3z/dMWOXpACLu18JgMjFLT3ob+XBd8D+nXebW6uhiBFXVGku4XzdLBJnxoz
XrFzNNc36SmGs92FibqGtBLXdm/0wk1333XDMnch0RJW+8zYyxkrCEmbTpxxVEGI7eTmbYo4a781
+MuEeA5wIUgPkSTrK1uNvefXTTuUP7rLyHdTLmWuldLTZxBZd22Ec+EXtjrH7l6tGnyu8b2Txmjv
wSUevCcZR8Q8YGYyaaDnIM85UByVSeSL7QNYPoXwOqameIzyAVkhocZMlYT4ztL8eyOrvDmcWbUi
YC9E/pdYvagFjit6QxWSuS3RAdQypBXoq07ZJRtFm3smO6RDwrdUhKguqSvXatdfP4cVp/QbnPtS
Yvct93iRcQrvS5bWAayLMKUGrV8e71Tu8u5CYqpzQLvqtFfZSGP6ricfFxsttdaml7yyuacGoj2K
BatyW1kXfcRZ3zJbUAbJUoeYKIk5lceuxTG3A0YiaCPRSqwrio2+f3uFmBOLThvh/0FJdWnLzqWP
RxnooPUSLvkXR/AexSE6NW0OVczQPHFd0jR8pruMZzpwASFSTL1DMXL3a0O458DZzQv8V4yBZRTs
/VyRL5o5NIRlcFu3NB1zGCuVbdhoR5fp9Vsue3wlVjpfg9nSY8a5bSBV0zX2qdN/jW7BLQiGB6FR
vZ+y4I8vB1WKVJkGPRwcwQIxcfE6WiX0gs5vVHuSnQz3gX+mav8fY8W7BZlaOb8xa6t8WEzxTqXa
FiB6TbMN5r8ZY4+xzIvAYQaxs4GBGqRzARvx+HdHXEoGUVm6GR11QLHqfajTpBg12znrK67eDQrr
MhhUEjo3Kzolonbv+xMGQ3e/xImyZ+a1CHbes7oC1X447cDDaizIwaoaXG8M2TpqhQ9dAfJ4k/gQ
HCIAlGeZpY1GUqXcU9PBbrtpXY++DkK8V7/YsFhp0s8fEwTzYGa5KFr9lrzaMu0APkUhS+ZfemRu
Luiq/qobHnkyk4wOEaRn2xnllq62OHftLPfhruE+GSswhpnHc+Iu2AsEJ9ZeUcxVn01WSR6a5zCa
F+2cwu/BcO0Sktrd/2+rG6ufuHYVrMvJ8SrmRgCm4Cv8/iW7DXptfhBM0wTCcbVTUoSVaeRkfzzE
UaJmGNsqnlf6516Q87y0l+Vt+jKKsinqydsRAmgs3oLgc8G8mDmQbWC0CUVHeiIk9GTOjWjwyPuk
xEombod3cBdEbSQUwbPhbPFbv2nkft+JVm4A3DWPtjvuko3+2/tGXZn5HlLqLj/zyVvswkWTOo24
tHlr858NNLjHeomx2uWMvykkl034xLVI0e5YlEelDAacHjozzFe4Tjn/AP+a8moFyrdiaws2UnG4
Rf0Hv9/1nLcatXRnMvW0RWda9u4eoCw7BV5NfhdlQSo3ZPLXW5SnrHSWJpgj2feBxJmLjwOIPOzc
ZhZg/P3lGt1Qy+1w/6S16XEsaYcSnF/g/QAmwlXJw8N538bz1p/Qt4IiMW0YK9IU4ZyBzxOyQmZH
ZirVFnSSD85nC322WLFKazQ6hib0PPxO7tczHGrrJffKGTUTl1sFwp53hlQrKoWuAew1wmUQVZon
8yZ2PpgNLmHrM2AQ4jmCKO+lDOAKjPWfTKsZGT9nqtujef4C0rDC4CXA9LABaMbBDQSY4L1/z3BL
/qGu/V11Vh1d/ufTrf3Z+2ClQS21Yvu7CKH1e/jUPGbnWbo/zjTb3oEP6TdPbvYl+Q7F1hMU9W/l
6dojOiBaL1bJy3jEr/9W8v0qeYrTz6L91FqhGJO2W7TiBXB8k4J20e/Vd0h+kKMhZvnrl+2oAsGx
76jPKs1phr551QnXSlNoEv/l2FQn6Y/Xu1E/UhAzJ9Vl9JtIF95gOujROfb/sqQXYKqiYPUVLjNZ
1kNvcrCR0rcBTsXqADvIvH1oSiREzZLOFTvlsv1MMggwWhapzN81LIU+iH6nKZ39hDCKXD9OWEz5
LFyzycxnP14yvSQFUMKG3TQvhSTSjxkj/wvvwQnOpvAnM6CGqaJ8nR5QZsAWhSEAcZ/hxC+1CiiK
upvv5fQGhoLoICwQwEROuXExAGD/Rr2ZhIeQ5E3hkwKIZzbDVNqhy9uW95B5Q+cA63hqLs5cQYtG
I2gUsjJf1JUlGxEot46pU2Ss6eIhI97UzcJcS+pzo+5P2xHxtZ9kHEotAsYeHOYjqc0tr9Uajth7
aPvpMc98CZwhjX82bPlqlmwDg7c0ckzju1DK90CidGQKojKulDK7xyzvAGw0G5js+z0/XC88pNMP
dBslhQvOSuCvuMs16SXShVWrYPx+njSxlydvj2suYMsf7CJ+TH1eJLzdt3d5nzPGMMfLOG3hqf9f
diebkGrqxuwd3RFnxhkmCB8pd61qy/B+NYvYgHXpPkZnm2/L8+N7J4WERJrhcypSQLXAxMHb50sy
P6lZQenmANSB9o7T0AzZB1DP1TlDXB117buJ3akJoZPuPi4cdGTKSRFZ6WBes3Tsa8VV8D/nAhXZ
j+9Dkgjq7Hc0r+4p6lcT116aYQPs2gWVCAUSSPm4Kj54dbdunYhq5ZCW0h377tg68udxzyMqVWFf
qt8xlnB6wQoM2heurpPB+URSJP1yxPstQVJ1CAK6RQF5+7+rKQPPaBOtyDcknxXaiZtKUYQPmhUk
7sITMy8CXkeVH7EF4Ymk+9V8nAfqYGsyBFDABm8qyEZPPyhFYpG2SMrcpOxd1qBlE8x5eVW52BRJ
Qa/iHqD36hSYDEHvpZd235v0Gd5gurWgT2M+UiIKQ8WizvEAmSGvvxZ2gl7jb8CmpA+efHaabTXd
6ZpqKCWWZBd3iXU2rpK3aPNbb5m7rx/MYQkDfi4C2jp8x5x4CwpPl9/oShLlLV7KNutJ3fZzLERW
0NlyV9c5W3kkWnib69DCo9aDR5qBMlPAdXZpYcGMIn5/4SUYpUehAIbz6+Ptu0bmLrvldX/Cl0yv
7iVWBWmYNWnnnAdZn5YeaYsIWjor9Zp7OQJSswe4xtF1pjWgxIHEwd/5Aa1eDnn3IYIrQcx/AZ51
ozDfT+lMwe7i3QAn5rQHVnGgwUoH4BG7zwf1ikdg4CRI6iXrpBo6ysokFgY6ZzKhsfX4SI0WiKdk
PHWrnHlMX4SM55SeSZd6O+k2KosrwIZXDiXRqfXTZcuUdmHKCiiOmF5M2CG5QFE4+Wjtg7wNqF+Y
E6TdbNsmiMiidfuurrD9L5GCVuxrnbf98K34m8cFabeNmJI322fq2wT5U4bQ2h0marhv3cacI5xl
ME5USO4yWIhLQwkvT+aHQ/Tbf1DpaSk63onkTId9bZYJqwxky/RwMj4jYsVArRdH7CYPVXzx7Rel
Q2NCqWPQ4a2WeFqCqTyqc4PIjt28Dj7TAZUkouFtZt24m5s8QtcZTbE7/6xXNlOAyR7WiYMxLHVz
hyGVxIHNs+OmIde68AMifmiuCp28YmBO0UAyclf8uG89p4vXhWVROMAtTocHBE1WtosMtYJ52KMf
949azXfhE5qySwYwOBlcnnPLGsL8ixREO+QdtOtFMrHzSeZOppNOSHPJI+G3knPBd1ijKRU47gt1
0sIm6SQOqiUPJRx0I4NcbiOwzIpRcc8DrnXy90qep1lWbQplVQXC8CKcgyt3f+NIVSX9+Wyjrl0I
mnTc0Gfv5WfhBGtD0jrYxanOru1w7ppFYQQxr+0q7SQu2zovFxeo7vtFYSWuK3VOpsjmuMXrYJS/
kcmebBS9EzPdS7FMM4i4C4acf2Rg40cCScvT/nnj/5Sd5jIbvx0KHHmxws216eWfpTgGQlph9bIs
PFqeO52QraKpVyhPDkWBs7Ehje2yP1G1HMv2P1K/l2IyG0oNAaS2QjmSSkxnXRKfgxwGwfnJ16bu
bL8MlQPUXkaFQ/DRIcSc6IifTABqHunMibhz89VhWQLRt3f4/PHWVW4Rj1d1XMFsWR3Z+SMG/ylc
y8sQxVni1AgpQyPdMitAy873yLtnrD4con6hW+KDaXVkncqYkncBG8Wr6fE8WrL1qvF0jIu7QUvQ
fFicnXoGjQ4JH81YDZBnrzh+xhKQIQw9W/+w05OgtA1mqg6sYOeeKmhGMiavtrQ/vItFLR/cNFyK
WjrNYBDlbsjJQV3EmTB/x2/V/1DzX9+AozwDh5Dx4PxgbkQgKybjZWPLGAwR2FQy70Qc1KbvuVr6
xfpgVIjy4Pidvl025JjYwn4qLavyrAee72b5AIACdFoFK8CFRvPbDZ6g1x3293VUG9IR3POjqroK
G1Uuvmoxy6pc4X1X/yor9YEaVnAa2+dL5l0xfhWTnSGQmC8fk2PMt4dIcskGYNq0bImoAhPY31St
SNKjWLCW1668iW/ikPHSSiAcSbq07O8bhHVVseeE6h8NbuBnanBguXIPk3QEH6JcsisPrq9nVYm/
JsSSYf+Ms/1JKWZ6njSiwcQ7dd0twLTKzatRv1QRsTSbaCC2XKxchuBVUTindRQkQmwfv1Y4K4BP
D98UTakphO0TeMl3OTfZWFYqQxxu1lxgs/GcsQPimJRUuJduonfsQI9tghNh8vrxrkRZzBvTyoko
+CtLERm1lGJizIRNevOSn9j98EkN9FZ3mCL42ElGOEbm+UHOcditX5XpLpl9dRCJQf0KfzvfEAZk
QlmaiM3qLdD58AGU3txlNWE2Zg4QG9+pgSrwz9BMieKA77vbU27I9GS3+5DDt5m0YwpZ1dt1eysH
y1btQkOmJhewMmoLKCqPnkzAqTqdLZMrTGu9sSaaWrUaxeLKJx6w80UrE/2n1FiBh+KQt3ibztdU
XWnXDkSGr7GidZlFi6tUkqpxV6hDK4mF7blUiWK0pMNwYzVtVeroUOC8lhtXsAdDNkgAwxcguaBK
7qJWScvmcpyQ2i2BKgLSrVdGgb/7rLKMvcdxOGI0QW5o9QaDt191sjFIPBmKDKuiEr8YrdL3W4t/
NHrqPHj2OwOdC5f2Ad/wl00dmX4d8tvEg9vnOUFk3VXC1hxr+yW6R50bd3vV610qGMt4Rd1nRUj0
YII37i444UhUaf3FRb/KzyjW9soegkA8mQRZZoYjaR//fFjb+lvJJCwmCuCBRErMTlL/KfTBRn/+
3ZMkMLyVPSwz08WqDIzwyC4h9Lg9Jc1MCfO8Toqxmvzq0enXTU/P/vG7MKwCQTchpKfxHzlHqcz+
V6JTlnF62HBVA5ynv4rA7UiuK5lzkdK5VqqyG/VnijXVDUg3TO//PUhwLmGDswmctTCe6Pkh9rWD
rrqFzcKvPS/KxLxfs8pmcdPS4O/3A8blNTDVRCbJuSWZ3RzBTsdY8HA4dUiKaiiALDunh3XA9QKF
oBUlVcvLX5hbJ4vWOYmNXZPlk94kR/uKXoUaysfKcKIi+8QiNgEEPRU0CD3rfHYzEwR0Q1LOw/r0
7fgBUyIZx7sgIp3PMP0ezmQSlAoRzj0wmWiPPfVRxqDMxJo+YUrAEQ8HDzQ311A8/4OAuxVcXUat
KyTtpxkTuOB7rQYMNFe/QVkkqk258a5Do6XlJ2Yc0hpp/g9aZhG0YxFsvjlkEX4vYBcDDGCu9TZX
+qkiBjTFihkjhzMQKsfNzd+hP15Y6oQ4ZqTk0dIX0mmnAipPd62XsgWJhQOX851UnsDNgyQYb/SC
dperobUWh7khojUMHVa8X8golzXUdI8hWA5ssvbDWFaWuRRnFFHY8JXj7QNUKJOVrOQjC+yK9uNx
uJbJSr57ATBYnsEodwtLOTl9tk6goA3jjJ661hA9OcDAPnGF2hmT3IORZO0tCPVKnlprxJAH3oSa
OEhLny7opo4m2oiCUjSausOHK9Io07EiLXLGJ6GCWx33fWbWdJ6dM/HvVlgW1OxGkVSVSlKSnlJV
UOTJ5hHhTyZ2MmAIGBSvI7fmI/uBamIqGHXXZZ/p9wUhbXlXBtpwb4O6Z3w7zvnSRBGAWI9dbvIO
xmjrihEuzJm0bsOdh6Px+HrlSajqkoWr8psq5nkRxYXAaRdHm1D4Hi+9SdzeVOu4ET1Ot8v+ILh8
Xn/2ZjvvNpdWICksl6xM9+w4Vi+A497G0nsJyiKk7OPwB1yVuaFxlJj7S5MFA8vvXy/rwWc15iC6
P6IPOduLKKrkmchvEM+3ccA0a8x+eLDVDqblHaVncMCdVzLCvbNqPJS6f6EjRQ2kf2/cZxnrGeNI
/BDZ9WS4Sq4WUJIcKdw/fbC10M+DgzcP8mXLKiNm1BhEDCApKSBHzJtUeQk/cjLS1oWQ//v30LCp
ejvuvli1FgDvj00qyhyqAZp4586qZmQSkUm9DQyJyYn6Ns5fmn3lnOV3A3B8SiPKdiFr13Smk8ZD
Qa6+5REgBBC+hFULmlXr/iEGrIVpkMtPRZg5lybOTGMS/ukq12z0pdZ72mrhpojfaH5bzrIxFzni
WeSVYEoUlwXodrx1H42Q/OfSGmdcDyozXVXIJIK10aP3fyjjt+hiBvUwgSZNYq2ReqF9E48o8oLt
KDHh24IrCy1Rrt9P3xmVTS0H1Pzm74OCKoVjX5tRn/lOQhi+e02E7+hxM91uFZbiYTnm3oySXJve
lfx6hBD1D3tT8LJ0P1mwKUfzDsLdSWb13T+WVj5JF2ApENaah/x00hIO+uNI5P0/dGqPMeId65V1
0xngGFJQ+cGNGoLZ3X5c0oFeTfinaYXfTJUpIwCpMCb225lq4A56Ug6//VmX/wKQy0YH1UtmdEVk
RDQ2Zm74+2qd5WEh668Fz6A15b/Xg0jm9GInZ6Y5mjQIs3ekNAGb41jiUxDznVtRNGI6VlHRmEjO
EulZkGJZm/LpCy7ihN19P/vC4+Ky8XIgsq7nSs80vzwHkKR0j/kfe4OIepl9XD6L0Ay88krRrddw
AJjOyADiinYa90a0ysSI+1galY+NJKDPudV+zZBWNF4ChjP5uqvSvqB/CuPDjHveLGb7+sGNIZVJ
uP35Lxc9wCwBCxooesTd1zqBZH/IqtYprNS/c+yJjHz01CoXdn3UxEU+kQIzUTv83BQDZYmnwFdn
98EKBKrHeHEuOuKt7oneINeMROapcjJW03T8y4/mIt1ikem8wyi1T1Nl3AwPj/AjE0QOhm89TluX
0+9WTwZUkvtwB69K0ammWRmDk9fbiIzW+n+lB+Bk/hnVja6HEN1Lsi+Ki8dNG9xqT4SCl4U9RVBu
Bxnh2VR+qrBZIg1+uc/pYToqpZo9pvGLE4dwljkP6O1rzVC1ffrW3gc1rSxsxpTbzBYGzQpFQKkP
Ef2vriijwPqdimrbHjm2ZNR6uJk2HGFakmRKR2G5VbMhc63ALlUSxBhQfvA2LlR2pfoI2otoETQr
SDsE/lko65hEwpCwR7qEYQT7rwptrhkhJJ3KWwJ5wvHwuHhUEqRYHkCXiF9I4/l78xsz9mWZiPrU
sgbP4Cfe24VICKXFr1auZ35zC5SSSQmKuFtWPwq5NGC52jPzqmw4/hzgN6P3YhpBcpbzXL6c3mJ8
J5Zu/UhKSM8XXwUdMqoy/r/IQizGDb2x0cJuvtV7eGbMvgoGatPTNgCs0cJiCi6QhlAYu3YgJu14
+62hqczqxrcfeXK3JUaPh3GfAg1zlxOt6CugWXvkshnDsX94GYwXEcS2qMqq+gbh6m06bOz7cP7s
8sf2s2BXgD2cUGB+GzSAhbIW7nKxw4tznuMvgzPFoM1voHuTyvMvXntTatGHfPWGNevXZ4YRH/ye
wYrQCBLLZC5l0U4J1tnQL5FYdddEtiGrn+vsCN+UoovQIe38u6Lm1Q8weZw/lcWHgfE7jBReWUyR
pIDQ41jJAY9na8YQ46Cw4u98FvF1ii/H5lxTKcgn4AkeH9Z2n8wU0eNt88fh/DAmq7z+1pLDvqVr
br+YAzJxsjQvIB1zgTSbLNYWMPgdKPyKi3S1XDIJzdnHrQwwx+q3khaDQ8PlK7e3GBX+gMHqWLmD
9CPnDifNB/DybAMfu7Orz+dEFNK8lpcW8IDkjSD2FZt+6kFhkTsBoPOaX8QALa1VPdllIPGDlLDV
f32tTAi7ZkXEZjPe1gstNgdPq3hrH3JF/rW0p1ZsExnmvVtM2H1SWg7Cz0IiW0meBl2dPbya8EZi
8rNyzlZZKUoPG+LkUX5jfU4fF5tGFW+vdX8Jb06GPKa8Mmz9754g5DIQJBN9zBeSGEWm04XaBaWE
ZqNOwQtS7jrRarXod1RjObnfPfelaJLIDqryppXo8hzm7sgdteF+JR6O7hHp0D67TrpEI3cI9y7y
j2xb61/Nrf7c8ayGTC9XeDX4k7tZY0dr6X/9B3emNOXXEI3IVDV7ZiDrZQepnVZ0RmdEuCW6kko3
m+MlGz2wTmOYRIeinTVr+xWE91BJslf6RJTTig6APMo6XwiGDXz57dSHMkEPMDBgDKxfvoeHEnJZ
0pxYcJ2EyjTiEtQ93Y2KPHOc7UIey8mZHX/1S7CbezRmrJTIkVamfwl4L6V3D+S/w4DdLStS+D75
1vb/DvuxeSThbLwHffGWVJ405IV/oqZZpWhBy0mS+aKI7hEx5VVaCv7fCyVqJQpEsvtoV7MFTc95
2zrmuZm7JMOdq+5MGt/OYTZ+UDT3spi6IkVoH0QAzsBQFZKMIm1QOGdImb7KAONkjJQhA/4y549J
StBStHum0W+HZdTgyo9TQtLeHjJjgO4RRtKDzPSoGIcSRNXwlezYZbh0o2scIDG4n4cGjNYt92Ff
3UquskTNvdjuh0I6uypAPDCwDhId6v2ZQKtMftu4aC7pQm/purReAgz0waLm2l2HqsDdBl4Oi+Tc
1VvxWrOu4hGfx3eRkD9/mVRG4WieI9G9gPS2TFvqdTTFPqQ2sdZ0L7qCLg9fjo409esR/rsnzKuu
z08kHn3f/UsYkEAVPI9wieBo4VIZZuhQ01Lt0DIYsvdkqA0ueC2mR+Ua6Qoi6b3Zt0yhDwOHNQfE
x/YHUPuo7yXTmy81tafg0tSQnbjZxKqKZhJPvaMzIROwLMIqvs/op4ShEaOv1yMu/qFbZ1UtEMl9
97M4OQGorHOFbdNEYODrqnR7mnptvhtZcNcGaJWcl5kqw8aJxyia6yV2aNfVbjrpaE7USbNPHvcG
RK7GfBxuP3/oRbImW/c9Jg3MXxVIT/uN0gsHcPHtym6J8gT+UduRn+sB9sLgESfTWoqCHZH0goMN
dsmBgXPo6fPT9bg7cn3icw6uYiICbI8isKOpXwih4ZFxyvktIeYC4bCY11cK7iKNoKTP9957FY77
LEV75slTKI1zKNTRvG/E98Pr614135TvvQbj+RVwyLH/rSaKHTGSYnq3UhAtr5jwUlxv0jcXDSnK
7pdqMhPt5vpxPfQ9DLxcfFMaEWQOelVBDOvPvL2JvRVmNmaN7Epg8VJsu7ZjucRPhcAOYqTrS6O1
E/EWYCGUC/823N1bjqfE1lDIccrx2IhpXEADRF8W7+nuYXVuWmp9mjWSlEW3JY5K8n9mzWMPEa+h
a7rwZWGSBjJQlUG7wyWSVFUD52IRLYMG4ZiBWlJX12YtK8B9O+yH8HoIjtq+KRQDpqwFdlgMtsTY
UjOPBfZytpG6YvwC8oqhGrJUs2rNWaGGpKmwuPrGVkQDA30dRldYPkg6MleIWqNGRhM6E/wx0gD4
56/faUn1GQMqaB2dw1rRDrHgzUfFQMAdE0OdgwO43a16RDLOtDPRHBe2JEnE0EkxYVA2x4NvgqW9
Wkes86Ba4yj/EswiHj2+IFgJKF8LNsFNoRNdh0dYiiHBLpJoqMAP/cx57GZ2Du1M6EmDlMfmtJZY
h8oVIK2I8Lt/YY/4txMGstOUzpAX0FPfM9OiLYi/qFC+R3LIyiMRgY+yNugZ83yxLGDwN/6vY4Zl
/3K+/6i/oDINECpo0DccQK13jWqlbD3BL1Wqk8L6aMgrW7Jyekho0VHj8+9KGLdD9r+TGtCi4Eo7
sJ6UDall1HogMGnN2Vehte0YW9vyQf8uJSplcGsgJ8TJXlbbGkQFBTjV/BtGPrzpsH7y0TlgHvGF
/01sLGrt2lPSy+7hs5i6ye7pRf1qYqIrCJJ//C+rUBE3rlHNerTytygHT0XWvkWgjcAZNeyMhFXg
QiQDkzbAFm9YGblarFdfdycDE3CkK5Lje/6Yxslr8FHjp4nGyqPjFDS7AHYXJcP6AUCQNV5XhTvT
TGOYe11aN1RS1Vq9Xs/XATjZhhHjNttw6V1vlLNrlCBbfczg+DV4ZtmW43HCW2fBG6g0K9Slumuw
Vf7aJBkukgwO/1q5yJmoYiNbxl2RF8JV0xF6Xw8a/X5bQ19LphUj6k9H9wCKJs4Ijvpo1ilyD0pq
dnzZXJ2qw96nhh9nmlQA7S4KT590NEXUZTT6AYhtGoTWfedp6IiS+/NtuOGtWEzKBUxGb176Tz7f
D+J13jzcqv/uFo2eTmDkSYmo8jb6w9s7tOWY6TsXiT9jd0O3L87C0CuRCReNczYAwT2PwyaN4LIr
qJR7mW/WwXeWIGEk7GNzl3/t7wuUGVxvGuOloXMlBnErdCfQ+oapC2FO4fAwEQwQ4BWEu6nBgvlX
EWN31gJPTsN4XTZX2jTnC+8Df99iHk8BqmS56SXvAXIwYjvxhGBh9ujv4RUwp8hABH1tkH2OgWzj
DP5fEtiH3ZiL1lI5NJwN0VEbL5+L6Kc+tsruO8PAY/8DSaRuN7P2JO9VIppLrL1Ic/crkF8Km46/
f3tcwDdPnqy9DVSBubeY3tqGH4ERhbkCfau1ghcGGf3n7l65lEhI7afX6ytGB1y4MSSd8Ql3Y6hg
FuZtNlsDh3ULbAHbImJLJT6D7OtsKKHcd0vTqFc69VqMmCov96jjp5a5dPztM3JWN86B/pROHF+V
UYW7bx6Qb2O1OmZeWz8AZBi9ZJDclfDeBIxzztS8gtGnizwVt7bp2ZMNlf4DzHg3A+pTF7jRAUtR
UpmpuBUiaDb+jUCmu+/HBxb5OMZ8s+EIRFZ0icFgiA0+S7IJVFXAWh9lYf4HxL8nhI2+gE7Mhg00
Kph4PLmjHuHAUFQsV+dASI2nVo9F5fd60ZQsBYl0PjF62EDH3VRzk+IEDvcVnxrUP17YHP1FiKxo
kzCqR+UfdJJ4una3get/ny1Kf8OHED70tFzfa+5S1+N/XyPS89LFCSf0/YdZ+Lxk+jMK1EolZEu6
+H9mQFmYy3KfQuS5TWp9FtxbK+GSbZtWt29kRXMz5NOOb7nWdWZlXHw1XXKV7jCTcEvIK3HaAH5x
2NVDxezjaviFqKUcPMKCg89cVD+ssEhd367rD37JL75a1gwIizOX1FnBSqG2fT7LnzVCSC05GW7R
QcyP49fzvPYcuh8IQsy3KAT4gzPDan77/Ou5M74yD1QEET5AJJ6CuDor1c171HfU4qNl7Q+SHoPK
M1WRV699TysA5IiG/maN4aHHqY4Exs+Hkfa5MQZXDhN5S4pHSiYtgcEMpaDUqIfjNPL1L/KOpRyv
d8kP8uTWNe9L/YSOAf8ktgeMXfq7Ww+xba0p1AA+gTNXO4WTVUY0i0dR3w9fCsO/stn867d/4+Eu
cIDUQCxG40UF9vtw09MLmZ7+KoFPnp2wDcc0fHXg7YmqzjS3Y67Lpz8+JoKeF+ACgLIy1zDpmymG
WSvJDPa+nP6BQOZJmeZBB7jAK/x1u6NJmDxgTvMy2+LuZrbdDyk+w/5Cld4AcGHkZxXVHNrk+pkL
L+ygzF33gpxTec+YzAMPxUkkOvt2ThXDH6OeC3afpPtJ/2sWL9ZMR5nDaeP2qptjPtjUciVYjcT6
GJ7/YdnjU/J0XFVdGXRM56heT/Eosolql9rMbrAYr5H9m7ukvYLQJ19XsyiWRBHsFFlb4f9kEo5B
j7bw68a5Gu0Dq4nLOqowCbF9drqaDhBPn30uLCzL35dB/HV0LctYyj0f89pS6InrjZHkqvALc7po
Hknmp0ug1GbPUoOX5fLE0rityn9wjq5BABuWzpmzhcMvGw7uaUdPymC4sJpkTUQFbwkcxnvDawfY
Cw63d6stiixNRt63I2H1K/XRGS+hpQZh8nnxxTYhWtHAlSnrVC/sO4RJE/ixS9EG9qrjmL01bBLy
XhWogH3ULP/Asc/uryRnXvdqOSSpuf28Kb73LgpVok/ai1jLRLPUboLtNMDsSJLpQhx8mrlmFOYM
hUbf3So4lkzGiLZc8rNvCIA4O10uPWZMmRDDvkilJdCnTg5AVu0MTjLvXGwW6MOv21RIB2HhaZ7j
sGWGbAjJk8VzhlF6gokkmE4AoNKHoEeM/f7BTqLx5G+nM9URwfgFXai4nvs2AcMvQ5GmqV7CUZ9S
4lt73gD3MdU+QuD/SFrDWi3Agu0Q11YfumICRFILNfTuPv2vh/aLNivBYZMSZ950u8sZEQxHsOkc
+XPPLYFkQ+Q08d6cXSd10cXcn6c6uXO+jxPxUCgsqFCa8BJHhhVdBc4CvNFxtdB/R5UHNBRSzmxl
YKUvDmB/FrWxSgNP0aHGzs4NVdItG+qpS/M5/8mt8VNSHIwFkNPZjJY/pcI/mbSxu4bCZWDNSFxh
2uzooBUoQC50ZnUfhNZwBMnnpV6rGDsDsubZ0ScodS1Y1sDEe6g50DOTXPNajbyGJNHQ8TYLxcWv
UJJcsUiwIu/dEk+lxmOoumv9p3AjwuG696ticpF4W8XooO1mEHAAQyxA0Y9TED6VSlayNgFRrACk
EteHoBaEqQYmNxMUMTZ3b3Zg0J6pUpDy2WD57/kGa1x576KzJGZQ9lIhZmGhRCq/RnuwWOzqoC03
wBvAJz8rW9yE18lCpwGZwo6t0aMjzEnLF4FX9dvd9yGREjJay7+q3I7xEt1pQjnwCBGmAw9Q/nRa
+CTCxL91KKYrfhcpYk58uYpb3WLZvaCBdbfL60cJh8th3SDbbJFzBhc2hzUgYF4H5vqPicHMHVmz
D78Cd/BTLG77YtmRvirbCChVU9OpOn5570sLSvwLGLvkhrDE+xaKna2v1UHnKTxLPGQQn+nq1xKN
Di8cVDKUW/2EFrmhLGBD81nVOFUfvirm3KFRx/YyqVgrgjrUMN4Yk3UiQaX6PrfREg0uktQt4cTr
vqIGKKhZQuc+GgPTfmwgwAOez7epY0ItLZAyQfMKUISbSV5nQNXq5Ck5wxmvjFJmb9gl2pUuxwwu
h2+DRvqWk1ttFd8/mkgD/6Lmz0a5KQz95WkT/q5+NDtPHC/rX1jOZgDR6o68zAY4evknPdxZGIbS
bzfvHNCXcJjGLoHK064Cdw1modnk2IJ/JrS++CQYK6oKiJpUibWw0oJhNCJ8+/PjhvdG5rVD0M8C
ssThLqrOUdk9Xk4E9AjeEwgMTesGOE/1SSNe9QJZDsaacla+gsx7A30CW0BH0Q7CAg1b2bO3PWNG
C15tUyjANjbkLRrU7HePDiB1Uu0623ivqcRzI8kiJYN0cwTv0mU/1w0+3zazhuxBoUO6NpTiJ4bg
vt2SmzLPmotoRRf4JsD+qWVjZ/8V5JViFKKT+ASdGYsXWpZtUkkV787Pz9ubo1BnT7Q3nislViBu
yKsPWXIO68BGkAIVCi59/zv8rF3xU3H6B5jYhf4ZxRno71Vs4qyzLT1oi16WtQ9Oqi9oisEDpBHZ
FSqg8IPdi4UgsK3dJet18oohkDFl+XEhysxsO1rCnLqtuWs5QCmZicxY+S+Etq02RJeujmuQCKBZ
thz5T0kvXznLYfY9LZfxoPfx+19Babj12ZeNM1aJajRq+tKLALNG4VadFBvtS0oMzcuXhXtrvWD+
BqremxdbCtpe9Td5lyqK7zk4aotPKCIage2FTlbvEDsFFsRG0JUdEal7dMcWLCZdMFsMsiobIGKR
rKTCxz8hhCISUfPJlAjl1HI0Qassc3P4qu91KBrqkw/rVVxKITI8+6s3Bebzn6eI1BCI6UYyDmuy
DkV2W1ox2uhpzlFJElW1QFxbVGDVrpyZyhWcRN72B33D0NI6U97jrZw3XouZhb84xiSG9swuuWgE
ieM548KO5MqQBpUpz7DpUjeWFrMz/h7GbHR48UlcCxznwKD6fHQBilDE/Ddv/B+qnEpr/1ArVkby
2wYRL9NqyLUITGk1BFhzgMIRgMpQbt3lAyHNw5qAs8lWzBV+bIQQp23G7B+1eYN0Ol+KHG0ItTdu
Xzql282b005Zwq4jyB6Z1jwxSbLuq4lrX/0f8NBb8bIJrSnVE7bSEyPmGHcg9vnhUzmCvSNZyHwI
thbEPxxkBS13ZVc1X+U7cnGZFVXVL0vMfqPaG89fcoJMhyH6nptPZO+tMHOpT2FkyWwNgNUV8qOR
a23mVnyJmn+AcmbplFa+z80HZDHG7ryoptFw6GtNSFPd3angT3v1TgWZjFtYTEXQCkJ1+7KFmkJe
CEgV023bOdkycbBjl9+pNigfHHemOS6Xeo7GQi3qcAUDTup+n5UBrGAwgtsB14y/sBTXGhJQtDul
I94WPOE9upDPsuz9VHTTYl5xRBZhpd/qm97KZJ0AIimio0tD7X3KbT4YKQMMa6qififovgbyJW2Z
Xcss0cj/GQHocrZjZdcxVOKpCx09AduFXiNui0rzF5hoNsLgQVUcX+4LSmM3OwgltOJ5yCwL0Lyi
pxHapRODBZuNwEQz0jnAExBWOUclSInHbHGsPARvixU1kKibuYC92Ok7kxB6+QSPyaZa74jDVASv
t6r8/HTArbFByDK2GIUZbTufxISb1bEMlLXzqZ2XvOCYiTdt0VWr8xicS2iLLusX1u1y4G0jhW97
bvB4Ntlqx1lGeHcX4pkCnnhUQ+z0jwoHFnu/KuYz0SRDGg6Az1hJvBoR6X1Du8p0X73g+j7P2dXU
+BkqjfBHiOu/3YXxtAaMEEKjw7kYaG3sGd1nYuaSh3hwhBsUlIKToExMmorOpTDD2LFHRQz+cVmC
jF5AvLCW8f+wPtvrHtrpg0CAeFrYkH82ulTdF8a4aoV/F76lP2/668cg1Dvrd2QL/Veqp1vZ5ANl
AIEXpcJS/VCWtnKJ7djHtyfI+Qk2zzXRNBGqKZk/JHMEVWKiXw2jPeBypmWFzPBPnUgN37tGDN/u
FD/LKNK8DVhVSBV75VV/phC/35t5YOPGkxu46JbE9fXXtttgYsBpz/ITc37HKrZx11C/xm0aCJSb
5HuMUeaJetpQzip/4N7isxhggngu5TVhNHnQjDOXNJb/mJ/STa+66dfFhpMPgfDupzTFmjJFRINL
4H1LgAKG25TAQgQpluW/KN6mPZqmY4iu5hrUYcTmAqhIWVOvANOQyhypi4xoGD9qvNxzuMRrB1yF
tKifUxBd7CwRiwbunDLLbeJUNbHkDQj/oKwvAmXsJ7SYywV2mnvox0AQv36xguJhnhTxY9hj/Gw3
suXazdUgtJprxnRmtBUQYgy7vxTWxsmth5/OeBeePmGK51d/VAt0a8wYbJwwlbs6w/P5sW8YP5Yn
XPt9Bsfp+7Sa0Xaq+b1E2BhwEpbQSYMIGt5qog4bR6EOb7nFcHSpv68PS/tT3hDkiJIB/Lgce1fx
g8LSopQzzsNeNLzhFWy+60O9k2y3/0EqQHpf9q7cp6mOVsE3YBsf82aclFSaP1zj0Kk2dlYDMZZe
3fHpQBz/0RD2COr2M1Tjb6rIaVsRyyIyc7qWj4G3Sw/+9faluoa20BtsFDKMtAg4GoFeN2UhqOgV
IoYrFDgQ70vRDgS6bXwWZrACQGwneyJNUvi1XCzwVW1rHssRub8XFwUosvu4FAzWxYmlWYftN0Ix
IDOYX5QEJyiI3FHgdr4cMCtFRwnS6VZhiiQUseGqBB95LdhrKuSIEZISBqD+ypA1h6a6AaNWW3jN
R1dA0M8HepTTLLEi+FpTsXgJ2S2xm9GhXYeAJLNlcfTFSZdi1SWp6qkZjPE+CK6QIRLRAuTPNNp8
JIHQ34eCoO0NCFPewUsZXyiCg+Oa/JRohxKIFvBuHuyJ801ld52rLomTsu5f+DIZ2w5Lse2XIZ1D
602f0BLUaoVLvHbjxGMQnozrF9lMqJKuCj1b9A4mi1LWu+NDXGpuKLNXVDFHg8dzvFv/m8JWmt/i
7m6PBLSv6r76hxgnUoT13CCfTW2DzVLGoLKiuEa2zAlK4FXFeo/QomMf/zocSmDC04NW6sCQgiXJ
brWWE+6YJlqaRz9OYJ0kVXLD6E3aNdzrlUmvKxOlct7ZrP48w3enqfOCJle0bEIZvhtbV12qR5zO
BZ3AxZ9CKyI/WQffmFe+aNS8Uqd2euhfC4QUaD/FxumPCZKZVlAmjEXIU8d1bOn+Hi3+brU67GeE
oPHdz6cPQurvsCIerb9w59joTDi0mIycGacchEaGROcOIPyLlD9zWwMQ+iJm3p1gs9a7Lb+rNgSu
EykrY2SHBZJOKX3SaY76DEwq6rrUiggBY9Jh4zwD9YzTKMRckbP/2uwGTYUVV1Cg2jXBngUq7ZBq
QfSie4dvsa8B48nBiYw9JXb21T76gUf9svbOY6W4ISznzqo6j84StP3Tp4b0Ob1I9HAX2460sKoQ
y6Gj5J+cm82Z15hJ0XqIhJSXoPxcVhO9dTtdzPt/KXXwVQbYnLgJqmcS0ErZMkrD7swW8cHgclUv
lIyKjwyP7NWeDlqCvPxD/s/9xynTDOTAwYoNvWmYr4jEf74WnUW5tzWP4A+QHucmOerg+88VDr3O
Bu//BJFORS19d7j0BXLTAztvEHP9cvcGHyjuL/1hlro3roMeOUhjfFwSZvYo5BK9WI8FalOlwsMo
9E9LrEbaXg0zMmjRRLFtbXHl/6xAf9KnGZvJeqK+oRTy0pVdy7eW/806E7z1HL+VC5JftsD1NaL+
fb3hquUBQ6284Ky3RuNxtYS3AcHKkAHRFIeZ0QsWdhGr/Im3SIBA/lvMkQAWo0hgjw+ieQfUhFg4
cuFctZ7wt7QILUet8nn2Kl9YE1ydN+Zzekjq4LINOK7/kD/HdyrRW8Q4AWn6yDwvPdg5RH5YkUe0
hWex1np/ABQaDKU/IEe9JOcL7xvQoui0jNXj5ij9lI2QuVdLsH8LFif1fI0y8ntkJXqMESFbrIB2
XY/tYfoqe6K1Go3Ku5xCoTZ4a0P2AzH0IsFC/wWw4L889Tgb5IffNRk5DlUXAqdYe+B1BmDZqkn2
MitUwANeTCKMPRTZS+OKE0LA4frMa0zbIEK8j6XJ1PvRWzijRhhwiTTl/Xuf5ZtQ2srrssKUYy0L
2f+uTh/huCUBxg85eXNGas4HBHuiipyTYfQ4RZWixW1dqVlmHmVZ2wIKASRVGf2eotPKfEvh6oeX
Hh40hI3mQC89MwRXGvHDEPQAcmnwai2HZiU8zKS0QsSmXi2WiUVXzKoDc+g6uqkP7HcxyM+CDUj0
evioCZccRW9XnNm5eU4w/N+NSts2WthNtMPORID/SEHSUCwhlAuVIghi+pykTCyx3cCaKXGQbyOb
xbsM9/wXQRVKIdi/imNsJq8GV7/Gqft+oj3a1J/O94l48PdKOG61LTdQsx5ySxM0NrtFdwm9GarI
wIXIwWNFMyGPc20fTV2je+diK54Ooe9mVu8+yZ0jZ1KZlsgaAxciAiXfhBd+d3DS9iYD3MTlPWgu
nVQIPAwKjCgRlosamo0dsKFwre12azzu0GQVIEexbVwwwU2w97UKg2cm/YYq5tJEGzozeFoI1fLY
ZRP9lWbmwMne/T5Q2/4eEUhAPw3ha1nADFhcpkdxg2RwoXO4MzaBhgnTbLsNgws3IAE2Gq59QroZ
hSH1P+BnTwz9/JBE7DC4jvhbQ1T0VDspwwhUdcOB3irtbLkWKh05Uye0ihnTvaLXp7MuqbPQfKZs
0V9QMBweQsbghzsn83SYFigyWFiUvs+rXJAH/fk+j6Ohg7t3j2DRlS8Sem8BzMb22Pdy0H5AYJF9
LfFFJQj/4XFfiKaupp4Lucw2DouHsPszM2g0Z7I7w5iaIVnhU4ov5mHHFJ6J5ne0Q7jFeIMp1NQV
0u2Wbq/0ko3lEVATiR60NADK0Es+AH6wHjpNJTdjEvJPLkOoTl1fLEVIrK74yi3qJ6BTgl4aQFQ1
ujwBbRtsQHWr6qGLA97PJJxXPan1UPJgd8b46XU2o3FyRTVqEhPkC67Bnvtdpka+RG5Y0y6uulY+
Yg+WT4II0sPUlvmzYvgXbge36Iw0NHXqSbLhmxdSYOoEglFIVkTxfHnge7g5GfZXHorLS1INwc14
2AEMBrDDfrSNithADEK75Sr+R9r4aWirecoRE1JzMKbJQDUT8ENyZ67qoZNmeUmfnD4h9gAKIpQd
UtumegusiwarkMKb8cHbFnRaM1Xqa1WeNBD01ObK/odtDNYqoNtpAS3SnXuaJ/20ecVAz3bwmwPT
pB/keeVmFQVfI8hBgUcpZ2mJ98bk0WQvIayXQh5xHPbPlCog/+zyv0mWbdJ+h3mUUP8z92ld7ky8
lTUW/TLZHOaH8AWirCInQDjbZCyT+qngqjwD9jH/0ymt7YVmaGl2FDHp9jxcxugiRsJBY5TW/GpJ
Yy0WIOj5qREv0or2Ifl57v44tiGkhi6RecM2ZNaCqlQrn6bedo++rdCpTH1yKLdgKU8zVGmeU1Be
1YyyHA+096fyAaAKj2wKGp+s9bD9cfuBN25F9Mh+rgx+3WMjvB8EX6F3liDeYZFwc1bzQz/SM9vL
7x+opVavPo+3MEFw6z4D7PhAjNnW1KnuS/7Sj1NaAn48tTYqYJT0HdWCz17WUZNOEj3Wai6XScCe
XuFlaLHWBE6yan373e267pfOpfH3hn4VMeDV12sw9+UuIentuRvpoHgmlRJ/lupQdeDSRa0wX/R0
dNtFqozy1X+SuNtysA01TtJwoSQZR8v1f+O34SExVvJDffeCitz9YJzU3rAsa2wpQ3xXn6npYFej
tR7ZCrZ9yIf6Q7j3YGHzYhNmS93Fm1aWfDs3g5LazwlyEjLLHh/S2BFkiFTuv6HMkYxNKc5+cXkW
NBMt+I/JZqGBlKppcqqr93nzcP8iGE+2TfloAJigGAzJi+5b4R4wcNFaPsmExvpGNU6Ncgq0ODv+
HqMbSyGONd95zExC7PftBc2+tJEVGe7d+Zv9TmnGVLJbsYzdpbQcQIUWvrOZPZPeFBsXcnhkT5pI
bGwtNSKheAWIZmJAT+/IklDQzdSNVdBDEEJrmyz0B+nWy8jlyLXQsFOrRWXhz76tS94E/+Ox7m4K
vgFaifgsg2SHPehEwGCYAn6Yure8txxYfcRosisQN/goPZ4AZ+5LSY35zisvkJvrjqR1fmsEhK7e
HdxiHclDeoWyhowjvQBZ02SFDrX0/IFSBiBV1PL8jkRaVmLjtHnubrSRSKW1h/o6we/Snhlzmch+
IY3b1Poa6JfWwXzu3HomQAMs63gxl5LgAigwVvffjADlnW6DGn9aIXL35Q2R5Qcafg4m45ErL4vL
MZlxd55vx0+bQmeSIzaT9NlEQQDSvp6HmvlHDZEGKHn4K800+oBdiClbfRsAFouaGcNRCRFzAcWZ
9zp7JC7NDabpdxb/mhMQmC6BdLisHGiNZ13NL+ndmakYlsxY9EureKSpUqCC2zXKDNxoV6r5uowG
cgBwe4lfSMBf/724y8o5IX7hsj9OC0l2+oItCATAb07v+TC3NAdd8GNBNg47H5yZT3QmWGbHlBUs
rK/xmCiRkuL/b6KK6EWdFW+1yl3gqoiGXkStFxpvPaRPBAeKkxicRiOfD748mX4XFpX3GL2fBJfo
/DRPAttBhcGRalyKGqNKTEFgzv6t4c8Y7jUozMx4ovZ7Gt015ciOD+kCt7AorY9qBrx8YRUb2hON
7kQsYy3EQGOH3x1AHH/Lpsg+Fefp+njx0BGI1HSCGBXifueqSw1zM0gJJ/GbG6utThShAdyE8/+k
4Bmp/ododh0zw71XHM3P9IXVEVVowKaa2tMk88tV9+vEPrz+cNLzSyN1O1c+ZrYMVvagQyUf1XmR
8PJon29IKYpmYMBhl8buqqGhOM8GDO268ULR7jXYKs2SYUKpXc57IgbPPt+OzhymIyncdNghPua+
c3pPzuJSJtfY1VhnYVucAAXMPhtvpDnJi3LNv2K925QPIRcvWcKFg8OzKolM3L4T6PWJ6Xs+wuXZ
u9Ta77CgnGXBYRi/r0AJy6y7k47nzwNwnUEs3GTV5fuUFQ828AHl589EmPqo0QY5Q4Hm6z7iEq7e
IyoJxy5B7pp6BWVVjZ5m3GrA+aJPMbi8k4RhQBUUnJQcN9C+3bpFVH64MoyxIUQ5dJNKKtBeW/7f
9ZiLR49ixIepxK09K17ry+3uiikpR0g8zTmXLKJvF7I7hCL9MSnoHrQu6oFQO10bhP8P9VCChGHc
AT6+xaM/DXAOmrQoRh2LtzGuz+Fs9epFJMjqyizAqPIvyUNW2CJhtbpaBQAKAawMwiZm0u4KNJc3
ZJTbu6x1+OHJZyU+ld0/v5dk2RZObmfPyjlBNd1Kk9DbscODFxpNUz28WBUTtH9FQh0t9Er/xYnU
vshRbK4DLpk2e1TrZtXtKOg2o0Ee9I/GBU0U7E1P2bC3R/CJS4s/zUXU1+MnBS/B3cqwCC1NAcnO
7B3dLZnIE+qCOaFyduJpu++vEt/R48wl3mwUg+FaPLPXWNxYBYoyZxb31OjdiaRGZqO5R51GMqMJ
6aD4vk0J9O8/3DBdDE62zZGyqkTzwryU2m6Cf35NIFtlI6gc/y7n9QjV7XbhEM1RUkCsJ7Te6X8+
EOLEuZk25nKOQAiBzM2B4Jntwb1mwJUvWrREjY+HLjT7VBgsUIanvjpHUY+82FSGuT7VQd1gwrZA
UgB4jIhnr64SxD1zAQsComkM4QoiWbaFoi4vE/XxSxtKTOcwPskZEHm8Ca9YvqwKTezkwBLLggfp
NIJEoYtSNEGdCi5t2oUPuAIv0ddF9vkvv7YfaUlBd5jmCIDlGPq0Jtrf4ChgvsL3U4czcqCy2T+n
HAYAxAXm7GGAyK80sXDSjoSnKtH/IZ99gzdPJIXNA0G39qTX/GC5TH8UAJyXH4dZq4+RY+HEP++/
tGJtMCPXUQJ+62mRxNk9UWVUCE720/9WEi8NEOAQ9GILOJpZw5cqJhjYEyzG3DvXd0Awt3aN1l+2
9kHcSYtfoLPbOrnft50VNyA/35sRpCdmnn9bTLExGJjnheovbNHFbIE4s2KfnoKJOPVfPpuXavRn
r8OwiBPQR3TQQKO6z9nJRYH5IhE6kRM3/W0NYtpxUBg6yReSS/VTlw73YOfSPwUtHb0c3pIlObuP
q4imPMibP/L0jl15GYpff/o/3V13DsVDsUseV0xYNVZMBGdVBL56foT83IZrrulkB/f+hidp8vFz
T1PAFKmcEHoRDflampJ2GQChIUNNnoEBCv1WqrwYDR3WChj6WB6NyVFGXMw5LSFg0y3Tkisb64iS
mAf/CwFno1II//nSOgoe4MY2j5A/z0OOWTXPxvIDnUSgj/dR4QgvAlefW7GWyB8uBkKxOCyI2wX9
18mGKJ92GPcyU/pm/pU6DvHApWXFOIm832UDDIbWxJoYzOnQN3TXwtZSY2hM2/V4qINPtw985nKL
yfhVBLWKez8SMqHLe7DZmvmdhz1OH7uWicR/GPPoE0hNQbew3y3LOM6BwMM3Yj6IFWrP6OIg0p6/
PfZURqv4rtvWoD20RHNQgu8BSvR7ugwyAzetgpipMVjnrFVGc4Ht6EPPVFAtfYilN4KIXR/q9i48
0OZ93VucXoZKijuhqQ0lB0r27TqYZOMkFctto3EaAOuQt0e41oLbeM91NrXD9rpW0sQsP/yG9Akz
ajNEmlrw4wfAHEgTyA0yw+qLmpKs3rGjregHRCqeW0hfO9FORJpWyv18Ypqu8G9To9RNHiMLtbTf
KW78XvrqYnR/meGFNQXIW+sypbtgKqkK9fKiz9nbZJeqgE98V1RymhKlp4cWkr7XpjGanyzujX2w
oVcDmZ8XgkvTHCUf8a4M6p3AuKV8EorxHT/pmJlQ+bCSZlO4pX+bFqWEI3+liIGNAS9SgFpfhg38
nv05dz6Mhrij+yQlAmCuFEF4FP7+hkpcYfNkXlEYIxXwc1o19Cce9E/J/gnXMgTI/OlrA910NxcI
6SWM2wGiqJuY3OGyWpeTkdjJzxpyhH612uh9CBz6W7T+QpHStQP4IVvvdFZo8OI26SnpS6xyflln
PJdaqlOVwshS7GCsWtzh0DMqFMajakjvugQTwvnLPKjSGtepgo8n68QWRougTTdV4b9/11HQLrPt
9dENZzkAM6O1/ejgLiMfBfth39rzYvyRsQVahfxfKR632OVBz2J9kcLOeE4sHVi0HoxuT55p0Mp4
mOP7k+jec0abGLTCiIgyKZmwT4aZjztZVfY3zcNIXZUDTiAGPU+mULY1K7QOHi+QB3D+qJCecc3d
9+QCsw/u7Jw5/bdKWtuyE9VjkOgpESrO63oJ7EZtL1kGzqPHrGFrl/xg9RGad8zmySLg3HiiQT8A
wLRfsWRkrzhJ9ZRAslqj4h6qldOq6bU09iPRxjqCPpA+eeM85UC1Lwqa8LMGSguEQqp4OJI5DeJ6
eJ0vOSPGV9IQUNtv8cE6QAJXC1u+iyZNcTaBOYwB0Q9G0/6do/o8SZC2A2nMyv4xq84Oh6r+k1RP
xhVC70Q14ZdGVk59dmATdPjGGuo9aG/6F4nkONN7gyve2LuQxj+iNty4s+mEeYrQoUS71jN3a/Zp
8PQjlIDnlM/vcxWuk1Xhb9gRF3OOpL1ko8cYcbu9rzdPXtFkLS1IIBq5WXUeQJlLDHP2B7/2K6WQ
qq1OdjHC157wous9vE4L0MKpwJXlpJghdAC00Cp/bhbjlu8kEhz8Swd7VtwidKc4UrfDtLV4siII
QxrxsGlx6MOycv7C91mdhDkNJQjJxc+5TVUHlW295U1Mv+otQpEnw0kudxZr33tyEOumgyxDuSx1
IohPYW92GWOVg87UKx6tQ10MxNhb43LpuFMLLGqRoyNSpbXIVWTqj1D8J3w5UpQBsLhoxXMt5/aA
YpZvYXZFMVN3R1W9JvXBd3UbsAbpbE6bwVCwPBMF1Imuk1qHrLK/Yf6zOXEg5pGyckG6a78Ykcbc
IekYFqmDecpPJtUqV5oSnZ/zbGGMo2Fd/r9t5l+7C0heMkwIERCb73ABlJOZfybmJjm0VGEsfIeS
V2bHSZ57VKGgB5tQfd85DNIdmTNjdpW7xhgb4HJZyfV01v76rjJ5L5CrbN3DlW81jXR1CjbXGFer
7irxD3j7uBBOadKKhzOL3jjhSEg/Uepg3Beeil1mOTWqcPrMDNf3CgeFVSkTqQMsJPbbmS2cY5ie
fJY0tH2qn+6BloHdjLZXNwDq8FwAxjpltGZS1NWKhWrpUriNCvBQeMpFpovsfRJCTd+yaVLkZ5nL
N4hFO4qKm6gNH7ifdJUP7vfrMY7nfrzryheLuUxDHpiNXg02kt8QDX9k7gT5D8cX4rBc9UqZEyVV
Mpw/Kge/762f8QNmihoy1f7dZyTM49vrj++VH+b3yiGlU6NJec27gntgy0/gT4f6QmSdA9WolZ4C
/WQMNv/vsdVOjsVv/WQwS4E6lAlZHkJxsK7f0xGHvetU0WHH/PrV9fqB3HKU70MjdnPgLZ4OzdCa
pI/VYg9x4booDzZvEYrh/YrCt8mjsHnKqZwE0gIf3M4IlCNnK7qN2GUfNx9FFKzsuazEncJg87I2
uWSqYzsWW1WG0AtNWpA4Ghjo+j3CJqfRBgiWZ7k35qeV0d7yEYHT+vGepoYuAHtCFY+lX+OUH4WX
JKep5yJmbmvlgOzTf7JgxypWnCHOLyHUgCX7EqVhsiI3+xt5R7XCRGQNWRQdNqE/9F7luyJvVjYx
oH5Pzxq7owh0AUzsEERpF92judPpJyjsVXQ/YpUZltuXTUmcLZY992XhUS579IE+W4CXchsHwou6
E7sVPTYc7Y0Y2miXf/eAgZ/JgcJtADU+oPnpYBd/OSXKbt2dmf545xJ+ozO0F3VX1bd0I7WorWBT
JaEib8Oxdn45KH/GVYVoP2sNF843ffqFRYjkkeCuOf5W4/dpZXK3qXAZ9iDvRGqYlQ2acij7BIng
Vr70bYys/3ZrSJYOWaLzKmVsU1Aglu4zYuGVKKc09VSWbhr9mXZ9n+fBfvquIPBtMJYNMxiOLtRP
x5sugi2DE9LRRNyhp/7ox1CiGdk2N3KSaxLEka8ooReCyW+ykNJMubyuOH7sMb9VWIONB6NUI1/I
Wkd+d2Nxnqe2Xe9r/tESA5qSn5PkdI7FBGVB9oaG9ZIq7mXLpCcobBOI+wx+j5vn5CYCgxROSVpz
Zrt2p4PbPb/Dld+treWEQW+XYglabsZokn/dk49A9HWUAAkzT0jqBQXJTRexcs2iUZ0YZ12nlTgR
yqaxX3UW3V4kUXtyI9Xgl2MJqRbAyrIn8ElIS+URHriY+1EtPIgUltgAKaYAoPwWoG7+jLl5o2Un
L0VEveLQOl+v2B5W2RnS7gbpIqKBlaepwKgAnTHsZLU+HQZFkuihZkr31UTxlqvBxnR0pMlCmIIE
tAdlXvVTKQnOkVAS5FuQvMB7PAyJ5qo52iEwhpMRwd89iJGGf3+OORogQVuLcq729H1L+hF8kB/P
ZaXjmv5yIFVRsbhxoqv2PduZS8t7ZufUK43i38WLJzrT/LOHlOMVpB4v1hgPjnamvs/e8/kmRUtl
3ViwgQ+KpNOCdp0JDgpDoVweT6r32QX7Z7yRPJ/Fkkm58UBkX3ZsCwUkwkStJYCLxZYg+NTKjBLe
X45Mcyg6OrwDY9EYIkyXQL8O5lZTsLT8r6C66lqkiEiG99UEUdVdubftcyyJYWTfavzbRXFXVFqf
1dxURysLdEGiJpshjFOeA4Dz9lktohWaIBklvlZwv+JYAt9LS638yAX+1kqNZLzZ8FFQsrqLtz+j
l8tglskbVZUOcw7QV5hoIzbWvXbX2heLT8Hl3s+3aZUOpyudZSsrZ96dlEEWycBacCSzrMJYgCCh
V4xC1mnLzGtXgecdd6GSF4aSQG9EHfelLeKz1t06d+DWZol05K9/jnYrWMRfLPKhdu28CaFKNKBE
1P6WBDOai8lRZr1urTmO3zwrfOprqGdB5JCW85BKxU1tL5DMp1eXrM3fLXULfNVOovk7MsLAQUui
iqJQ/lDQAMtbJJEnrKeAvaiqv7HYXcpD01THEJj1efzREaka37PoAfM/sHirSr622pmHuHqbSsNP
gTucZePvJAtypHP3HFuyhpH0f5Fq1om7w4SW3w5a1trkndB8iq/lulXbX9oNA5PQyQsV1DR9gXPn
Yc1gDhBUuNI4KyhfnYPVlWsaC+/RTlMQhU1q2vwOYHHyB+pZnCBSovhz/7uV2fQsJuLTPSVg5vaB
OVW/i9agg9Q5iiqcWISTUFXtW9LoYMTUrwdkWvXQXHGJfo+KOHEiquvZP2d5HgKfJQP/q+fnCmoC
gLT/NKLf5cljak5xAE/xDQoDBlauGn/5/b3bN4ei9gg1YxAD2LNi7Dgt18Epk28E05ksvWXav1Ca
wF6SQwpMax37WOl3Q8VVdaVlvHua9IRMKhvHkL0Qy71kOJz1zcYbmlDsw8E54kbvTKpZusubGsQy
JGMKt6vUf+N2jHs+BOwcgHCs4lACmZkdH8JgC5qzol8VLdwxpdJ3rsGMbwCydFpsu46cNp+bsaYE
zwTopyRglFbHnxortN0zW7NPtTH8xzli6PhBHiC/A1tOhP06v07cvUG1PbwjcNFLhZ9aQiZWStK2
RT7zTj6gCGc74dsMH/qbxyvUjvmf1B9ENg5ssxuTP5UDBGWwLNZZGqj0hY482qAApjuJ+PMHiKak
Bwo9QGtBVyUwmhlpa60qDyr0QbkVGMwoB6pa5LmycWave8dgu7a/7h/nWPM6sCr5omX8HqLvluYv
+kI/B3Bzhymt26gmKllY1UG6neKty0PtZB1jr1S5Pyp95a4oRg8Bx0UmlxOSMMTElWeFU+akfyMS
hP+iPpgjqzedAkMptknEBMktAxyOVJFDg13bUcyvR3d7onOMO4aKi7byjV4d64x4LIppUiMN/3KN
SWqJfwjIRYUwrkLriPDlc4lbD9gHutMRNAmqbtqxLocgZafrvGctN0WMy4Awck7XcE+6bYGGXZHc
N6BdWVlGdR8/AUfgOnKGg9f2knpXdSU4LukRPOQihyl5M42CMpk6Lfa2X/KVackoHlm4fKikFoMA
Bo19DV+Z0/wjOdtuQNkPACk2CMyghrrSTZIjWPVcwxQFxC1aw8vuTCvWw8niEm1oTkHCo3WFhHeD
3ACDBklONQRPPHnVhp99INZGG/r4O0f09B5KK4Adkhjs0y4vnNcdbWYMAZcY0+cb0T/JDGwH97Gb
RagVMr0AzZmIUAlLwjekGhkLBR8cfR8Op5PDDLwYqWToQtLT9Kngg2Sq/6beaNcvzxlyNmTuRSg4
ElfHXhL6tTlloJntlNadtPrWSAxrLkkMu44Nrd5Km8NeccaHdp3WI3BBsUIgC4JvtpXbrcyoWVbZ
XqxPMnxYzWWnliyJHlwWtsLXHRSue0uQiRYM93b9s427ekMXgmGvLXsIS1xMv7XG3cHo3QFKd4Dw
AJKT1TPvaZP/RF20lPhnspjRsj4MyZRqC8InBB4ED33bUcyx21D9GrG1PnMFoVreiqaIrFVQF1d+
5ZBzJL+MQkP+Sk97nWgcYy9SfJylm46eZvuMXXJ9OHZ5fhbxg71A0oA6NNT5InV/LA2mBzwhcKfg
LOUMESI+YoAGu0rCpE16uvqeORView8WS6IruNxVTJGtPE2OnbxXX3aOQtjD7DzV4TFwAQJLVzS1
z7Hc2kta0Zsq+uHe0vi9Rvw2Fc0vMZnCttcyhQ9CRgjZUPNvHWiK05itE5fZtP71KmCeNICAL0Jf
uP3MvD11luX2NJLkB2PpWZD2iRvsasZQ/QGABJlZQui3vQSXQ2XO3PemPltrnw3zRnAM4Yl9RTOa
P5q512zN4ClqcK+h/ahLpyKPT6BLjwqIDJUTbB5GqdSiKU0f/Z/beUglPFVs6UMMG+Wu165BkukW
wSVTuxeb5KLrO61TCfcFfHFdrOIhQPa6auidb0JRdFMcGfUvaPWASVuXcLq76HMHLdpWNLturFdI
rVvKSDrGp+NmUXc27VVqwh9vjVJ2wPUGj9V7Kp4RtwMxeMmGzn+nBiuGl+eqEfwEQB6Q3Cwxadf2
PrTaTaH5sdbIngeHE0q4vRx1A6KIsFH+YpRAecLLsQB+AmpmtbYdK6xeIOOQLEXld5/7NOc/8OyE
3g1cfj1W2Ms1uoRjlbNs7sxDQQJorKH+6Jws5YlthtR43G1lJa1Hk1S1hNjhg+8tZy0vTeUhy4XH
Y4K8prRVPFlfyKGQmKA01H4ML7BoLJBxr/yxLSrAnDJK3ibp76J7mssiBPF1RoSFm7QOkI1VPEr9
rp3/HIF637UglydF0+W69p1oj6ZXldwmUTtfnZmQ/kUfwL81y4vBFMre9HJV+X692r4U0NVI6FRa
YVa9rdNbm8HHKY22zArkR2x4ZdefZJsVKqcufpyo5WqILr3qnJ3v9JY0bSfK/6TffpfR2U1S6Y4+
yM/wcqC0UIRfvYnODHZBN8+IYzVo8wA5TWDvDw8H3Q6U9PWYXHW97LVjaaPueEzaCX6JX3SRB5jE
cvG/8KgHv1hoh6H56t+znbQUAVCxDNDlDoxUvXSNHPjUcTFVLgzPDceB+puan0ssph0CVUewWlkY
waIa02I3O8PClal7ieLqD1lMjAO2Tttg3BJDJN+RjVT4tKjEVbCup6svEan1+nzn+WHnQpHiHuTX
6UyB4Da2zJD1zp7/9hP8HFWgUd5mMpMdHpKxi/i/PDCRi2U0UjRZGjHhXYf6J7gGHVgCKtP3Eeuo
MZyzb4UIvssO1bxOUVAUSV4vOpI4tFUT5wcldPJUpDU7kYq+/rW3D9QP8lbNN9SKc7JTi0b8zjKS
Oe0Ib2trp4oTf8zv5V4rGqVocPVsi4XcRNAnW1PQJCE+35xkdYUw3In9xp19xZ6QGrMk8MAuUIza
oy/qZVD+0UT5xN7sEN4z6fVoW5DMC8mCX5pv3d4CSDJAKnfrNc5fD8qA4WjzKIs6rNcKuji6U2Di
1AqL3QaXfqD7OIozwOftxQp0ZuwL7t41GVAX42WGu/Yu3yj9FxwUrTZyb+nl/YgFsfQheakpzTKB
eustN6xlrufgtEcTR4Qd0ryjHjGnYxmEH0uqIFQZrjxiPo+YA5oLym1owgpVnw+EJcMvbhRNVBC6
UK9gxLYCzisXpMrxbOyvuFG+VgcNhutL+fuFAnwHIqbZhR8CF2CI2X/5fGcs2AoBirfTOFJ5RB4T
ML/+t11fIm7YO/51f6lJFCGJYML5TnK3OC7Rjftm908RFWnbHM6RFyqJ4tjGNxIg0un5CaB1Rf7M
3ywdf4RZRERSVnuPy1ArMX2AlVCyrewh/6yK4sbQIM1s1/dCoJRdJ5l+y25S0tf5OdE+fv2WwkCP
FGgWXyCNPiQXRwDeeGROeJGAPfVCGMWl70MJ2OuSBCrAJiB6DkVame65oD/HwimpKIqb9SYeBbHz
4cnPkwJfj9wwoIIVdXVRTL3m79LI8lT8jBhcVy3A/h3RdbgbFm2gB5Td+HX3y3fUda+CdQpOAkJr
c4EzDV3e+e/iV6srou9RubYdPQoLmwyrh6MtQV1ZFWpJxmQdWR1Ro00lmGt75YlaWQ4h8xyijs09
Sz5SiayoMkG6BZVF4fLMsDHVxsGHp/hDWqk7YccUI5MdlP7r/sy0tLmIpJ+q/qnv0E8MFOo/0lWx
Bsmow3DqI5Uo+iRxZaoLrxETcQWLQUjPR4PjggwjRljN0SEoKkA90YHa7iZtbtkWcADXzfJUX0Cc
Jm8KIrD9NjRxIey5YLJimWFABMNCqiTck+/VLdZK4fll0PY3/wZimImpQ7XF6xZMO5lX8oiQPS7x
k/sRWPyli2pEDJZO9zumm31R+rT0mX/QQlxQ/WfoD/qf6sPwnDEVeDnm3Y04kGHhmqeDTOaya7Q1
JaO+pwjgGtxgw2s+rRVKLbrWJdDqnhw4IWLM0xCmdMdseVptgDMypnus8mtTsmQX5gmUVwhGVb1h
NSu75CIEcC8pTFSH2Vj2a3x4iommgbuxa567vhzj2VwxGhrzK+8wWHcjv/nQkt8K7xgdf+3uAyVM
kWIX7thr9DhsgADOLouFHg1X/x43GRxkxFN0Ymimbx6Bo+sy24+MDLVpt8K5ufMc+jjYxAhQez8g
iYacO2wuvQJs49x0v7/sPWvrb85EBgPvOlCI0BwiTVScNM5IhSrFn7w7emneQWr7OsSqo9IIIyFx
nxtI2kPuC2HtTVZdKmCdjSDRIPk0vkU48u6Wj7lQ4i6SFoc7gNDLczCaFITn/4luKDcqDNZM4IW+
itJXM87Do1y6P4+eWy6fe+FEC72tbwFTFwMf9XWk2Hy/HjuqpUjrCon6QVXMoyCReALRINgy5p3W
sYmvd3sR5dvLJu16mELXqh4juRedrx9QvPNX9W8F78xyP5JxuFADOfMeR26PPHcr6AxFsc4gusQ4
FkSBVYy5IeTMBNKfdC4OtjCSUtn8nLcs4TCn8nZIR5T464ASvYqLIo2cjeasb5dnSaJj0xFGUUWr
pBGdJcYc2Rb7nq9dbJ6xoJo/XPCvNpGkba/sr/ePvZztgnGhn3cIEe+xC8J4qos5N78PQY68wyr6
UWoSnBRP1tnCjAr5b+Mmp1QwE7Fw+aJ7TAKVVjatVkcaCzaNz1BXthAeJbUv6KiMjRnc3cDN5unS
213YsmbSMkEQzRH6rd/VTUsq8mfAZ3G49xnThRHQ9YZkarkoa9nFlzVO2Wa87wesSMCwybupkcuC
2vyhQcpvmIsDkAl7lgUstsOmZMHtKsUIfxAYeOfAHDl3oqb0zRxUEy24SZGLykd/s20prhy9oC3B
HOahFj+52odDeWse68JL56YC+hUZFG0z2QeI92YvNAo0pcKJxeaOrH625ZltbHbmZl5wofM54OfV
W34mNJgmXDTzLTRm8jbo6vTRNrLgRUPc7nl2U20qH2IG+A/dLsloFUQ788QJADMyJriW6L1FlYPt
VECclkEvsTLABBFiUeE5LVl+RyaXir1PHHf0Cwfo7Y2JV4lJwTn8CeRsmY0Zkoy0SQaGF3lL+pF3
j5TIpARf8lSSKc0BT+CpLGOBI2TQRsBLXGG90ZihEJq5ou9UjkqxO+0u1/U7+rsnY+VBSIL0Rmat
+FtVG77luqXEG/yN8zIIfxaxUK5rFfiaPexX8s0tdpVUbBjsVPpTZWLlx8T91d/US1dHozL3hmEE
+ndkLqfPqU1OHg/aO6jWxWP35KxkXlKSyehfopdAzN7nIMd55vsqcyRDhTRYBhhvyxOCgVoBH2Qd
LO9h+8rSCuB4YcuF1vjUCO8yETEhp2BB7TfXim98ADJ6QO45dd40jGbb1RKBKcz+WHvmdp+987Nj
LT5vOsEVwIzgQlgfQO3WSoxSDys1rV7HQTcZxEob0gGRRtx6WUe2SUipATOv/vXSEB9AsZcbLhQk
G7e52duHGDeWxtmysmy6ChIOjCLnDG8VWUF0eVZr9xlZgFzIezd96arP/ZyT3Pvhol+2cvgGQeO5
O/Huvhh2IHqblY9dx0PsUxTgJwVvmPi4EFyC6dGHk6lvxedbH9jkMIrr4vQnii572FLg2R3BBkPv
c1DoKXBSI5Otgmhd6xOAI3mr2cY9JRpUaDBq/cyqedr9CQmdqKWARNqvnWyCW6cmcWQxGwTt6a5P
P3RKFm4IwG/slQsS7j33uS6dddlwMdfbETCN3Iph1lPbCUByyp0Zsn0UECaci5LOqnv8F2ECxWr/
ZmxqWrKa6RqXajrbEMzNVyUnYqaaLobw1ZtKQNSzoteRlXpWjOqdW6YYSwQK0IO/meTByREKzRC+
upB0/uL1TwAYg3LpbXi1NDKRdGjyUUKcA3KER6BhVmuR4JNTFCIiYz8lCsMJHF9F/tWUvnydGwi9
rGCD6/yxB1fkyMJuRs1o8MXxA3QIR0idKczr+llh9TLMnNnjTdt5XxlPtG4RpkM20Mu7rugFxfpF
+uhU2GGGsiSRtdSuumR7HDCIIGFJM5Psc1JypjkzCmzB5cggkJdl9d0/P9D5fQfJHt5ohrfylSEC
Mf0ZDE/T1FGove3FN6BkSMYbnb024GU5kb1V5F8aIZMyR2zsAdZDDYXAsrLJe8oLQYyYiV5F3Lfi
EXf2COvw+AIEjQ3WNrxT9K0NCMtZ5YgrmhF6NmN5KralOsqavCUNvevGGTgnoc4waEXxPSHqqhs7
clJ1SDe9g6GB5A1+1Yo51fBdd++iFEePIItpIh2D2iMuoV7WK61Jd8meMTgOzi0DcMHun9ZAFuCq
I+XWWA/+KlR3bXx67BmbZRgtidfx+jsMBfqPV55lWr8SrehuFgpbWjfEawtFGLL1PmtgJq1EwiWn
HKYK2Oa6GauPobZBalrhQPQRYJ+KdRQxqlqVIyF55i62Mlzucl4B3NouQXMD+QarJ4sFUgVSsD0V
e/KQUmGIwYELVWLzLgVJzQ+kFLVRiPCOGgMByIuDfjjc5HzUOmog+EYUerhXnsmujaBHjyZc3nq4
uxQWXVUe76nbsId7zFBLtW2F2vL0Pt2pZs5Z3dSpO/Gm3QvkvoLpBX00refQ1WHpvz+9rBXJynbI
MzlQWugzFV6lg/67xVhSDzfdVMaDId3p7+EtYva46FYXo2+ayVptiEDDihVq2OnM5l7hkL7FFhdw
nCVsJ9vYoLQwDQHnayMvA0GRksZVxewf+hxQTuDM4uLwj+5qeFV7BSspxkEUyGV+FHwzeX4xpvI+
KDQbHfGLZos0Vp6zgniVCY4HNm2dgoXAVpNbgE+SoppGLPq36kIgzUe5ZcGuCJ98nXbncMfqlPUx
ThOtXjZdns8SgwqcTT7Uxf6+2N1cP1rpV+NOflYtFA3s5fIfy79jizVTS3kakpOZKE/4RMZrwM0x
k7YojOUcRDnKdQqFS2F7YXM37AxUCl0ZWXYl19AGxEuW/C+QvKLcvdHM412nzYtk65uNAOjMav3W
rCTwiNH/HpElBK6QvvwGPD00hCxZa9yIG406u+AkobyH5TRzOxw684zS28kYVMvkmush1s9rLNvW
27yTWd+iMrui3MbS1fC06sryabhoMZzH5yI9CFkRL2VHBINymOMrJBEKjebzy8lvbn2adiCPvXgh
acb/BVyck7EDrLWtUhNokQ1W9AMFVVj+VtMpr3TNTALIz9HcOa7BFALlMm0HeaIg1xVVJ03Oz5Nj
lH2JJmHOx5JuZWBMIU+wl9RUFz2EGS24gVbCV5V8Fp7xj6KVy2ihB/jc9WpBm5/Yr0gRBVS+KGHE
tVFfa4tmFAh/R6Ker2Z4cU2uzTJAjsuiDB1nfvzFIz9FdV02u0NybAQUyvHeAX6Rc7hL1QgcTG56
uvcp9QYVsuQYIrwhmuAqhmu7eGWBu+08mOQymScwpnly2RHTbZkYcZKCwbCmj17b3TPSvlskGpF8
18GBoL07X2ktSU5uxaYRD5XzRhpQbdeHrUbA5J3jGwUf2RvvNSWjTFZb2dQAJZ7X+ybqsVHpulXs
U7n2N4amge+3vdMJJsB/sMrOndYPadKZq897w9+duGYX5Uqi1WjkQQQxaA9FHR+cA5eZJQGbQ2lK
Yto8XXIKVy8HzSgRf+VmzFW2gtQpnwXGRFNukcYepLKMLKNRi6r4vFJsdYa8fJ1eh1qSDvkihvBc
VeD4Bi04VlBgj7PYh0iFLD2P5BgLk6pgMfCuAyUwBN0zecQdeJi0x2bGjJr9SxjoEylTsajlxQMU
zHdHssDW4wOllhysHinHeONMe0tmfgSawHP7rwgpYNdWrjsprqNCntLdux1xxtDqgolYsm5kdYk0
pbEL1U6PLcI3l13nTeoTo8j2AbuwmKQDRWS6U+/IRFEW/wYW4DJZKL8H3FrPICif0MgArLRVqcBv
21AM2k8dj/loImd5TCYeU7+JLdbcy3GQANVOaoVVh3KMbK6JM3wNVK/S+/BIZKgn7wU5sM6voJPC
532pECKrr+gWZR/BlQBLqDx75vFcSG7UOjfTxbtBnwKCgXsv4zIM2+NgeaatBf4iWXoRmwlNjJpP
coNYty/3tfjntkmOdHXM334B/2uEVK4SpwhvOUwGgmToy6Xy6NLy8NaoEJA2KwXLvWMH9k8yIk/r
68QmlzF+Mj+/uNvtjxFWQ6vNfWlkxht7yAqGNgGeqfGurB3GUSNEH9ZwkAPgH+7blhHyETgICv3G
f0F07tnyaqreBZlOt3LfzZs14OOI4fsRcN+qa3Hxerhmqg9K3ds5KQJ9kRwv7kKuKL7TR7EsDXWD
B4HB9qR33OtB0n23wkAcv+vktKxZ9hRP8t1fXeuzv6Ijc11/fZg1B+8zD0oRfIpMbfjRCXGmqSDL
qlIPK9JZL9ZPS0zudn7ZcKzT120vN0/mLyUqV9Sxz1K/Eo6LcBOQMIXaBfugID2eFe9li1xPiHDe
JWtWHVTQZwnMAUZWIAdoem8xhX+Q59pBGk51wvRCrku0CR/uYgAnhKrj5T8JhBjVBT30yvtNKcuI
jDzaenmgFKlg4cydwe0FV/Exfh3Qlt+tX/kl2+uki7BPafZNJubVTzcWgU3gsWMrMNfFtYJP/WtM
dBynbXftmwgfz+TBcu6cM4nOpfPArWNyPbP8npkPcfH4NS8Orj2wUnSG+MDbYM9Amw12vwn/GeIH
n3neu9AcKBMPcChWbAbZt3K5WWI+41qrJb20av0qxvNfXIRbUdTP6r3AawGDBoNYaGtrzg7tFJYt
W8tmeP0qZbrvYMU/eKfcIczjetviozx8ksjjTlMEQeSpzrMWPEpy9KUE7A0Yvc2oE8BuuMvPxkPj
urXd8+56r3o6unL8aQHPY3wkhcGrVgQ8A5zMekk2TqniHJkr4AtyyxWNVkE6Ag8f2/zfI4tO6oyV
l526jnUEaBdHPo+yTvoDyH+AKd7toga/oN1LtX6l+vxF4lhZpErATU2GKvgw2qqKs2h8d2g/5ZHB
pZh+6jFBtgLnFFFBll9Olott7vcV8kjaaddaVy9BUapyc8kAtkoLQv7ufpvu4VzMyOD8nCROhWKs
eNtO9tKQ4h1Mi05Mq2mRdhoDZbXghrl0Sxk6hwx8o8csE/fnhvnBzzUAEMNkhAAy5m33A+mXiXIc
XtxKMzVzW6x356ZOQMpVmxN3Nt/U96sD7BJuGA78Aeox0Q/sYWCQEPjzBa/tOsoIJW/IV1wWX3Rx
L/NYulv0fPpPpexcBjKE8CgsDXoHjuVMNrC20AJeiK3YN5YAUjSiUt+Umo9IWMGyAT9nN1gELb0J
hlW4pzU5JGoiXcl9Tt6VHBOumbEw7twWdRoaeoQcqzhhrXU/AYLAucJ2AdrkWbshb+QUZf7BLhtA
a7etejdP4Wt84NDQdw0sfwITFkKLunCH6zU6h5i1qJQEQjqQSTFFVY2uEsKa4PnrwGCJGOVsAnid
tsJTUfThp1aPmxD5boe2eTvHyqmc9dgE3/YJA9MTsdbp552g7BmG+WV7B2CaN4gXRj2NUK0vZfK/
mG7jedvQX6m0MK39dIl/eOJy66/lpffWPHzOGFGQNzmKqyelPk26o/CD1vbJ6zEvEO/tr8si55Zh
zZLhjGm5vIpnU4ueWYx3epAryNmKK8zXiMnHcx0RPOebanaQSOwxPt7ff98ECG0u7SkIh+FTRzQv
fGUGK9tifkp35NmwfTn3LDORqVX7widV7PI2X6xfR93B4RZX8iOXJtok2IWKml+Ar//lyCFn8jZL
dzmTEObR2yxhQlIuo1wq5ppCN8QjIJ9PpLiWs+zVl4fmXxAKHzHp3peMIVW3s2pIEsKcPnkjKUJI
qrKFfQOdtgJfNHswO+lGVn5xuPFaH9wXXlbiyRyCo/NQPbqaMJia/FdhWyluzDFJHJtU4ox4cmqH
FKQb7TkEA5XyH+gAL9w4ukU8qHq61q1y87KLk5ZrhrJxaXMskv/dgeVtJT/3oxldCtzuXO+XE3vI
2fdhZZasdfjFkUzxSU1DsmmUWD4BHqWEB6lKPDMOfK4xJeDGSb+qy1HYGYl0bDGqNQsOBu/2z8tJ
nk29R340Ef9TT1kn+f2ayFHnhGqJhg1VvdHfXFE+a7uYvYxbIGUQ8XoOEsG56APG+0Xw3FJhiZfw
x1Q2KPbtqyblsB1shISFfC1qKs+97uNs9sc/DNs+Gg4K22k6lPfmE4uqwcDBOj6I77zGB+nO0yU/
GLLOxqZ4zZVH+K/kDQuV2VrGxNktPc4YIiJOocfclvtxbKRLg4hvFsQjBhvgPJQ76JgZlKFJIPiN
ALhwoBdGYY4WEXfrKmMo5Bq3DMCBEu4wr4xcspOffbh/UgMlPnIqDJZRpYM69eeWtQJqiHtCQFX7
P3Q1jEq3tL1Ke0L+kkqY8UMrbAHe6kyCJclckiLy48/1hM9EqQ3wx7Wn4ydXskpbgQh8ZXqII6jr
bsiCY6Sp86WBvVLdyKoZdimmgVS1/c0Wqv1HrbsMc60YguZkXRNbXY/YcDSSTkSbuZE/C8OZJXqZ
7hQIcGU95dnaSi8ETYycwQxSAkmG02LQM/Ifc3zBxTzNqIPsXe4FcQW1IasdXNHKsTo9HD4ztQSE
AeqYg1tI/4gzPuS66WxI8DRaRqLZ1Lx3ih8iHwC5adCvM26ht7dnl6HKjnUF4+r6ushKiJ3rJWQh
X9CC3zb3JukR99OqsmQUIeUoUic+khPIrNfJ2x+cynjDwByacBmwVNM8uZVXWl5iTTMeSdZAzDXY
7NjRTroWvKuVUmMV30R6b2QN/HSfSek2YaGLtOc/4MWzyprPid1toP6H/Gfwveo8vQHakhZGvFD4
q1QWXfaldtX26hdDyPkhVznXb1Vq0XKLuua9a8fAFIV0RRYvwfwQ1T1jg9JHLnL6i9C7XiI3GoNu
+RRGQj+InP/1aZAypKJrE+tetKS+SNd9o9XSyveGg6R85v6hHEJaJGNjML+9srRE8F86L0tNpQcL
ZTE9XRIJisBC/39Yfgqk9s8VUEVuFo/3WvpLquxrktEojttlgo3O9CGgLff+p/RqewCxGV3w7SN6
g5CEd1Zl7xpmr2C7n2Ps5LeJ+tiEkzR3/wTDOiAxe3dmay2NecS45SCRqGymmWZUjtYpHNtE31rL
bozeUXIcNusyK8Hf9ms8lIJ7jXySDShJHNlDKVUt6g7Su2qsNUIU+6otak1n07fGEs0DCTzDlcTE
wmk/NjzbtqwTu2DcI717rxfVMe4jfgMc9+IC17BMwMm50n73YRkZyt6S2q1x7hz5F4ir5y71WfqZ
eIGLrFLjHP7koCOH6AxP/a4N48rSkpqvsGNPlinNDu6vI1avz22mouLcDAmrzdJ7N/zDpIlZR6AQ
ZNY5elLjhHIX6L65AFm6p+NQYAUN0ut/yDgaVqz1ktKbRj6rgO4R7ZJCF64GGVxKQOL2V4UEIrq3
6NZEdeS03rbedr4lVCVBBl6tpivDXd08qeCNEbWSaijRA0LEopzDhVVJDSSInYUm8LbPi3c+7fN5
pe8qF8C5iHTwfAGaA6HV31rDtUupKVpn28rbQJOCkjdB2E2t+nsI/0d1XEWv2of+daqvorAcFprB
Lzmp2Zq17VmBH4ykBpc0DCCyeYGCZjQvjMbqyRfUerbyw2cGB1KFSwlMhK2EgyD2LR8J+hHrcZoR
lBchIBa9w9j35YAv9Ym4gO6sm2QawDlwiCdNmSPyfvBKN5XgiwYWgaK/Scr/SH0WaAVtRKPBj4NI
7UhbIUIENu7XWa2wM6PayIx/yEhCtiY+ZNo5uW9yoiCswsrXOlIGwfskhJcp1riqqtwm2I32XdKZ
xcvOIYKNoue30qVSHWJk2+mi+ShkCdwzi+8I4hzV3d4HfNqyudVK0c2L4kJmociwXQAhTvgIt6kS
RrdIQjJ81oxxYVX0XNCHKLb4aKyGr+Tez4+vqBcD6TUupmvlAMIwl3bSqq+GD0+Ttjrhi1Y7VsRe
KD9GfgRmqOSrpXDNIvMpaOTXrkOP4KsZI65cP2Y6hzVxWFjB35Jv/Jf6WMVvC1UqPx3xDMUtoLnK
+rJ8IurOqushDcCy+DwtFK78zPqv74Y9fXrMjzXeRRICmA7auScZWaQskd1wwrNmIjP487WJqWym
FtJPDGuCAOQJ1vB9sae8+LiQHL2vCs9DF8vMzlk3GtKFqg+HlMSksPg6f3u/2tOuMrQc5tYU8XmK
G7h10akQxTzTFlX06HlWGk8CkNbeO7UvPPE0rZAlI9B7BlP6ZuxhE2d7ob+db3UxLWSNnG5xfVwT
YUrjdzhRRY9ckhCyR5bmh/P175x8eBi0iTTkYZ5KlF8Y5RHSNdCJ6F3Y822yjhIIST6u/Ey23ZdM
KWB9ymAtQjPm401xHWu4Ojs53sh9PMQiVPYpu1rTnbRfsxhCxX6cqfGJwj+cV8TX7/toDQgZjxN+
JwZxv3FCji/YkoAm/VRutbawEW8utO8E6Fjvi5tpUwZBSkjUgb2dD12BmKdBMImhwAk9iMB7OtR0
X7evADtWTmvhV9KqjrTXOhrKK2V3hVej0fPrb1WhNd6Ji+6GCmJfgpF/5gov8QOY45IbO6ymTXct
nH/PjlcHk0kaPNmtcIizz/Zn8BsAypH/BPZkpFW5l8sxcEbJpd0fRya9SpM5BSjMhiIE1cnEkZCw
iZ9KkzE9F33ha0YM79J5RsSNvj3Cq5nXr6C53wizKWDKLmsjhwxIDeCu/86KuI8iehsl68nusJPW
eaMD2O6sBVMAiWYQYpjMRDN5IJdXWXrZ7vpinCn24B26pF9KSTYFxP64IkjkAJFFal0FZcpb1c91
KeZyE9U6HRzJ/HzvcusySnKJA2oRGHhw3dxqwg5UUgWSPmVLlfSHuLV/Oh7WXv0xB//YUMthQA+l
4tcfEJ1yx8gE0GUOF4yav7+bAL8/P8VvskVDqJh3s7lHsZNyEXECTY1WGPzvrN7YhcGzjPUMkfwP
gKLoSNPp9ydBHqVm8T4IIBFNPc09177i3nXK3W+LwvchKKA16CYc38puQRNW/M1bhXGvSAvrtVfW
R4CZJev7TbFoHJX7iKBddBTO+LhSEeL3/2Kn/Fdt/eLqHeha2+iQaAdUqAFlmCgMOySQdYZcPXZo
WMppcpBOGQFjHrtlV52PUKowh6WUDX9SPipwQmw1Q2EGu0LSkNqoGjBTGOpXFsrpxg7S9QGsRtlU
rjaSzx1gYmdpy6BKowTbsytQ6MoHDprKkQkv93BSjLapyfQJAMcBPI/ZnAfQk60biWgEpZ90dFmT
eWdqf77wPGTeURDkuCoCAx56rDru5hh3STBxtTsmrTIIoi6MwEsGkpD9Lji5qojt1Rmioultrphu
JXR3V7G0ajlHqNlZCVG6sKW3nsWQ3rX/yhDMzGR1+AktYlobi2QVourkh7HJtg+un0XHjDWr67df
bTOuULXAEGG3syKbetOPmdjkxBicGqOTPlIfP9QIQMkc+eGVTv3W4M41G1s4mo6RiduciHr2DNOa
zjZ5i5fqnAZ0e4EQ/VqVekAJc1cVDgTsatrKozd6n801ijSLmp4CJTStb3Rc/WoSYZtr2LAMwZqZ
2L5UIeRTlytmLz2nQqE2ef+j+rQkZGLZr6a2+fRXcP0vvDTR4Jx7DmTOhouE7o9aXzdna1xtDZWP
HFVW5T++biDSdlRFnQGGiO7M3y2KwYW4fY7d3KqJuA+bCqK4T5xktBEwjFLzEl/3wj6SflwyCpMe
7qcSh+1z+hlAV6GgXCRoeZ6cFGPZAQGKLyJ7cQqo2MQUjm/bGv5m815qnZVnywCHuAvyCxz9kIVl
ivRSZzhsiXjks3gBYL4+krbVm2vehqu2KZ2kV+bW3Jm24R9Gy0YJJ2p283UReyicFr+3bQw9FLAP
eb7QpzEtne0Iv/j8g5v65OkDcy18VE5eecJfkHyrqbTyl4PHRHulgmIVGkS4kB/RGleHSRC4GVM5
VG1kXIIrOEffggeb4gMJBubOm5U1AQseTMisqQbU+dCT6wSvbO4O1FUG9mmYC7oqj3vhxFAIgz81
pSf//82IKIlqxPF/B07k0KmQ5TR9AKLCaKU3D2T7Su3dPJHdmprzswvneAX661ORLBrFN2Kud2jL
lecViLh+rtPn/vMB7zxPlp0o4Ne6epTUr3aP1DnIpPk3F/Vb4sCDLDUW0WKTYvnuNKouqj8vVLkU
SZzclVfb+Tp5N8UEvAFFYLmbtJUByJgi6/kLD/QDLJM0I+sXSOqSJXhitfo8bfHOOTAZi0vpRwsQ
xUICrGTGlg1mIwcTuwg0u9/kYveZDhV2oVYxeQ2nw9IU/HhVeId2OZz0GFhn0VQ5Abs7zFxpcBjf
V7xXJ3/5ZLyQLzN0FDGAO61LhVPbcEP+DVenvFmKcLPQFI3vJABl9lzHiZHPN62QGM4lzopXWZdN
HxaJOpImqVQtB6cQEumkdqREtg3jVFYTOypY0z+E7OHVTfHUTaunILhqILlOJ7/rXdRT0ZR6vWf0
w2+IAM8T7bzbwo0fKCWENe1223xaYPSqbtgX/SZ28fyCmDKlj4X/7aePjB/v6MBXb+jGAh5fvaEn
PXv06yISSD9s00kTuY0kCul7Qr4nJmbSm6bJ8nNA4MrwHtSg+wjr0aazVyr07B5wWrmjwJUnNtxI
cSsz+BogrQpiey8MrBMucEZp5v6ne2qM0wZCHpHY0KAgOhIe3KacZBXVlySJoL4F/Ue6n+XEkplh
Knu8y1can2cXQi8FOL+ELBgxEuRa4lm+Fyu0rrY7PpKrwumYBNlADraiPBKgfeEHNtXeR03iUJWd
lXKvLE4JIC4xfxEIvEgQmLLHJIzahLMSneVL4CEf+t7Ega3l2+O+LHIJ5L8xGidYmrq9fUzAFNJ6
0DDa/JuPbyt5uoxaMO+yYhQDe5pStbGuwYjwPijbVqABXBSB0xbXLdSsF0jaOZ4snVaZPRFGEsLL
1C4NcJSc9T4SNomZAgJGBVTSwfAtJI6wpInWsvQvMQ84OjwpkCftI3rZKn1ToXCDyvJUKBXzNZ4S
LZGJnQyT9IMuxhUU3mOKQewyoLP1UV9AL5ARhFAKne7sjys5LooX8b7YOkw6jflzKnYCaMboyj9S
7cpmX0BtQN+cIYYcX/5r1dnHV5bw9jiygBOQ4eXKARPpDdH3c9pY/MJ1s73Hlxh9Ik8XbZzwVMty
eTEXkh5fOipcVR4BEtCvUDiSzJONB8J9j5EI5eSC1mW8ck8SGPgiS3lc8Otc2BiUsaXMaJLu5vTd
vCO8yoDK3+O+SX6WqniAusCuAMqAx8QboyTf3WGL5qleVEPSdY1zc6aca+HDTpJppn7KApF8s/Ux
2w3N7TfQYfh4HjLHnQPbGJW/LE/69tM1lMALRtUPM/qnYC0Ueqksyj2DPEr0C2KMCbpPH1xjHBr0
NyhsROuHb3KyB3ZbrhvQ39Sv3DDmzjzqFIHfxaIkKKPmVpNYAg/T4I7gMNN35k0Jr0JNXx5vsaZP
B4Rshw8jFqcmCTs7v66lTHars6F5i5ZD+QhzHensi2MMlbavxCKWSUSv7PwHKaIrUVEP/C2b90KX
7gQmT4HUgXrEBRtsGOanBmY8zuUb7XhSGtEHThJWgI6Qu/aJmVNyzcUlezGB5kv0jeXuOp2kNcIA
/ZZBGWBOWIdtbtvN++QFKqN8zXUB45XFHFzX8KiGHIvdhMO9E8bsj5hDjb5SnDuC+rnpQyly2FtT
+BEbIZBacYkr/8tlJY3fdkGqwo1aIeur9pDjjN+RmuZTfocDdkdBhE7ucroWJ7CcEPR0d4W7/Clg
V+kQOJCiqgb2gUP4WNCjbnSvHb7CFGnnlSomIphg67kdl/FX2PDyTy+rTcYV56YPgnNj7H0mum3c
Ew2T0r2bcJH2POnzoSeOTdp+L1mGTYC/AQUZ+S7gNYQCxRGFhiPuCthAygUCyMlE3HqOmfnooJi2
bGFhEpTyRvg/QmXHq0t6STjjsRGpq3wV2jyI72qZBXFSF23EwQsVywV+Q0WVF+Doxl02jvR7xQpv
qVKGlsjIIm3MYFyWXIImzICbb2s6upTIPwqRgBdZO5adXF9iuMLJeiyjBegLaSs5+iSdeWBt9j28
/ChCeccFgiWSneE/PeDcmYSIo9mpfCjxrQoxhaNIVEfovloKe656k/fq+HrW2smy+5TFdQq3jy+V
vGaXWZ3DGELXlleRf97kEM1hoZ+sUkWM7FUsurC7IN0zxggXOPWA73yhY5eEM989oWvUW6EWb195
nMu+8AQhwoqhnzi0VZaPcvG5VVdrR8Aj5xa/klYvCsbtvdBF/4HCNE/ImyAdywityaEH6CtfVVTw
Im2RDKYDPuQ0XJpTNUSmBGJRcvA++xspnWjgwE4dn1K3TcD6egg5mA8p5iKeGP8C6HZVkGBn/Yn+
AbZVH4spFlPyhCEpFZIu536uwXBcKBrSGZA7bLqF07iyTjY+Cyu5fBxzcPGNN9zQqZec1sFn6IaH
X8RsfH08+jxBUjxniYdQyqqB0e+ESu3S2bBJGFspdjwV2kmkpI28Jhlp4xtEcYnMd5WxIgcnVfWD
k5iPOV6O68bBj9esV4Aautoza9ImDabPhgmU2Lyr8MqJzxv3UPR0//L19ILtuAQInLJYWoD01jsx
InPONjW9dHZ/GlmT2Y/L2nxvLt77ib6rqHW/hPEwZpeF8EFD+ItDP7uZCo8cnZgmmKDlHZ/Anim3
kOnK1xlvsiRGQaqQ/Rua+kP14U9YtcxzrKzde/ZN26Icq7XH9FusHjDiEaGkFTb98yw9Gt0y4asB
/JKMIbUzCQeYpt+ftYueai9gAv1jym9fjbEF+myjgoIDhta8fPCRKcWHovqXgDI+Or601OHgqstq
07Xc5lEhpPMF4tZfdZW2I9Zjct5JuNQ/t1Qlwt+ijR05k/Ya7RUU7b+8gCi4SNlNx9XLJQYesx+P
wCcmDQTeUm5P/xvKRyakhWJ8/kKVNjMOwPzTom0mL4j3W95NXx1j5Snq8+u2Fum3jzi0TfVFbNVq
/J+hH3/VrDsEORxGJb3TiC/+GXg7S8nNckQuG5T2WtBQU7pxY0fjyKhiWvhmIlydlHMHCApiH3fq
XSy9c0AN0z4ld0HEopAU9GasACgxO5klytwwheHZLBw7MCWXGTkm2mJ6rxh46HtytlMQlxeaQtNe
ogQ3z0lZO72eW7PabbAc25fs8FtTn/EmPEto40ow33tIIqD8gaRGtzRlyVe2xYEh4jAg5RrCZao4
KsFpI3BqnLdBQ8lwDHyQ+FY6NFKSy2g+KXY25dfm9M2qxJbxnU3+SQLkZdRFAqOyhSdgBg5d4HL8
+4k+B37cZ0HlDdrq18ZvD0OuPfADzLcUDNL07HJXmsRaslhLhFWOiyjgxkql1uSiRfq8HeCAvX+2
+mxVNbREvQ/VyEIRMe1r5js7UsdNi+Nx2S2eKizyWqddW65+eby95BI81k8tKjCtD2tWw5VisVtg
g8p8NkzbzdwHyA3QIIxJUhdWL1oV0PLGla8wYGf0OUGOHJ/bUbMhZcXXY2Z/3ZLaIoDktM3cnB47
wzQgR2juRWiXguYA6iyQgoCUU2SBDOTzNCiA1AQZaM4SD4R3zizRPu40mfx54SAaVEjShHOTnq+w
+H/42HeRaWejujmPVYeRdefJ+CSdurP2giC8TF7U45FMveb03ONH+P1w4HNuw/wRww+k6c5ONiIO
W+kKLEiELkDdb07CzxJXq2F5/RDhvNibM0hYvQo8KVy/QQIaIVCOdhluej96UaWcRTfKe0p2Is2f
ZqaaLg4Zh3VhHPuBhZgA4KYsC5gbjhypDbjUSGe8ICrbluqlbYdxHk3Kr08dhkK4jV6WJZWrT0P3
Z2+i0uyb+Ylzj/LCrtHOheNLbYgHgJbS2DoO3gh6pB/T3p2QVkTOsvQ1dcsDxN27V24b6JCV3cD+
n15wv0LlFLOmn4jswN3FQc5/iIgOsJxLkAKUd+njIlY+KfWYR2H93HRhvCoiFwPtKboGOBlQjQAw
cGWXiDkO2D+sIodkt7CD9MGI9jwfRQ/c5ZVTMIxtk0iX8PKBr7CxKdh11QZVxLXOB3zODk4h3ymE
EyX95d4seQY1LBxww54rpdYk8oCYjSD03enDFPgTGP35eGG7j9x/OGBe6M2iHYH36Pq490gN2Iq2
RkdxvahPCkauNvI/OwmE0DbTBk8Bw+pi1xdzAhOFGKarZV0A5PUhvpx6g86BcfOC8vvkoNlTm6jf
icT3ztrW3XyNhYiiRiPNYCTS/CR56PK+QKVIH7vMiheppyfh7lgVddJJd4jwBybvI2pfDfuPmpQY
q+XshESDTauARsYzlWWPBACDKtmlOFsevMxEfwH2f6grZ/VoawONZO+qKuU4urt//faJGCL9PSk+
gxaZxfENwkivqG6x91Bar2mRkRDeijeqFlpa5B933Ll9TSksap4RE6Svcn4RfSv8VcPIqZbsxV/g
2c9FumgVH+Kdl92LgizZvgCTiv+Z9SLAe2b11W8n91V2SZwzqTEbV6ZBnYXfwEY7WOAPBRckUNtz
bNQpgI3rZfnxpsNmeV/DcqU2782HYfLDmfli6kKv2zbkC75Y9OdHXBLak+ghorMlwhsdU6HUO0e0
9+k5jkYxLCW6SmAF6dmFDmd2PTDpxolVcBzNXIex8kOy0jXkDGMfTVI4rvUKB0sYSl22RIWFM4en
qJQW1+V5tNipEfWIQztP2mUC2kzb6aq/3PdgiBdzovChUf99jeo/G8Hie12emqIoVXJv2k2/wW2n
j0DlRdRze3CeJwsDpV141tZNv2JUp0HfM91xuSbNcHlJu06m/id/4tczbOH4WBEV+m1QoEVN605f
shoFYYGeqwWepPq/INm4FpsWOg565xiXbwOINyxCF5wwf0QcdzsygZqg6nqqr+CKo6iv1MKrCI7l
R3dbo4qyB4/h9ypEBS/X8Du+gDINDOb3DVgw1KmW7j/lSTg8Isi+VFQkBJhtlqpOZtpv64a+MuK1
WiohHynK1O//8WU2d8ykvfz2QTgv5B4VPUZC+hRQjo7qk1FcwwJY1EWEPl+6zOPSis7ciYwHWshd
WsVIhHaXfZAAc4g+OC3OhFnoMs1YIiW01I3RafyZENn49QhciyALawkBA018lliG21TK6V9YLFIo
+bvwjgU9V7h2LibFQ84YanHP7IInk8fhGI949WTUsVI9L/2GU2wGhfW3p4nn9a9CI7Rq4TTjGK+5
yDmVIiYjYc5jV4yOSVYulOwDvrFkJ0AyZn9isaC0Dbh9LH5m9ARj2QW0Iu/yUA6jt1pl/CpwDO8S
BtPt4HNRKdKJ2dooeYhULC3N5PKZ/ShwA2lwtqvvqraBc8f8qKqwCePVjRzkMcZGiriqzgs5dXwP
qcx5ieJHKLEHgq+hkv4na7TAZ02ZWQra/7r4wDLpr/N75sP6zGS3nKMvglrUQMK/K/xGWj0tXq/f
ll0ZGrPrO5tV8ppNdm+e/4TxGS1Y3ID3k2IfcVL9SHYAVY+yKUKIW8uUzLRDOsNFygmqXmLM3ETV
xAmKiwgqasJDtmVZ43lN/91ytNAzAp39wADc77wsDRWI4Ielwrfy44QpBbdcDdRO9P3MuRGAbF0d
TRO3h+f0s9Ythe4NBUEsnjEFty0bTZ2zuIRnx5/MC0suhqvFzdrzUKJo1norcthUlFutyrnagbQ9
lE+YkaYmTZiu5b6Kf0iazw1S8hxI4kzA8zarPmF/IxDyQVteBJ7Okx/Yfj1owWMavV+eI50SCc16
xgdPTo+7hKDjIYghFaJGQRaK7DqohphIDYZuPGCac5bmv5rpWpK30bF7tXJMP7LpS3gFAY9Dh2xC
Qzrme3Nf4KGAb5nWl4CqtpUC05o+AeXHDeei0NjuIo9PmSQ6Bl52FkUei3TgCzoa5cqAcnshGc52
/GZc0bP+SkKZyLUM6aM6EDE3jSaCrzORoby1pkaCJyCBHCMD/lEC2OvbYw+NnBpRT8zn8Do85h5n
SiDURFe2lulWeb9t5eU1veP++nkaRHxW9ucNlTWt7Lsc0gsCm/WyMrdpGET6upMB8FfUBKoxfZUz
KxYGkgQMZiBJ0lRG02BeidZKDAi8XWLZn0Q6q1ej8DIXjPmfv8uHVdPA/vB5OEQTryfPuH9acyLe
PZQ2tYafDy/3cVEdrkf/aCeOBj0rKPz1AHtC/E1hOuSmGZm7Ci/bppvaWjGgJBC2CSbI51Ffu80J
hKioz2pVeg/H925W0COxaMhCsV3BQElCren5S2OtXcc/zW4sO7gIRZHfqc7GCrb3Uls9wb1KKCo1
eownoCrIJtinhUgbBuyY/rXbtWUFZD+L4UyXqsvxlU69xtI/akloMB4ycDfKCBDrKHcov5NwFDsk
75yYtmPBgIhtNQjkRW2LucDkS1Qhbf5ZO3EUldO24H6H6xQatq7h2ZVih+094u/XOp55wfvdW7ex
/RlT9FnvJ2wUywZLERpq5idsV4eXS1tY8iGMgygtbeACxT/ceQylTY/BpA9gGz4V2Vy/brxXmYXy
9ngceFQdyWOVAgzpe8T6Y0r5XfW90Z3L9HuJTjjgnPEy88Oepkp2GyijlkBk5BPywEQ8bsph6rN6
IfU7RXkWCUMLfecLQW8CQKoZWjRvcxvqWyo5rVY23LtZDh2qKxmfBrUhpvCNSG0QM+uqXj6FYZdM
wRnZInXDbdm7THs9CeaQ6bAa5D8Zl/wj4bRUo9h64JNJIdarvtKA7z+dlI2+EoyEVqU9AS9jyBBe
AbYl8Q1gIzQStZjzJgy/8t+dkv4DMJpp3KZzJTmyMYgaKW0q2ujnH0jQE+bp84qie88/rw7w7+b2
kWYkenAvMYc2pGrj0QRc0eg6c3Fy0pSIV880tQ1lb6X2EPRmjdpiIAX8hpJIlI9mXBGCo276mSxb
00EEMwsqRCCcZkuubvJ8OfZBdIb76sI8u9SrXqJiZdJFMfSXZdEvdaF/NREKtGe/wY3GBYuIoQ2+
dm3FOctZTUIg46cXPZ5T2tRAZTTbAYsLp0a9eR6stgZHUDsW3JOuDm1dkB79qGNY29UgM7jI9PoQ
x440IEa3s5wDctxOPHcg74fskNhAbvDNHoNvWjnM2wCmzN1KYRWn41cj8RqOiC0Wjb98nhLRnpE6
rSR5wdpcDWycs7dPj7YUwP4BrQE2N3PU5Opw/hV01PIWKWjLeHAlpBXrLPMly5Y8nyVixGkn2GVM
6vn8OEz+Z8cYHmirrUWsQaDgJlnNgPCCcptvjREcd7FaZlUzmTqOK/sbdTOc9Z8Euheg5nOV5V7W
1AW0GHT9eMZ/ZXa1VypQ6/DkmfJ2Xw/tvkf+C+Ve7RtTJJZfF6UnfK618IPkyCLjNnE5M4AHmird
MXy/9rESQlnSYmomCWDJAIBHHis6pxwC71GfZ7qdx7MHvDHCD9gUn0z3UHucj0cd/ZaHCwVuPc5v
yZSrHESS1dddQHokR2oHKchKCKAqWWJh5vITt17iVNJCSxk19NUjHJqhOvlLZEeQLi1+1CRdnW6A
BJr78Fa9yfWnNAjlGUEpz+z8MRMS364qLcN90lPn4PTpV+50nlDJk4QIetfzsrdtaevPIK0qhq3c
I5OxG4jiQzC5vg6bSNuk9Ongdi7OtjX6JSdhxOinkuZ8n4BH0T+amfurforvgR2k6001oYeaYZMi
OQcU/yHC5tlUJ7ODH8EyuV4o5GNDrBvLIfJWsDSMpO9Au8OkYuHRxEKgO74xUsyj3gSjRl53ufFC
4MThCGgVth0Rjlmis+vS6FwqmFPrMD+IcVRD72kIGHUt9mTt3gkgrhdOmxw6YMEmZdGM6eEAk69Y
S43RAw9PEUGcHkIrQiyx0+TOxgEy1lS74v3ByqRKXv9X5am5shXc8KnR1iUZ5QTIwa/SZdgkS1lL
ZeQpJijg00RNDAFsZMd8rte7zDYysyf8Q3N6SDVizmmTBDM/fyjkpfguwEomvJiycNL6TfD6oiHo
axBr19s6rpqMNrZocw5UKg1K7+J3z10DcIZOAid+EtXlIIGihr07FFtngssJrvNAcn04u+oXS1pJ
sdWwZi9mVjTfbLGPr6AFn0Dp5FgtZfdx0v5NlUBHpEM1qL75CXr3UPndo3XjD6JGhFRx9lT6/YKe
TK8CKUukFCqYos42p6ji8cLgwOX2FFZO8hq3jgL6n403FYe2IAPS+exYfDnXPQMP3XOqJQwK2g28
TeY4MWcbY2yDNPT1K/g2N8Gd33txqj9FMd+qI0grJZ3FBNv65sXBXT9fVD5R0ilc/oIN8GSAPT8G
D1g4ocA+ZVbbVBs3wSUytA7CwF5iCt8TC5dJTpg+TNKuZcmRYrMQ8hzr1SZpV1LYZdmAKfOt2xlZ
mTquj2ZqEG2wb1InQzNAX4JdC3h6fYNRNtRwXq6+PiMh4/G9Ln812vDg4e8P4zABNvseOM/Cs/cj
B/OFjOP7ALi17HmaNvoR1HABMhWXHNe69CEduAhYFako5T9Y/hPBCVv9Nqzajvb3JRos952IXm1s
uG7SzyhKL4/BQ1H9DQgDd6f1TSQy05MKrhHpQFqp3+8A/XixDpzsmBgq/NBWgwyHQu0Uh7CZY1Sr
LudrlK45qWx4265ELzxszYypmPqeqsfjkeZInV7kF0Rn0+JQwbyFAMzevgnYCDqPJOBt0OHH+jgf
6OiJ3brudMVyKPTlO2CQVNASeQSrfH5hgS9NdSw8OX7VqG/gfGNWk8047gWVLAGZDusaxZtVQfT5
pNM+u59luvHVA9ZF4OTYfRuLI7Khv3qPbN9sSD75MH0uysoQYQhgHG7QdmjA1ArYMufskYyv86Ce
7bRnNpJzIEJntyucJ3i190kQ/sN3wLEnH8VGgJ+QbfR3l3NqvcswxoxOEfBcXNEn30D8qRf7PH9Q
vs+l3W70K+HsbNE9xaGa3LoFY7AFOT0wlAwtbufy/6PJdZbKAd0FZDLew8eEbp0hLOHv6lJoM+M8
/lBEd1AmipCh6qbRfR70bZoxT+v8jtSoDfhEEILBdCkamTHu8GcoDgNIgzKLKeRbN2qlUoz9/vyW
HWYBVAn5aYQbOzW7WEgj50XJMUhQxgRvsO7/HQwCRCpliYjzMa9JvPsT36GG95sLUxV/g1DVtXJe
jtx9aEPOU8+bv9ox8bivzzYgMjHu+W/QMU5u9+7YXkPOUzaBCySM8m/deMaAavWM8pojagbic/WB
ZkQhaOiFtLWctfrftf3WiN+WHgskYZq2duKg4hX159nyXPeZCxcPMlvH4CmkHVzs57hmi1dSbZJC
xRt148UlEJXwqHGVhVtAIdpeEwpMeHsKevBD91lyIvpZ96B5WtScxK7amw/5qOsUXjdGnOZToEkp
51Eb+UxigjAqU7VounYZaZcSI09pLR11ar+6fBskZzxi/7s2yRS47CXc61ZkiXEHB6g7tM9JESEN
V3cPbTVc9tk7voJrX7JW6DuHbChbdU2moKicFsRHF0CKaqzDTfVdlGtDEzNbCbslslufeET50CaO
QkdGyDS8017phEtJ2ppPt+kUTlZIrteBMsbuoGq0mBbSQpb0i3txSfjnwbYVa81yYL9POWjnMeOb
Tl3muLW0tzqWc11VvXvAIlZx1gzNvhc1VcuN1Bk18ypRZ/FRInNrdomB9WVZN4cgDfdDqoLbVHSy
5Kut7shOcTRIWIVRIWGfogBK3tMUl1XCEtfIDwiQGfLly7BV2JxWgCDmEF52TuBmmZQxt5Z49Wum
a8YPEgOmPlB1HiimTa8EInLLY3zhLaA+3Eqz2Q1yeoHkMNJZysaaj23doUFejTPGoyz3mQeziEpk
bTyrikSEOO3JTCWfPtlAZRez/nCX+wOma/rt8Vn8+JmfMVxMimCBGkZiLhFDXKTFhwRLjF4P0ERd
f2wTy/TDydsfZo9pTY7jGdR3bSWZ5Fk0KXJX2puXanbRuR59OGlwZLjiEUwQzbKazbtkAsvj0vDB
ycXZw+aMmCf1/Q+6frWfmpIprC1r6tq07hQKdCl6RirDGI4wXOHrKXny1H7DBkfwdP437eT0r/yU
u7jTH8b6dMp6aYl9tpR4c8mcHOWYYrSV+VgqPzRAeVmvYySP+Xz/8lXLUQaZzqKkhuVs0welPUz+
mkyUiWRyZmp9A9rNnE2+4NkZu7yMkS/m3qFPWeY/cOPamRh2xve+mTz5Xcvbg0zVv1Y3qwZx3utb
kfZHUTvkgfx+dOY5X9ZVMvBhJXcFr/Cn1Ni4kg8HN8EdbRbxQYOXM0+flc/F1BVrAAV86PGGjIuZ
ppR6sSib8EdkmgAoVNjz99yPPzZtRVW53fvTzItlCDM9H3hqwP4zQi784P/BwBJ3mVxyPe0Nkukb
HFhJ/+Isc8P6spp7ZbYlkXRPUd7CTrXqGjF2SDj2gtMEoq9f2vWFVaRyJ496UKbhaWMwkZAZ+Ypc
QYfIdlRan63FdfpTuJ2C7SaKxEWxGk5iJJ3dzczIpbaB/4QS31btLzOcJKOHtkn2yuzjNmqEqgWc
QgZAVkD86RieM4BvEwOOrWPIwt7sEMaXUiKFANSI0J3H5zgYVTic68lJE3sZgD1sDeGpAph7Q0Rs
/vfhKIqjzFSk6tFopCi0HDPsYVlj3NUjgRTeTHlvrHhfyG5w+EYX2BYid1OJSbVpMtEcRf2NVvVl
0fG2+bnE4sGLfSXkVtE2bLcE6JqIVubZ8S6f952oecWOJsA0dH2qlWXLYlEXSBFvLVE9llqLfk9e
wglU2nesAYqDcti4oJGUPY0YfMB+YhKhMTC2ifyefeHQai5JnyCQ+rWRbRn5zN1jmt74jC9/PM9c
FpHtFv157kNyklGVC4H8oTronv1COwysgYN6XBsK7ZhOv/7n83Wrxic3U/nbfP9CfWNY2Z/zlrj7
XE7Zf2tDgNtVpBZPdF8PsO7bwi6l5fUIGQ4hfjY9G1jcQjapwub+AmOGHwIElIohDx6AaAEr6JEa
/Z7+zp0FETfQH/vSj41ZJz2gTTfWftPa5tj+BeSp4B/4AaW5nSe+N6oBzZLKk4YHlQXWAIWssiNv
f2Ddq5z8Xhb0a6BGasPFm8s/dFQmioSuGk43ICb2osYZVari/EpGV7p5oswmhjI/oY1CPm5ww+e7
pZwUYnzsGmZ2Si5eAkUC4rRJOK5utKuj+wRWoNlF0Ckk/y9WXj/tsYfAQeWGo7lLHAmEewDMwG1u
JbbtTgFC521/rwp+LWl8iQ7sEQrRP4rGgjUuB13kupQ/NJUloOawdhqlhZ5C8XmdEUB8EwX2XaQU
4ZEV+EqJkE7vQU5XEvVnvsG/iY4Hvuy3X5yY6CiHbpZn1OFrItWqW9wY8ZFlB52txjhMprwE7Yi3
Zsf+k81i90qoL084niXVRcwibm6JvtzFPxl38dffEwPGdWb/EAhkz9iTcDtk2WRHlyGjy+e2GzP9
xbVNifE0y6vZIo4TWGDtXnBT/tacloDCrENxdE7fkaa+qzfOo51k+wu7okLtBstB4PzM/rU3KaVz
K0BSrHRWFgKEAU5nJGC6jqUXso5gtF8JpF8ecBIZWmRC8Zus7Pfi3GbrY3muQKrqyafd7xqlKsWE
vvg/n4Mw9s7I5zTcevXol8mMH9z1f/RG2VsW9anmgDth4UppVXXuKEsrDz68oovISkIXI7997RTh
X4bMaHEV+H3KL216amqxP6iT64nEEyKQaEflsquS35t3GyjbhVHWfoLXxAJOMQ1mo7wcOXvyJlTw
fb4dhRWSSqQh/Wgn0sXUllij1Z1gIhM4wslC0c0a7s9lYZkqUXg9HjUDvwvKFPKPPLhZpuEx+xPS
/SeYkdJaJ8eWu3ZpUFuKd4x0vaAoacYo+dNA0F+ySNOCQbxu6hPZrPZ/Uw2ZGRQrMlrt30XMrwmo
pyiu5mN/tJ8alnzwK3Zid4Q36avY3l0O+7T3rRRezY+HAtgV9cyoOD8uyKbqnBZjXBEvHXgsMbSx
+Sywi6TKfQu7At4u8ZraY2xVdUfcy2tSdicPyL0GDTunT90TuUc3JW3Zf1xinEBbRVDSmv1lNa/k
DIvx6fagoajdBERbyg9LX4IQ6ZkwgSDcbHj74zw3HG+MNq4NO/pYr9XKVvCg7e9NrFb+/48OFZ2k
pjszf7r8ig8rLuIZcEzJyqjvjGLoEhEH3l2cVotFuaHPRQPfagvxUzKnzeT6kIfr1fzs438jZDyr
WaofauX1frG8hzcG+1NJ4/TQs1U62hO+9/OGDwb37lzd6SZby0X3tYEMvTygp20cBY0oTqxuUlm4
CXT8pF9+4TERxqIGdxUfjdSIrN2vRxWMTppy34GkKptUJtj/C+MElwVRB9fb726zqaPyvBpZajgY
01QHYcO90YD5S8GrrEC2eNREZP9Igoov0GD4NpYtgRj5vZAXZfA9VNCfa6jCUlgDySUEIPM4hgO4
ozdsWXGrJcxLUk6ykYAUkpfZ+3/6crfBf339/6EWYlsb04Wx6UCEwb4id/c/p5gWp5FkTiosoFnY
wfnc/M0IdhL17oEm4zTDu/EVUp3wdhoMupxVLKuJgRkLMFaqYGdtnt0eTzDW5I/Y6rRVj/Cru5Ce
xdLJHCSqK9o11p/u3qy4T6ojza/uzej2ERCa98Jsxn/x+JzLOteOSmBM7fk/4JeOgqbxS13zb1mk
e7xf6uX5O4nqb7yOeXmchbH6s7+eR7ozlYqiz/hdcJM+8zojVyQfOO7HuA+Jf9pGqs2AsWmE7sJF
sraT29ZO+aMcB7GgGefEV8STbiVkBMnAkjoUaBNnNbLovo3fK7i/rzvj8BN2jyBruHd6lw1C7psT
XZs00a0e902iM/Vxe9nxKHBc9jN96ja0YCluy9DwRxAikzqGDZoGG/FxQytWHMhJmJ7GfOMtraBl
Tuz/X1azSPcPb9UnxN4pIFrrYrV+FAM5p7xLXVNvfw7HaWBrHLKHLjrKUV+oRRBZ3XHOUVGQszkq
NOgeYWYubWq5+bon5PVAjr9pUJJZSIuBwsEtDraSZ3vxUUQ4j/SiBhpmOkTiYQbnhllvnCiWAcSE
dmxRGxFdDTNDgFtY6jb7LtFQJOxTiWS1rITC/ey7zHmV1j+CuAlp/s8SZ/b7XcX3JcNkRsWnHgzC
i9iEz8Ge4c5i3nooIzFcMwu5qpwbHEcW6nsGnq6ITWd2sewZdvBiHmpNDaWYWaTRJMs6NoRXjgjC
orlgS2XrZBpNytUW7xHacm7+TDGD3cUIfNYY9QQWlJvgD1pmxwjmSzgJUyFRD9HsSVUkHIMm/W2h
M2FgkWfuapCyw9UBeUnnvpyvwvIxtxHWupbbyhKisz7KXuIlTYXL1jbC0e/ADKmOSl0Ygzx5grQw
CnejUaISsK9fPPU7RXFQ+0jqvzGqwuXTqK+0tDi2bHEg304n5XSNxI/K3Aaxxcyhsaqs4qMaLA98
jpQCSbGoHRwdpofwesEiTZHziGkfZ25y6mdrbH7DXBA9THGJa6dvFJBJOHG8foEMuNebExluhRGg
uGbH2oBHH1uywVcoPTjsDv8okRTGEwlIj69wgpIIKMnqn281Le2gYfu5+fopDt+yJU3gJZxPPaCY
Zgm+NU73GJrjHwwtXPh6Re3/tPK4QWuCk/Ew2lpQVvoK05J09qqO7Qoanb6hR0ivhRHy3LwxZjqm
QRGGd3Dx62qEz0/YhsjbCG9qW7h544Z/3fOr+WRNWcB4P/DWx/7bhWqTEwSLx9+ItCUSsraOEpdd
xDo6qP83hdjauOICzfBbqVh9tApyaCxBexQCpiJEHKB5Gaze4iN/4+v6osOYoAD91BuJWAZKt2mQ
HwJjNNRNB/KbUmPM86Z7lLTs8UhsmjcCw/jUJNCpapJb7H+NhQNzQYIBENjjpOYZATKEZS+hGnpM
Wb0F/zfqKadH64lksEqLFvZ84YV2OlB/Wem++m2XeWXHQdpIHeTUo26wLlTTwKJLhpZFAG+a5/B/
vp4csUBSPKIFsBiCCkL5QxdgNHkzy5tIbx6Gn7Y3UU5oS41vOWX6DPsrRl7ZMtTRxkwval3rGGte
3/QaiS/hejRDywxVQGkilcaIUE1MN/IUa5a++ZwxpV7LXtu8mcB39yzzdkmOoEvf5+JAmU8yzLS/
ribavWqIiaKbJ9yjkmBGn6NSAHQ03DWvrVXpCvGhjxmNLDELmVpdzSIIt1w4OMO+9FRjyUZlx1Qx
LDr3CJTb9zyBQuSDDLOiZwuTLvUAN3z3mE8/h6vC60IRVcEa7nM35rmEqX8uMaTNrWVEwKUF6RKD
ReKU8MhyX9RiBHy6yXmfjgJPAKGtXCQc26R5Bsjoa4yVmiXRM35CM317im3EnaNZGpNX+JY7Kz7v
2TbXsZOCDiRZp5NUI1nXoBsxwzFhj58cNkeK3Z+x8Vn6Fw04Xjp9Fkp7cpmv2auM3rDQFheZUuIY
0x9+C4LTM2HJwGbygQvBCv0FVWizEDWRa6pop0S+qY068ydHTPeBTPZ4oreF7QL9AT6eNPztDitf
pbVi9hHyJyaM4BOqDV20fsLm4bZRwsYuCTqMedeC7TLfeCTfOdTxP846ImATpMiMVrSbVm0QNa+s
Uy6/F2ZTmghYTKMGQcwrF08xajH0LTFIntQSUP/Tvb8GXGW5mzdJ862nviHHzUfMQjckt5sAXzce
L9px6SrfVZ3/qF68By5DrV0k1PRa8w7Bb/K/kBFtD/DYWlwKzseIKY4iMU51GJWgWohRJY7EUmf8
eUia209B8lLplG3NAIYKCxltkinLOYinhUoCg2sNfx3gwzVIdgQhM4CeNoEXLziT43E2220M07Q7
mXHmpQ4x7jPSepvoawDWIQWxNO6CCN+8X3sDWypla15dsiEo74SivHLGnsVjXJ+94QrfjmT15K8j
18NMQAaGXycYGO0jLaEXdWkqwYtrt/W/Y9RdSqG/6OCFDXxIxE4kQ/tIRiQ5o9a/kQCRCIe70xnj
0GOWaXV7P0qP3uulaj2aqxZoULH0IpwLPEC+cFE3wFbouq77sLh117r4CASRkTP4cMCB+B4WBw/3
IWHkSkMf52zHw/n5F0V3r3mGCL2OWEVlInT/5uIL4bZ/rXHxdkUC8SZ1P4dtFDPJDOUdZiR7/oM4
ctiiyin2BDJjDXFvNOLlTVaOM2a+1wVWp8HT8WoU1oFACT+EI6nDKDJRzpR8+wMUBKKPe/wvvzlU
jjDsPqRYQ77Fqg3dZE72zMWG71PqMakqZKyTrDo1sxeD1SJPpKAnXP74yYuhoME3CXxooR/SeT8Y
2z8bdfCXlz2vsjc90uGMX9tH68SPoVhDM3VmcH5SePa6acUkuKl9b0+XxeIs0fiQW6hNwJ5N3STy
D8jAoErRK5q/CX1MAXXn42ye4vUJpuDbED72vYoRietPGWQ5mEbNH3UrCUSX0nBVNukHp/Vfj6lQ
4qYsdLfXaxu4CLDJQjf7tKBUH/7M2rNCmG/6Hk+mwumQljtW09u/zIF7N8GwQqnT1wC1zyG0Se2M
TG/vlyJf/4SYiajIjabi4xdbHcUptIQfkZW7CafFONFSkUXjYUYoa+rvxJWXlT932r9q5A7H7YfO
8eR8QJbOabkmCoaru35qIU81u4x3J8mGcBXJtRVX+lXJy7LvQ71EdBgPmr4lKbQz5PWE7A9iyrr5
PlL6H4N5dvzQf2alILK10bosl3zG0rSB1b6Me/jqX7ZG72U8YSuc5DQ7+IqBWMi7AFAJ4+uP6Den
3rEmtKDnlCV3/oaoE6/n6FggdYkijsrBHi1BIMpwE9NRUJEYJ6MbaDu5HvuUa/1eJwB6NjjYyifk
lggMJ51cW+5qDqnSBlh+dgby9frWlFQuBZVwWCBCjkD+9gIQcYF/JfNLHNRecphnRejc7aYpJLTL
JgAf80LfzXN4mKCeXM0g7u8r3gDUBlJpny9GKMyuRT+oCBf3wuivo6A6AAtLerDVVtJK14TVb43H
RwcM5KtL1bjGO1VMggfPU/SKunjz8Q/X1ngtc4+yyJRdRhe3lH+83rgRMrBbVHrK6u/HnvhuQKaw
lFUW3G8PgRqG5H1T/T/V4bdqEvdhO4UOJwiKFIWVl2N2PaDDkFWD3/h89+ft2upzNwTfeKd85NKg
7UtJbMrFQ+VNrcGS6KFfmYAKC+9mfxADBZ95LYzQNu1fbQ7D//gJvCnkHqB8fZUU0Xksk/zhDqSl
iDjgtmW3Ce2Q4GrZqIJufRudCI+hs2C8kFz6W4tgG1hOlOblI4ZBVw4VdnVDQ2+yUx0lFjI/hcli
pCBA2X9XA1RNkMYB1ue1oMxLGPeF9TExCVnk7DXw6KEUMT8sjdbvD/bjkBmLvg4GCFEjAus4kO4F
OyDOtKqoopP/118wz6yJZEhptaJFhloHCSgbsvjupdeCY9qUDt31LO4zbi65HjAWiGatV1qcBc3W
uaXMlFv+o5dHPwmniZVSVjInOs06kVKuZCHtE3+ycmFmM0v3flRqzQ7ebZ3mIjsKlCAAQNZr8wvw
OCLnH9Qd68V02Aw1/ISCWxXW/Rp+V2nk+4+tWzDbhyvsiW06Wn58fw42UBDjy40aJ9d2oPAfE/59
B7Z7bqUhhupqn4BxoGeJGP+Ye7FRsbXhS5vQeLIVDlvJM/wDEHJGHq/0j1d0sNjojV/VSQ47xPJc
1e6RLEaECb1F8NhWl/BIly/6nOU2a5rAYI+w5UuRZQ6mmPtq8GQMz/fCNejqsKJOjS+RFObsCajA
9F+BnHE2ZgaKWm2NGOBBipSXSyX0gerbEBaPBlrpebczhKyT2yrOfvnu8HxJVvzGssPvwWYwccO7
Dm22jqIjEYYh6hKVzHLQ32LHVxRVY7NvWr+xyqpUEduD4gU4SgR81NkOexqtsig+yXVU7KcBH+9o
TYk3+QeKcZ1817IoYUKGV7noWM3HGz4ttqHkqPoVdV8w16pJ6zlA7URawDCd0XuWNUV4LDv63M15
eUYftnWN32uUtkv14UW9vLIayNljvXQfk2RvMld0YbHPc2YDZttF0srpoUxW521A9KHOlPhVB/Z8
ydKGVHxgnKIVw9Z37qX5KTzTlw8yMfCceVYI6K4hp8fab1/ld11OqbSZEWtQwAba3dO8I8lzZQKB
2tpouwYABOvdAWWPmpGgEV0b0j2dDz/+LcKt9fIz0gIQ9IVaa5Uu/3yMsQOeY2siXnJ32lDK6E3r
DGvviOt3dFGrxqe0w/JU8SF9rTBA9pkUIe3ZFk7N7UKxrVKBWHJB8jZ9ly940rnSTmT+UpMd2E32
yy/LXM9YZw6p+QGJrKxDIdx4M/clrN3poC9+aa+vmGMZMkyoePZdPJGF50qaGtVLrO3RT4a3F5mO
q2qTbuqcnQ7drtejIFkTnV9iJmzbA0cERlfdfy3EnmR2C6TffFpa+Gqi33F95nRICUHwRjCMujE5
NPtWJBCyeOHsN0e/A+aW8fvZxkGA/OllJ+vvMMisWkRfPeO/xnDtYvUkG8uox+Ey4mCB6EqBYcEV
ZyutBY+oTdJnJmZLikG8tlkJ7YN+5716ftW6ebf1Enq+agSJItBt7E4jaMZnTktt7PvP2WQG+zpg
OEvfjCe9ScfAO/qYOumDtzIxgyiSeDsfg8yZFpXGpEv5kkGbiwzzGMo9ba3wH/ZenLmSbHz4g3h1
30PiZqL9+Y1H4oUY0RbPuvmcPABJdmRZ01wp2NPHxqItNo5+/HKuz1zq2sYEQt04+rCLneY6qMmf
i2X/LoWF7rs8yGiuDQQ1vswKfm0xjMud4DflD61BPV03B8pz3fg8CxW3EODYmB+CECkfbIuAGK2K
gcwD/1j4FzWPyotEx8X9AKBcwxiKgsh+dDvGVnPYPHNiMWFqFlGmJmQhQ3p2iO/7TFyL0nfCJFO9
bDvoHh2UPbsLFUU642pIPEHzBItJ254zqPdQwwptI9CFQ6GXarCAaQITc8sJ5kXFDVBB0SZYZZhL
STwOqXlKgc2dedWY3FCbZCi3WtRl8mfiCu+/Vpg5gpfnSQfKViiE2EhC6grLCyQDMUf/oM3Z6FsH
H44FoEanNkQ9DTJ6flonmZwnyQpBTxrFk0uirt4vQklpUO5x74eWjhCIV2Dxr58Vy/QDrpgCPN78
DRswGdpsafLVfDGj+GOLQDF3Iy+j/eou/8vDmqnMyB9l8ro2G7nOSdZO8dTrtrarJbrcW1m7Zi+w
35lCyd9RgzYfIPW/JAc5/biVMMbkLBex0Mk3GITqn3wv0jw3vDhe9zf4jTEplFk2fPXAnsvlmjtc
dO67t1nG/CQTZzl/JFdkP5+2qP/sLrywVG+tt1Y6Ea5tmSSgImwsUivUyMAY75hg/vv66gYBgNlN
BoRPTJWNziVAicB+EcAEIU78XEKiKZatYpH/tcHMO+ujmuZCcxJFHjW9AthxWmbksKvSfJvLoRpG
JMrWYgweFQOUnsF9FJsXIZgqLA3TNBtxa4Ew5Ko57rXWAeubkT2V/NQ0F5S1+9zQpUkn/SvW6N5M
EMmElLFUi93S6ja2GRJ3EvUG4nbKMuj/ZajZ+uhebtaKP3XpTuM3VMhtdU3YmyWz1TfciflhZHtR
m6cP5+obKPLoxty+nWu+OFiOMdLzpRLvIVcmaV3RbmH445eUEdTCvxImMS+XrWOYZSMFCJGCuiYb
agn0hs96+mnq95BkbhcU0haCE699VJJeVLYagYnAr4+jqhJvtHauMwefO44LgRplMd9CF0MKBFzB
KV9OY20tSD2r/dH8jyiP5MGqxjxCLAXhE1c5KNNxFaqXPu2iy4fnjG1AETcdsBr6CDMDPjKRuUhv
dPW26b+9xYwHqbLNQpwNT7M/142cNMFShvbnoFnSyBrQZJp8e4Y/WvI67xj4WUmco0TOikSHMHM5
CRy1HPU2vtZf/MjtLit6OW5AST4ytEObipU36rKIGULgDePEBeJhGwugc6+3GT8o4BwxpJjj8sLP
sp/TmHUIQrYedqoe7vbvbXtSMexMkHoprp2r0dSjtGsoQFIz2MAgkWSYLvktfDCV7YsBnK654Nwg
QiVtv6h0WXQOaUyfZbXwIlooTFY4xQDchJwZrvP1W/Qu4wMqqollnQ+eHQ6OcCTdYNd6heqD+ABy
dS9pIzlr2fPfTfAS7Jl9/gs9ZNppKfw4kUIKYiVZviIPUemgRLqNhKvV10vB2Gnwp/m0D5Xn11fN
y8YAGPeM0g2NKksmmMJHesfUDmPTz1MZn5IxJB0fpX+Ec0520qClkDYEx3HwAHOHK4dwZexMT9iW
7JC0ZexDGFEDcnHFbjZqIsi6uUQvNbK4TPGPf8fTfQAmlS52MzcB3C3udeZp3Nf5Q99rKNIjkBfR
LD5Uho04O46OpS9ZGS3HDxy5i8JIjg2Al5KtSi9enJBIkxIylpaD7n1rI2wJ2bBn4xHWO9UXJJkq
X/t4SiYpby/n+RdJV3fAcQv49rJVmkDoq/AQgJY1h1nq8dy4LiURzImV77Jx9rMopuWgg8d/TVw+
+OVQ8V6UzBN3KViHs+5q4eGpZov0IBFydFymNSVfWSkXnwtmGNIQusAPinn+fEh627zNkUfWPqjI
wwYUQBZgnNrHecQK8kGfX7BGG/PY6oLLa95JyIpJug+ras3yIjb6gXtSfAvXbaWP3NgXeX36zddV
FRfP2vfmAiqjquwPn/4d5F7tPdEnRtXQKrIOhSyTJcq68aLU8SDpSNwkyUJXHp1+aw4OLVj2/tUh
SsOYXaU3uu9yTrBs86zjxeKtUQ9xSdQ8qPxaqZ05fEO6ltmjodF1AHOGSaboR9H3W1+M7RPpPplb
wX3byyAc1XeIIAlcYH6wPOk8gTvYSdN4VuL6PITaEoyeXr/NcRLmrwZlT/Za3/8lgvGfTfzxCN4l
/WTTvhQnH5PmRutX0kOa+qAIfJztDV6RvT83PXaDJID4QeW/QnX/IuzD5fFWCu9k7ivJeDfTp4R9
1T8P2x4W+3t8jbertClcHW4+3s/hOSQqqPas6ZoPKAQJXYzIBFUH74y5NkElqXjehFvJBRH/Y/lV
u/SYZO2faXzFH5aX2zoJqumUbf01ByCias8M0d5KmdLNzMQd2mle4mDnrqNP0fBhfZkobM5bOaul
+arSoJ7cCVcwiZ1KkM09XXfbR+8jGxIErhPd1dTQlAHBwpFAJD0n3f5yfRhz+U6KYFXbJlZugxQS
3ADWdiwkFTh4DyltDzWf6DEnaVWvcS490hmpc7WXTN/cVXXkeQhW6oYRfT2gs/c5xN3NOnxzFMrq
5rLF5fRh0NvW52rmB434PNpy3uKYxVnH53qo5M5x56o5br4VeAW2F9xUcMP/fFzP09oXEVjoHXZ+
73+0rziZBtHYb3DJbPaspXIL2MCDcYLY0JUzZD+aELcLRpsxGg0jc5wnYBkmEVoc81cGpXLnY7Sh
IvEVomIWkZGrR3kgzxiPZhd2ntVHPgkxSEzHF7sjHcJ38lbVc1woKFqpIK+rpPqUrDtjKpsZkO0w
7OIgRn0A2Nr170km6VPZOCfAAvwDWwscMvHxbDUSs88uZVPsqsxO+dEkazz0XUsuP1N5KUkLV/xB
aPyqWxFPK1xGfju58h/qHX+u6ZXyN4EVZrz4Avf/Ho6kLvMfpjFKKoSjs33xKaXtJqXuX5odWkHh
yZijbDX3QR086KGpZgDDa3QwqtEp9Y81/+TDc91su/75GFJ0ixGeHyH7v3S/JLeWubX/bljKfLcg
1rWb1ZzdTZUvPeeUN52q1LyasBwsc2pfK7hqpkw07qwlY7YgWsa9mnB8LWif1SPR3YXTvPuxsOfp
tUC6YD40P6XrYUAhRtLjNtHGl0uhO2jlkBfCbk2JRY1lEUj8Bd6NqjDUbfyAgLAw/9wddRVUEO8e
E0HLmxzykS3HblJKkfI080sMIB5JftzGWfQOwVMhQ/LUCzKfLsax0kj39KOsE5gaBFFuTPmSOfZx
/2X+crNv2HvtlOicf9jsN3nzgp8sesF2L70R5sNH+2oRkna7JmekKNLWBDvmnU5U3B7bpU/LMxE+
G/7nGIJDovCn2tJz1tYBXtknzIXDYxgCzk3xDDDVm8vLm9syKs7FpRQmsQEguheHjiLzGNFv/OKk
YzU2Y2j2IO5UGnoC1imLzzYKksPZcxXWnK9RQri8KwSkbIkY9UkObkqoc8BwxYBGLaTWLOS8ofex
Pg8gHCzVIn4WBUm0hLGOVv+xf5NypyUni5AIx4OILVTcxJUsQgwrDqMeUhwUsmCs93eOD1ZDdamD
ZwUdhrAP1F8P2BdSGutajvXXfEFchU2vcJ87k+IR736yjPS1rPX99w1UtxapasvtK1oVJAmVWIdX
pcyuS6STdJ1o1BPvB12DrtoCOg9rFV6yBH+oJaC322O/Smddbt5/RZCIzIxBC+4e9r+scQQ2gWhS
QOS5LIA7Y+mYo6HNxTCb1VRQ4C51/pIBlTBoV9EBwVC+R3wMao3JBpildYspOhQZUFwegc6Y+t53
URQRk8iVnVuuMdcBIoIPbDwDZhdRKvbgLJ93KzP6id/tmw/X0D5p25eJenbGnSQal0oWS1MOkmgm
GDOkkdpDJq9uA8LJtVzcspN3prUEDE+n4TRM0If3yHSt9wCYoNPcZHz3VtO/xgWkqNj1s/oapu1c
8Vlc6lEvTsweXvlB7DmKqPkdxh/HYCY/309a4/stquVYZPxEkS+nh9jB0nf73UKADzwEyX+mwVB7
4hxo3s7fpgPnTS+sDZ69ckh8NKMlpSauI+pvqC8Yt57iDQ61qCN6CpWdRdZvUo4Lat8KU1I40WP/
7R4hae4WsaQ5rTmRk3bK5eYMDpHs2XhPv7RgCZxagy6NB8TlKIH5xcXmEGYYbw455Z6ic6dGATKq
A8aSrfVVKWFxh+K/h1RUqL22l4dyszJtOuZQjsxw4gFvFGX2CCIuELvvXb/+gEwld1hNwQ+eG+ut
oeKMuxqbV+APirH+sR3IwLRpF6vrvreIn4KxgxBM1MjeqKJ0QS3RUmzo1rz04iWr4oy8E+oBUmKs
nc2A5nttNTCy7YSc0XoAAXWLF4F1uT5IBvkbUNqbSHUa/wGyS+K/ylFW1Ie6/6zEz6aCwr6nK5Iw
Mll1qzuJm9LDoR4GPTNLh0ubZoJ5fTzcTAKTfA9m9Q6hn8RVgOQmPH7YlW6E4RpxBvbqtxCQgrJr
UA2ahnvKnE7cJxsco3TdOklPBga5KaWzpFdcidU7XeZ8zZBRLuc4F3ZZQ6f9LE4avaBsDwvJiqlH
54hVO/hyzdQZJpr0MjRs1+hS9VmRx/QOkK7UA45bjLKGqes6XPPQ8bOJSWLQVbNFsXGmHIQBb74s
7pqGCSUeFAWn2+m2rTtRRcO761jL6kfin8q3tajup+UwtoKOjJ7B21O8mX13Oy7wko+s1nZ+CoUP
GHtK9A6XQ8e1ayXc7pPx4+p46dOBE/Mn0UeNM9foY/zFD8AspsUY2ycConCWIBiTOfwR0e9PYAVp
S1wB9rSmz+1toTXrBV0t8eL+AMEe/Jpx5olxkO4jv/qHkPJrg4ZldMaw0TSp3MOGy4LPkO5vU6vy
i+S6YNKvmXVV3oR48eAeDuX9YkZnXg2Q4x/V6GVUSmA2hJSBUcVsoABKZUMIJJYwGKcteXIPmLoe
r1s4hrq8bwC28lcFoW0twtgS0I/t90GSPAd5mJQVYlFpWqX05EHj+LGLABLIEKLBEavlClJmO7jg
YhMd05NZKUycSd8kJE5YLfQZZhDUm2RaBFPCdv/YXTCVaghT6gopadQCKj9QJGbqwICcpETiBld0
uc9unlbAtym7l2HLM5OvI4grePdKz4D79FpUtqRL0PIyIx4s8Yc31MSu/BS1RJNLr7W5UPzeCDFW
R9g4xJ8a/j4op1sATi5rn6nbvxKG9gFYVodPYy2xlbkgAbPPYY0lV9EgyksRkmYvtL7i1mO9unkx
8V09EqHKHbS2aLTsJbjMTE2ROvt12+L6o7dq90NIhqGhHflVu1PC0q1iOJTUfg6hjUIUyce6de6t
RXnMDdyX3Twqis8HUlMwX8DW4svatMMLsqH9aWcqS6GfTKAMPlGiWU7uC6gcPrZYEo/9VHE7TbGF
/KmN62ttfEjbC7hb2EcYqn1+p/2TJiqPm9vrx4Ir5C587hMFM8Q+8RMp03EvVESWB5s15IShuBuO
muA7KeNO4ekVMZbFWi6zAnhJFwzA/O2ouvS8sJFDsESo76+jyxuIbGnQ2rq2SvMyxwRTn81WJzLw
dqLcAfVro/k7WffUND4qsUVtcWNTtlXauyTQclnpPG/6T7b6WNaKSnnsBxFCBqFyQEmjGloejFaj
1Y2in5CPMnDkl8d/4/behP2hSnak2xJw6wDBix3vW4fiAnjFRL+/c7xKN7+OBdoc78HCSecHmKsh
g41HknICNI1rav12w4E/D+AHbtKXMJzQSZsydB4CGokdf5EFmhypceVTtl+NoKUznmDIrWv4LfVK
iCgr2PLRtcyp22OABXMJZNHzJYkgxLlIwWKXNNs8hBw/zNT8XDM8ep+e5vc+pVZ63S9FE18H5jG+
jBXvkCP70G58GCnjSUzmXzl6zHKYZHRFsX+wB5o/kUwdX9wwKI1eWq5NrZ1DDWQrwqEPB0nHu3QI
oKarFuGY+ptPsX2W2tmd4gnzeiiUZ/femPLoKyodbgI+qmBi42SDhu2HtGewuMPQeL/pbYHT1BcS
uP8+oMm87RuNKgYngdnm/MNoNjfWxYp7KzwAUHanau1xhfs1qlZld6o8dKr/8r/OO5Eaj6nrFdk/
PtDHl6vfp2cezw5Qml0a6qmaw3f2VqvbBxMhJvLMki9ce6QWd0d0e7klc8WpiSIunVCShwae7LVr
t2oXuFZwf2ww643Ok21iG4djNgTqEeLZtntuaFrb+mrgbn/0UWeKEebN3WeMcCmXJ3OHDcDdpiNX
zXErxNnPQa6Tt1xZs1vTkqQ/834HEpU3YDCYTjjNUzcelMxHlHTNDwZcNyJnlSXE5vPykVLmnhrJ
CLoeMFyE8ctia3YSTVbHW+YrIz4I7WI7oO5Dtb5y0WAXFETP+qZ+UwGfloU6qcQzX3uTxWUSyID8
iLTBc28RWIbgsM6bWWhFXJpD62YAIRGLiXb8pXlL/jPvWntBz4PHqRgwM6nojjFyGDpBz/Ig2+MP
34qVqcXsnufsRDK7Tz98ZUjeNaWQ9dWmFseQ9uFzRdUynVDtf3Elj8FMipQdW6Cnmqv9eWK+cH+c
O0Yef08FwS+mrEX8UQY3i71+mgieXPyevzsdpYQYjfbRsACnp8Aiitq1b9x8giISgzlrMo58Q65V
HjDlW+HPuDrPZGQZpyt/S+MhT2PKklL+y0qbHZ6nOlNAR8YJuO1tL9RS1Nu57GDsu4N4NApW1BuH
D2pHcbxwmQWPnktHdQBUaNKV2j4ZKcwX8vOucVfgAeKUziWwljiYbpirIqusg5YVNIo0mDxxazIs
OWwM+0PHG7Vi50RFJ4MFuR2UwRGjM20uBMCKCde0jeSjIdcTr0wKXb80K6Gech7po0Eg6lUAanP6
XCrFWUpAoFNR2M8mp/ZsciuGhqwG9XYGO+goImJytsb0BTDvVXYx3FhcQw12JsB+FVa55gox3ZIx
zAplZzze7wukCcn4oo6wi5/M4kZPwmE6JpinsEWWHel3P61IYFKHlwteBizsiLtmBkeHpEU2dXFu
zap4WY7Yb2i6zYb/y+tK0A6poLY5fMsbM95AvetEtSC5W05bKa05Sw456UcZzxTLz7Wpo9UeyrbU
Yt9JsLDZVTPRQPhe6EhDekv3ia3tU5tp9KCh66hH164jCCVRbdoalKVwN+yBIl3kiO3H6n84vFnn
/C0fFNESsbkD9uhfoq7PFe8zY8xJ16lo/+wvXmVwXFry4HOXM9yiZ3kz40v5Mqc6T1GCbYuC64vH
0O08+UvYJF73NZ3eE+3H28byaCZmub9StYQd5ZchjS9sTBqJdm+PX1NeT2qPIeClDLi4zItB9K+u
HaJSaDjrV+ZvLmWb5NeiCEJQzVWnawb7SbwE/aJ+7Z36QgYVmqLxupeYyBF0ueguIVr3NPydXHz3
2BKHaiSJMcnvEYcgLXh1x3QLUJLf32uMI44wBMk56HqMwFqcyZOGH7G3MFEA8VQS240zstxcmQQp
szUu1Jf8csOxMS99Rp08/9Y1FxO7e/LL5sKTjQvbIKzDBzxzhqSDEBtXCHb6mBwyjla87RT59EDz
p437KnMXZDB6K+FNesi8rfbnQ7NaMcOd3EzwOUWHKNqr1iHQyg/Ot4EB1VkEfBMi64VNQtuL7+NR
3v7V1nnwiDoOYIGPsdHgBK+YR0onj6PZJwExHWQK0TLbk8PfpAjqXadLnOPDkQKuBtz90dKFcOjt
6Da9N52Bv52/m1rJFwXrc8Re+kicjaHd/EgYVl86jBTabTbHhmCWfGppxLlID7qMoV5Rglu9ou/9
SsD7cXDvSxSK2pYths/v5M+K7iFu8fdnkzbHubF8GM2f3vOYBv4MpOIHyH5N2L2NBW3aVIwzG78t
84k/CZgJlaJ5yZYB2Z42f3oTz8R2A1uhE1FZgWXxNev5XGvk1pf9gWIk2TKbWC96NonEhxvSV3vx
5pB1jE4sWmsNkACWwh2UoxHoIMymLKRTiWkE/Gm5QPStTIw9ZzlU7aG70gIOHxMqRBh1MmUkkAtX
tbysMvUH9xPYIc8G8g4Y6/ScKXvpxikJnxUOnyvKo3wqy4nl7EIO7kb7jPhtiKxutqwTkzUV26pV
YfJGbCUcuXf9zVLux2HbivWQEZDBkuYB57S6tQ3RkbHASl7Ry45QqZMKeKTIbMIZMUvcy2HiNS+l
bo9jlo6yPbW9st7ldbERUSGBa1R2G611SRhUKhQlcqJ8Ips94g7/oDJ+iT/Oc28b7nb5aVdB26ek
USF+H9N9cH0ypIwDnqT0zdyw9RvrqoY+wbKu/P6YM5nokqPT68ZKDfgjCZWHiTQPYcGuFQW4mXfE
7aCu67NmfesCy/N31Xcu2pJDh+F1vb7Cz3QAqwcRbQxqIc35J2xsm2zujWaJWEjEmhtDGIuFTiVK
ns6LarZ7x1BZnUS0kRlGSZq2HjE0MZYo1VFbxtY9L3TzK2HsRCY/6yDlH9+1tJ1aAiUwEQ0paSQk
J4QobrhEKRgQGfTAOFy7WmAxQoNl2TmU862ZEayTXDHG5fLmHZhIlAduQyeU1G8m6kct4owchEJi
p4O7+W6LZfKZvgmk121J6IP1qAcXvyTVEPzJUq8228wSjHZWdJzzdVPAahzEQaX6wvjXeAOxtbxW
AMaz0m1TlfrxVtNnkNvS0xUBi+Pv7gm5dSSzZalbxie3wNJ6hCMwhIDuWiK+wFvOe+0Rji95i+vt
PTljC6+gYpfzNCC1/lRIDgBUq3dz4724adU4Y5eiC86BUcdneQQafeY3oUajMzMe86Fb1Eb3XvCU
0qBfT+Zx8Ol8N2WoXUYQu0A/udDk32vAJezsQzCbNVLDTvnThZka68zLZvmMvRlWpwohwN+ZZsWt
LhwJI8GjS+kZHez6OqKWSTENirk/UI8oX5kLNwjUmBCnJx/PPc+Hvn7lTv+TpzFNRZI7UzlKcY46
i/1D4dkAQ7d5NutAn6TP26Sp6vUvGD0k0aMbWF/4FAqIfGJwJPIt7qZuTgtHkAx+TpTipXkF2W1U
zSQq4YIUT9dQbqP6c1XkCwnye9jzHIpPUDJRnCuTSRtju7avbZzWw1i3PooBqgPkvFjLmdE0m6FP
8QW7PHX9X5j08ieoOz/N+k+89ZScHpr6endgKBfP8iK6vXGa0A+ki+lAqqN5lmdl0hmbq+5eM70E
YpqbcfnxiZNLEjgEVmegRLksFoyqHPz8sXgX5IM/RWKUj6r9cUjSyRWVAx++WYB5e/NNru5qQlI5
HS39L7plMQRaWlej+bTba5rGRnDQnx10AuwW/llXnDS0XfMXi+TWE6IK7LAEbTJHXy3BttDoe61p
qjJxrmhP1LMSkurKKpeLwKCzklY/blTXLdB+GU8Zc1gTsqzxnEk7oUOOBv9JepwkDUKIhLW5BhRD
BnaLmMUCClDhzhRXuE4IESwbS1mSgMIoyqH7b5hmCzF8/q/yMMINQj0hfjmz53lHUu55oyMWWKLC
p7hF36Az6Cr3ei7IEaiW5kvgRiE0aa98/c4DfPLbx4VHXKk3gfB5RA1c0YqI+jXapq/2AI8cuft+
Ckfqr0rBEZi7n8W8biQY9na+wCzShw9+VUnFXoAtSt3vh0FWbrT7uoAeirgGHAme30D5FISz17Pl
EFvsQHgAMEXZuHaS99rZF2cZN5FXDRJ/EMIwyMr827/22TYrmnmF/IrdQLcP1sT+hj5uJnvHgLOb
68a96fogkbOwb/o0IlZQ6f0CB+dI06l4J/ATUdoZxqVjvDFBbPCcR3CAsntt9G4oKttp3aSXigqU
2fV5Gv7CQ5DqAVF2t0hYQgWDDqBZ6rmx+noNEeo0npbPRbS8iSrSgiS4pSBlNheIgamyeREfpri3
w2E1cXXWVKccGeCet53I8ldv7PCu+CEtxfpwGdOHe4GlT9s9tQshg+Dw6S80SkP3EADv9kiWIX6q
bblwCQRba/2j3Uo+OJVt0jsWQ1FK9kCQMf0reRyWKVo48tNoy5C+APwEf0SpA0om56xQuQcLWmdu
dH+w45w4vhnz7tC0DnAQ4M4Cl0DwByGWzFffNA8PN8KJUJPKHfCtpzUyulMZcAAFUopHjXtmRRgH
TNmflqjWFT+5uukusFPzAY1SMZus2H60tpuo40yoROzB6vC/YI3gh05yqCHOuGEr7FeHVzUP1n0b
N6Nuv5pVyOB4RURBEZNpL8cZwuLqgPrS1XwMBh8t+ZuAWPaqybrvnVLDD+OlGkRLNZH1P0tLfnjq
JKBwLHtHTtX2FVySuRew9KVdFx8bN3YPisMgihY0bLcjANNnHJXY83bsDaPW7GhY08wsaShyVmxP
r42Zcc0yPDxf8m2YoWllE/R2xmlXECdLbBLabUlnO+f7vwbZi3veWpTgivYGttWwBJMu8ZdZ7iUX
jUyYBqXdj54q6oDJ+q9fM3arMrgY2xhsuTPVaZHPllD24huwDXk1dkfn3S8HXBsc7G7oI9/lBOs0
8YMtjlu/oQImDSItAf4eHjx/2uxqg9kzJ80MfhGLpF7QLaDNJTdmtAEw0kkHg48tTblVK0Ph/rtN
VzC4J3ibPpoEhvTUCQRjj2K3CnhAqB8MvfGRRKh1UYxoUQCkdXtboQaxhSiCWl+EjZ6bSCVWRfQs
lrz6LLlkLRnjiMSFm6B3g/nehqtbHxlNTF6tk6mybr42CrjmkxOPO/1SH9vKPvXE3480inURwtw/
EMG5TFSOBY+RTeeaC+rvCX6NZntM3qarMRDQkOS9rV0JHoe+3D+pclu/MWX69cs2pwYu+ysKjt3m
+d2VyM8lKJHwQeE1r6m6/FIru3tAfKd+H5+SQOegqVKO5Hgm+iOTaE139BX+5HTGB2Zp2rfA+IJI
+61d88ZcjVeAAsVWyXrSoc+0fLMtE1YT9WiYbNAWJzc2vcNu4gmu9AGpEyZrvxcQQKaV1BBifxTd
s5oORM7sF3peG+Tn7m4uHhz6X/PYV87j9bef1J59/PrePF7WrO/e9P1WVAHxtaaQXvyj3ev1/vKB
u1KYIqXMx/Wzd2ehwYyco7owmNsOXejyw6TDViIxMlk+pFNOXL3MphlRcq1SDOWaIR8jX8VsIdzh
PkgFnmJIi1dfwa3E7lCRSkWzAE2kyhtvLrItUR0YrcdMewOUOTUxquLsPl/vjp5H8DqUVQH1L0ki
DAIPAu4+iHOrowbDGuLRwTaTh0mCjjypANY7OJiLJ7laLq+nrK0tJ8xeuASS8UXoRRCMxi/EZEke
i64h92l92IUtBISMbCRf/2+cHbwwUSTdYdhjuzr65vtbBHmsNW2qRFI3XYwwcvuacYNQkUdsd83W
JmhAVLw2/B8PvkU+no1kHgYrp/rgPHADraSdcqrEn5LcHIiyR1x3HFM+NANBwrmUyjZZlbbRQMuF
dqZ8gbFI1krNBqvd1sQ64YvT1nKYLj9Ou52TVn2ffDITPyikv5KO+TuBtFwrNzCQjnwl9R/gZAn9
R0T70o0wTs5V0kJEQ6Fs+gfQ3dVXq+cN0wfoJ6QjyIw0nHCYW7YEVo0ekE9BYP5QXyaX2NP5VXog
/zhrZMLxVvPZ5ZxCVjsXxLNHA53R3xEE/OwPAXUrDZDavKEj33MBoM5pJm9iMS/Tvw9w6IyrwAm9
nHKFsNVQ+jteM5Yx3JVxt2VV4PBJI+a4f+9aF1V4OIqJgIeexTwtlQjqMfGHSABB+Nlv5kieT9Kt
hrP9Ay7DTXIcxX211UAgIocpb7boAMKBultbtNPGviG80F6qIWxi+CQa8BByKxYyyH5mNhO1mVpy
TXyV+e759wJgh+iDfTxW0mQPJSHXER1RZgbsJxEAjByF00tBRxJV+IyCtax12GIL9fjJ1HyP1d8Z
wrvjeUiqeFA8xMU6vMthOe+KKzUqKx2TVyGUcUUsICjPVfD3qCJw9FHeaUQYMqdGB1dvR1LuCXlU
k9oFH/e3FS/hgyTEGRf1c/Nw5b/ejBUaJ58a4ZbjKQ8Gp++2n0vMLkLvF02FOZwLipRd2UtFOrvS
67mFoeesO/dZVeJo5AfUpkw+oHcaUagp0FBVTFW0o4NmAP6Hm/HC/c+I9s5ez2TfcaXAMG0PRfPl
0l6xTd5nvhFIkjLYtu7ptt5G+jImXg19yEI0b6/adiFqocFCXsa7cxZ/4LuIQD1Bb4ZdhmwCCs+3
1dSZVawdMf0F8QvG7/nHmy5S+mgK+epnAXguSDwjEqixTQWKTD8902gblbAdz63qLojlfZei08UK
jTcA8+GgdIwspaMankALcdgTCUdXlWA3nmExekZyXqY2XeIXKss7w9X7MAJr46gW2JQF3hZ80n4A
jCPSQxDo4QKSkYwQHfdppNeJkNqRxnFiMoH7teXN+iu/jA3rVbGyPwA3Tc8+lHO7uXWqCa3FdEGQ
0EH17Bq2GidYtDm6vHYCZz2F/1qHHDWv/Eip1IK8I7kItc/cIaz8azTb0w2zi8Xx9+TRBN/uBqmP
LmeQXyxtFyE367HQ1cadmlOjy7EjOhUKyVBGaBODRC0STUJs2XDj0lqjDo6rH7YTAxGMqypYK/nl
u6TDXKToeqjMA5NZB+005q/hU6iHJGRwM/OscsI8QUAD0BJajFUtpZF9eH5vpQsIoZK8ca5HCEOj
7fSSHXhTHMShtUZeV1MsfctENATcpeE7Y0FDIw76mq2pGMdf4+sa2qL8pWi6eTA54QzXdyvwMjUu
F6Av87/TuPQsem8nHiIzwIar56+b1dDIGTQNgMkO2qHIyEsGTOdhLVOkS8Ae1v2sxeTrbppqDSdh
/IBO/4KXz+TIzOFZOyslC8QSvZF12WAaiVd27L6U6zr/D5lS+XPlHK0vAi/wKL1jFXQamaZ+2V3b
rwTooUTp+h+pxRKRFk2wkXjUz/Wh0I3d10XYMdYJkshomAD2CJMdgcjwtba0rBMkTtEidJWUdtrk
g0Q0bdt3UL6wye0vmhyzRR/ctRfc/BDTIqCOc81f0bsj6PM78GTBZCDbN5F37tg476vv1wFfFsom
aCtLJk5TmsK9R9cEblOfTVDT6Kf+jZ9I5oU+LcMVbAS00QeYaLWxIjRzkmnkA7j7tdSBuEorBqWi
XZ3T31hjPjl4l8CmHVTpOL1D1dTuQmI9CtK3CJDxYBdbDRZtK53xf47eEECyxQPPa4fBSpSkwCiH
lCgS5ESycczdsVkfgHNwV+baDgBMg1ahnIH/2M3w7yodWVmDD1xwdOrYYIm4dBovbTKVGWq7uPHU
YEy5T4ZeM9kWRceH5Ucdw/ZMF2Tzy4veMdJtNYvfcVfD6NQeOX36k0dOFRqFT3/tO9VZQhKuRhze
y7OprFmo6SZVryX2fHPHCjcdccGGzf13qmZAzFx/8+smy3rW/wE+p07vexTcl1cSevlBqDdK/qh+
h0N4Esw6QaaFURAWRQJN3pPFVPTrstrxho4+wL44knFZLj+lt6+nT3bLBqa2viQzVlT5b1OKflf+
1HbxQTngjiXtBhpR6XqxEeuY4/RJNnJ5v3A0/r6iS+tXAnTj7nqlvBsZ3A4CUKa3i+DyRDUGoB72
gvN9dvRVFH9wOPEJu/3zRQIG0J6zXN6kxw6jcbSUM/xljGQEf7u4aB3/E7mzbaESw79nMfQFCzOO
yC/92RsD5IPdicxS22DkAiN2rLSpw7+VwXJREKm5okqtEs1YpWjx9WBQrJtQvGJyCYJvlYSwn76z
JjM60/q55/WR2KtSc/scY2PEkhblG/qB+kZhRKJtW+omSo5e52aJeKStk3M17JDj29oERbfOUBUv
IQB3bx23rQejKknuP01nrgDqK4PJTYLFJG2Tk0uEg0NuZw8ryTzPtb5P2UOQgIaVSe0Jo7z4zY0m
npk5OfI0b5sIf+N3AY9oTZGD7EH0Uc3VqUt3qi5uz5gT8uFJi2oOYuSTbFSsyMH6clFgyQQZmvii
8vPu1gpgNB6mrqytY/SaIAA4WnwquAd4b+X415xLm7qfI14IlcwlB4JqP0a8FiVRq1YFz+WjInZB
XCbtgTu7qOMVjuEHu5b5sU/3Aw0ixYGJxly4uszEozBCKzTahlWwdOC5gizh85hvcQmaJvEQvXCx
bhc+w7wdtVHGWBUHnkZ3ZD8lJXz6Jn1Jrvt6BPGerD8T8fDmwHkBrDeQYJr+UpRVaRZct19L0U0j
5t5qfDqdveDCMfLQLZ/Hn4noG2cuq5wyv0VGYGvmaD6bAg711wiwL6d2BWGUMLO+m59sEM/lZcqj
s/EA5nviPdAV8oQSpMHh4wWRHc5oSGdcY17lJ1N+OpO9fCgWkxKGoWBvV4KCEumlgAvIvbSLGX2S
QwPQE1CLO8y4vInzQZSyUW6wZdR7p2TCsRF8n4Xx9Lxsj/YVBa3pVD/0j7PR6CRzymHr/lD8WRVd
VUoeoe2XkxLCcSKmrPsVQi+Nn72kyjJrGohh+R9rnzCFKnB/02bvkKtJLiRyF0UKvfXPgTLmpEF6
R0wvgaDTXXDRRUAUDd/i1PcLkVNf8CNc54JvHVpmBj5vd27W0YwnyeMqZITWKPoum1Flhz5T4CqW
zeqGKx+U2KEhdQrUDOmoZYL27XNL5syvdimTqmdQDnVkU6D3Uxz/ObaTfjmvGOGHPPXGO84aD6wD
Izf6rmjJDM/YLPt4dyeckm23Y1H4VweaBCdB8gIbulrEgGKmjnYFYl2J1opLgDkGHMf8b5HhGFtm
qL1DHhzdINXbSIbX5KqL7dSHx8OBxIOXaXsEh8DBn4PF0qZJvx0KBy2zIYnhJeBEkefn66Uv4XtU
G2q4vQovXLdAWwSC40hoThdQy/VW7peMVnLq1fPj1B2StVAAyuLPUrvoLj8bv7TAS1WHUEj7xklY
oMCP4SSKDQVhoZp02IahEN2fU0ix0ryzygFHxtDWpfq2ScyyYkXcsiJjln9htMKX82H16bKwSE4I
3QIFtbUoo5+02CVRmWwxcntwoU+dWNrsXv/ZuWKkC+DOfV49BF1fFY9hsusERq6TiDgeuy/S0TxN
u/Gubz+rmnj6+LW4PkgNOSPSTOD+nKUrctvOVA27lHwf/CsbHzjUzkJDBYtXDSRM0RfoqKGbZNEP
ejLhkHn1+R7T9S1ckscvQOOLzOmKNJDTBP2WAwGL5JK9OMWmiRmPP6Lyap2kUABTbmKA6C0YR+yu
MmNTm6vys6wF5hbTRKfUjp1RkPFYjecNWhvcPIDep4y/yWBWRXBlPPynV2L60NagcYtfhjxuGod6
m3YYq0JagxO4psIiT7XUQPM8RLTLpRIMM7bDKrYSA/fmdhBzj3xFJqv5qFjRx9kfveIAPaRfuu5c
d3EQlevmhLpVqH2Q3V24g8TsPV4wHaVhps3NIDbqNKhCOxT7CuQoRl92ymiT58QVcItIXkgCXkb3
kEcrr1/wCvf0JW0upOlTcNmp0O3eU+wlbreh94SWWbYKBCMji4Ep4tRH08xrVLdHvdMvSlTXHgVc
UbHo72USlfoco0VM7/y/L3/uB0LRX5gj9bH/s9JiufxXIOOE3nrJ/s+mIuShdFpOPTeNWFxj0DXO
o/PiQoNtrWvX2Iw1PJtTC5NoWZQlfP2OLUWWeTvZaiio9P/HI/jkE2mGzBEn+t+VvdSp8whfPMfs
dvNdCXffQQ2NtKxvggIz8rEjNqL1l4wGauSdW7sEp4G1tK1sWkxJJiQIW1UgWs5nAtxZ280ycVdy
nH2wPlzK6EmOCrwvhcvQTaHp5JOP7k0Dx/nqgH6FSMbB6Ae3FLvfU2sLYc00XgGlhnVxHjnyM3Cv
OVp91qGtbAxuN0bpj/uAk+LC6M1yAm66I3PZ6wpq02F8xofifvUXB50A1528pmAU4E0zPLdTqLZh
LNJA2qVjT5oX6sE363SV1hoaLgNo6oPOPpq6udH1RQgBEk6WyAHPlEF+UBvCcb35mNp0Ocpn0M7w
BX0CUEW1ktzQ9tzRvXC1c+ir8bQvTnJ6LGiJ53jBiNPovI+UGyqsnR15TXg2YtVZ422a8VSMUZJ/
KH//S62LBsZ2f28bq84xigxgkFSl5vpoZHQo1qWs+PrKHwsDDox3AqjvmV4A6gCtOcmQ1tggye3X
QaweBv0JlfpmLz1x6md3m9yIP6pIeR/rLGYCYqS0DQt96K+/KTZDPUeyEa4fesvXWLiDNEfAZTbA
H8SXkE/739GDHk01VoISeCWCoH7L7+i6nMcjuoMd9pbyBEF2PRw6oWvm60gHU1Cx77V5RwPeGTgO
t7ATjp9dqOJOxZkYSFVIHCl33y3o8vfjevAQJ++ZCdE1r3JlB1viZi7eXS2QzLm5QdJU33c9JE8q
LafyzI4a+2tIix4XHLNjlklLDOlcjPo7yQGPRVicQurO+85vCMtrXy33LVsZCEyr4vOyxFv5V/IA
mrE8M+rqk62ySXYvMlIDqpUUlLemC2rmh/sPPU8PauQKtKNmUCm3ptkwiFbuQxTpOrB259NAUppC
w2CSBSFoyRYYB7dnzn7aZZ6zgrWU+CCD09RNgPjcLTGv3D89tE/s7zmJ0ZX39V3h2yS9ZIcSVe61
IXDOwNGRsyP3++4CMiexcnHcWxxct3FzF9ioLHm1NFxTREwHjpZEZpCQDcmOC1uyBgBKe4LU/dsx
yIkzwdzV2n/CHU3Lu4jyObnzfHyDwber7wIYT1opgDgKFjQOzKRa5bZjSuxwLBc55I/hi5Pim7PB
TKocmw++HAW5JJw3tV2cMNCgxsJSS8Ut/MnbJ1EUovKUGhD/0J0rReHELZsPe2F766Mm3R2wDxzD
io3znspWi9a1hSW4G3TYS/RfSmH614/VY2oRydS2nVd3YxQZjmH14CT9uEV6X0JP3HrP6GHR6qku
I6aoJIOEjzwS9jkrE8zDCRsCkaKdJodyiBIzhH3WUmPDUT7Uo4YSzcl7ao2qN1ERatMKDQOQBW6o
AEl45gPAHunRnEjsTS9WPfDiEDgYtOcxhsn21TpJAGrW5JGD0cwrP4G0wWazja8PHtAakA90ponD
yEUmMcTOR/QB9njtPXf5ID8qjVQeBq5fEJruM/JT5JpLa5zG6k4o2+wM41P/GtPDlAhqFxA8EquK
ZAopyap9qdEaT2a/3vpT3R50yBsD3u6FUBzsoCnBE20C1ST6kFZ8LYk+rO7dZcE/HEwY2A5j2qXC
N5o4bE+29dTiGU237/j/Hvy0H9/288OiNvYpmI2vvUFeuAVRHBnPVOfxcHZZP8BF1a+mjN1o45RS
qK71rybtKyI/qsoqD5RITMQ5W75wlJSDq7gzro4MLEPWpXQNTLD0zBzPtCz21MgnOs5y2T1ESwla
UbiNEBCO559OAfIbDOvTpsh8uRu0WmfbAJlJxtZscc76gpcUVmMrm4AgO8jiOhasdkSVhG/8oY9A
ofQtal9akjMT8liXWWRN04t0JN/u3076kimVTtbVdq+mM6RLiZCF7kzTDw8ZUEX1P5WfduPWXq0w
SP3N2N1lgaFSoFLLwK9CWcOjNWBIc2L1aERaWYowh0AkwempyVcubLy40CBsA/tfjjqp8uR6QDAt
4WavIrM7p3LyTt8sDa7UbexjIvqWKZLhMjKYqgkGas1zTleGFLGbjcrEqDdhd7mmO8wcp1aAlSkA
vJ9gMHaH4LWphKcIVzfXTfspkO4zG1eozG4HIsQrbkYafEpN0dYtar9OPriByxkCiHg29O5ZIpw/
fcghgV8wZtHvldTkQi28/xkegtWBS8EvXbUfrrM29Yv8QyEcSjdXQS6BIZciE9NZyZs/zIHyp7b6
/yn9Z8L8swvVYO/3weS4fZ1LzBSCkJ8puBTKoMZXoh/3H7fH/24FQZeNgRUZzqw7aEgrLFBI1nCG
v7viDYe2Ivhe6PsIMSEG2BDCnUdKrLVdaStjPAxwm5CQKHnFwPd4DHd3yd8kmqvdNx+F8xvqafgC
qDy3Mg3NsQazJ/+YHDNLv0FudCONEgLGd1WvS6grd076mtJWlo37vQ2SkLhF9gLFAaeM5WSpHcb0
nTI21vU5wlV9qiei/HL+c0NqAi+Bw2g6z9G+hNBHWxzQgXs34+5KP5x3H/Rj1OPxBv9FONrbR7WA
bz8D81tIhdGLd1g7Vq+EtETnSmN+idtNZ2N1QmGo3lbdyfJWsJLgWf9VQ2/PPOACHijDDnY1+LAl
UHUF9GT5ZzHKPPRVfiheUrNA+LgImg7R/ab3kSdeDqr59NUE83H9I7XiEFs9WWUEe5xlBFG7eCew
epf4CUm3oebR+r+QeB3Eeo7Tlt4Q28Mgfu1GN/w8IFHE7P29Ko71a2gRcIclXz7sRnNQ1u5Yyjf2
/xGNsidIg08+dmQBzR8TR7sPdB/ME+6zmc2aKuCmvTk4sQbn7xU6ZqUaQt4NZ7zcAYx3jr53JnAr
nOefCVW474SZnDJlhL9szcQb0y4GstZRNMlB9quPCH6xLFFjDEvE7XDAwsWTU5Ukww9BW6hb5TYL
E+vGLg0iMIrHz+9Ea0T7HEDZ/VU8na2wie15xf1SFLGXP1Wj6VEUXSZQygnYkddxdNAlYDfiNzv1
7+FA6voi9pfY/6QkOhBZITMHlRBuowArHjp/npz5555OuJKU5r9SNVncbMu/u5MZfBDWwQkQUXkt
e+6gFTBuNNHMZctjezUNOSyF24QftuHa+3OTT1DVwl9f0vD+0vU7ytcHLOgcCi2AeMblZLy6A9zq
dOWP5gUtk7zJd6indNdAjBbY/DkZvbKVXXdW+aFF7oAwjmkiEVXYhy5laBFBPjDynSPDuis+ska1
im+M2e+I+MdO9JvEwGUbPBSDL72RLdYHu0J/AlRRAQyA21YJQudQThvZBDO/QgcgdyanoJBAbFyv
0sTivfv8jXJMyfhRwzprNgBvFJRnrO+A+p9WqcQvG8mKIxOAx728bMC5olGBe5FzyMSdMDNHGYpq
DnryH6TB7uS+9sRqrCBpr+pKy6EAVjmYZYAJtpseRtDz79e+HNU4IvMF8vSFFsA/IkxNWN80o5Qm
ZvG0efCsPZQMmcZRpsasixNJLmh4/3dLKX6HW9PgTgAqQbzSS3wi+wm+/tqfXnjWsoy9MXfpPzKD
tEiQpZb1IXbZn3lW65DdJKBj5zDZM8+WcHwUKvEUyfRyPKw9KvN5g/jqt0vlG5/sgHMAJrUt+ugu
B8uisFdMYG8RhN/SpRjzHrIkFvWF6E+oRpdF422nrjz0q5d9wzu9lJKlkRCccMdB7NTYM4DN08me
dTpGTRJt2A1H5j6VVjYBZFL24MfPJuJ/+KelE0tpimrXkscixcP6vzIDkp68GQxO86ug7ksXqjHX
m5eywv6uIbbnuiX4gG95BVZI4kIv0te288G2vyaCP1hywGRx9psY9gX4zwcTcAM0HlizNbp6RdlZ
6/EebCLguZASPS1BOEhTyKPKrHJXglNFzGp2YwoT4iWJH5BymDCAhGCGINNL8SW9t7kT4xlqeugb
Ue10Xy1WpV/vaxum7GBOXF1xUDSrcsIRmwk3ZzTiQJU5UTZmKCoaorTAF3miDQPkb2LMCa7OHkpf
kBoZV6E9DBmBdTkvkZNVI3YZTfhTeTq9d5VVf3aQiPLY+/oraiThL9ubi220lnc/CbHkgxBban65
vR4lzk3OrtWKAK0cGKp35y6NmuWlj3DQs+/jvme/zj99nK1LzJaHQxKtHXy893xR4WrTlkEX76jI
D/6zlyOsepQ9wJ7Ozk/E5LbXmcFO6+Pq9zmObMZPWIdYmNH8mMrsaOhf9y7ECB0POW6ZXqfQauLE
o0LaePL3udTgrhrcpUS3zEaMU7nwQdlJMUWnMuPQS+paz2sulRzkdytt7MOsQacF78+U0Yy/piFj
QnejK8ELU1oNZ2qcxcybGkpA1DoaxvtbtNjrT/vR0t8aO6Ydk/Ih4UMhhiI2BWYwo8f1XsCZBv3Q
bObaz/VsRAmK9ECknXawTM11K72wN+6CHIxcW0HXeaZPqKZTOHccefrVz7h40DGUTlCSPkqANz6u
oKwcesKIlqQxVGsgW5gUEkfdZk79y4SX1dKnbyNeWmQG7UKdjP+Al/GNa7o7nIXVtkknwgYlaBjS
NBKYg2P9XvMrL+02gqrarn6/bCUT8ETIxKDGSj3HhT608JUV5glQzgRUMB2M92aCoBoUgeJ6FZfF
ig4L9IAQk731FgILn06Cko/y/yuuC4ZkDaF+uyQ/U2NGq3fa5ZQUQ52TzyZWOLnyDrwY4uCkE9iY
OLHKL8wh0bZMtf/DOIHcVSSxPvS0ohHQdDmmDNzOT4IgogC4PcMQb3/xmjs1TLeS/WI2uUk+p9/9
MEywW/5KwTIbEal7Q77GU6hEJkQztK8OszR/OounLzd7zI27RCjWzzdjj1uuWFd2PSMbISnQ7DVE
PbHU7MjBC3aq3jea4JkGqDX+Nd1j8vryMTMRO2bXu19HlFuSpbNLU/f4mFPwwX+nXXYZk2BhArub
Yos+ZzPJA/NBNedHmXKKOvrEeya/3pqGW0J0rrCMIBzA3Uo4syhCdShEXpXbi3auN/Ec34nFNxrh
M5XE/v1/Y/mVfh59hMtB3ajlXTKfsdksTDq3R59M5iLVC7VTlRqIrKAYIAqC3BBTv3zl4F/hjFuT
zs5qXCEy8SFFetpAwogVY0iXOjxV46Lwz6LIDJkLLo64WHKga8Yhxm1lWIhVgaKyfaRgBZ72FQul
95/YI8QbYLIrvhki7lZ596sYqQrHZdVbYzsBspkGLWe7H5VRx/Ku9U+1tFs2BxAuZOwCUoy7pmaA
jWjY34pLMHEN7ERj/qKKgY6KCzUV+5yDWoHp668kMn8uMTLcz4dte1tdtY8ZPjEBT0+zGAFrsWYn
OTgE5wz7BeNBqr7XdaKxdrQXtNXCz2jPxgLBn/N/kpwxGsfcDpEERasCnaUhGlcBgFiF5USw0xbT
4E/2OzQ8i8pm0v+oRA34XZ04FWUr0QqfKGrGLghDyW5T+ogQq0TW1jTbwzf8nhMDw/9c2+BaPFHG
ieY0j9oFbog5eonSSWaGKa8jm2/kvjvvlIAN32sIE22GKe6Y1i/weWMoUEAWrQmNZ0W+hyrDXUfc
Q+NFMG6nocNPLQHsz7eyWwQLtcX/IQjvhit68AQaUniCus0SaTY+9jKUuG6I2BjS/O3/74xJtcMn
dWAQT2pU+5jPoAm3MpOrNWgcncggFkbgomN0jLUv3idaETmWRQlNWiGNNWEjNuB5HVcAewfLOIrI
08cjwvOw9+vObzdkizPwC926Lc894NWqcHZR1gCGOOPP3ka7JROwh7+IVs1GKmvlWHJ4ibxCW3K2
dWDG685KVpVX8hGk0QZU0JaPsOnTBs9RlJKsK2RdaAQBD8A6zWZxBLMkYwBBv+8MRE6qVGyElYAg
BngoGF+NjAwm2bVv29gUFVhexjavi64Lku4H+lmsvDeemF5+nWLw95JwV+xM6EpnNo6f6q46epPy
T4oVq9PIqhge/VoRmJR5wdW/M6r+kRWNETN82vTSRWoVXjOc45+VUPDPWNzASoiqrlXbDnc7g8Ud
alm+KFoY/OM1W2W4VowV3UVizr4PVCUC2qX1fbZXIHCuBEp8rLZc2zFOz9Us3jXR7L4oJt/C728V
ftQfND0mj0lQlgsleftF/CMbFQiCLyXV3itf1B15S0eI28DFBGm2hArhwWrDQihFNq9OKYtLJRG1
VJenuieoRDZev6yNKANRjz7Ubaa4Kjsqs17xcVSGNPRXgU30lKH52lU0tlEBrTx816/M7Cz1VY1x
o/ZTTtszf5DxW7yuJnJo6i8+GIiPz1Y0Mt20N4YU7Bll/2/kphExTUIzGRjaoVHYpdqRG2laC+q6
IELr7Io2cpgPi0+v4eFp1h1ReHyVXvBWJYCan8ZvlLfZsvCGbBbJmdXZ8z6Lbhq3nRiEJaldSMaO
7QAafdMxpATu2ktLZ/TT+LhywsKYs+7MeUNFMtuDPk7AhxFGSNLU5bpQNCdgLtLRABtdWaZ3H9QK
C7qgvgWr3Vrk/xAChZZ0d0SERm5WhxnoEuF+7cgkR/34/xJftXka1KPuVHk1Z0QxTKtf8YQqao41
rTTeUsmJoUY4Qo5hME38MrKDoCZHBpowP2jNbhBQWECIHqhsjee2SC7mTlPNMCIVQzQIffnqCo1t
fB9D2FeQlsiJRL/FK8Is2m4Z4ogqWHP0fe3VJAp6k7HpkFd3e+sPLMfRlCI164jVWzuHlTGUDW3s
I5x0N3iVZ9WM7CPJnOUIIpwRzIGfQAKPdBADcE4MNj1lbCnwnXhkJ9LNUMdlAUMpP2rUX3WZJWF0
/J0KBOXCwT+bHVKyEwkfn4d45YEnR8Ke/8he0B+KWqTk3KLpTVcATh+e4hJDr0GtwziRFZ3hmPQ4
7YnTptsjs4JvIt8Eclwv+6NHo0E0fJBUFBL12BcK5f/fBomtXqjHFP9BWn+/gnQSo6UACpmJb5x0
Lk+APz1beidLZrGpv1gIj2HyEBdEv9w8eo+oaV5QKcH+8ykRjIUKKc/zaZWDiz6pRDz6KEt6taKl
OTuA2/AAgzliJMC8pxpq2L1P6lgJcyiXhi1RdDuVygS9tiwFLsx2bfhm8bKgDoieqdScYb7uzjin
m1EiBUxMDQ92TgB4D2wyjJj9BxCut1jjacRa4kW7eo3ZEfncGcctCCxHJWHailfFMaEclI76UEAP
8SfGHDzAlZVwhKO5KBZG9axRSMBTmkhr+UbQdUJtDeeuJUH+eR2SEM2m8yBFKeDfuxHsBRsVqq1D
12lQxYV4Fg27Sm4yNpDEfRD3vnfwPdUFCCqWp2SUdNeQ12EJAuyZMKUreXm0yonYAp4re/Eyx6Vl
Ahm8YpKHzqNCYKFO8na96CJWsfYNI8tAKR3WLjfYBHS5V+452WP9GL6g5nJExKkkSkB8Hn2XbyRE
dOivaEV/zyaVrgt/203TQdG/Uvjn6AjgGn2Nh9WPAcoefu+EO8zwiDoowWKJNtK1ETDlqEJcEJA9
KmSCMZG4aRX71zxiRtKamvektYiD2Cn2VB1bu61XBuobIv/E8ebpfaBK8R0CaJlOPPScHKWWB5cK
v5iKDzqXHbbF7STcidNLJomO8uv+qxEaYiCTXRxvEDr+99jIIPXhSpdykD006/L7KvFY6dMXxxVK
VNnnbplH2irT8LI2P66bID/7H3gNKdFOuGxEMdJeJzN7lncPQ29DZdptyQhAnqw5RTnNDm1mdnLC
ytcGjK1iB/VdKvjTRi251B1UCgYdhX8DsgvoPDUlkjemqQPRR4AvFQnlzti7qQtQzSGR1MLxjxan
Bhd7tj0l2PFWK98AbICruKEt9gL2AJiKyMmoMHdoXLN9/mk9oo1YGMpRz3Evd/fVHtgkgnQXkzkx
Bhm+ZC9YTxEmqqPSxTjRGBX3EXQ2A0ocn8B3Te+JnZlO+w0X9lfjuTtZ0XsFalOD6nV+Ua6ugK+G
1VAW8XaxEGMre/Bc5bozejSiK2nax8BKE+MmHLJpwvjK8TEZTf+mFzFE5n95O07yaCGVrI+NeI5L
hUM1BA2wW2/SBAvdkvflnQqnHymEcyRN2wfnGPlYQ85FRCTk0H76YG/g9GUvzxVqrT7y4LQv8qRJ
VZhSW/mk2yTOVEb8geRttIv9LJ701Lc3zC8/0vpUxIW9PuWQddlSk5EDhlbvybhtqUE94kojjpQs
n66QRoXx+NgeL9G1RjqgJU4Y6LwI2o0QWjdekLp5rS0ycgz0Yv7vGLCIe1RuuWxTfVIByCS6jvRI
2XKspjMV2OcVWk4pkWyezmqTh44mlj6G72x6EfOGodM7uwrM5AYPZUjcnl0wisWcvFeB31FqFxbV
te51803Fyt7d0Jo0NsNwX9Itr9OfaR5kWopbif1UgB2g9gdFHDEVGhSl4PL+T4oBtO+M+81HMlcG
YCD+uJdM7MUy3PKsbUiKGx6YysenNB40PJJcs2Ogp48oDVD8SqnsQZq1TZGGOcF1qBZg7ejoOV9i
g6fQLFMObBUrghH1s9kziS4HNnG9eohySAeqI9v1kpO3Dkd2LrvWScZjZrF2iqRRwe/dOaJdveNb
2laVgF4qvESYteid82bG8YU+p2Ec/n+Aqv1GkiFcDo4xMy+ClS0N193vY9gEhieZe83iwY5LvRHG
GUB7Y/PIKw1wmv9uy1tw0+jMra6gz7L5sXSi7x16S7Gs8kphngrfpgXEN70teEQwACjYXWX57mwr
OR+x4KYHiYtwiuP3TjR3LFfwIB07mvVdWAWrx8XlwzlCWfuCoFnQrFdVxSzA8ebWWkU1wmA91mjN
rVF80xdanOANTDy+EDBzopMDTJneZWywLH6NKIFesO/uBbKB+c98N9HC2w6eGFA2spAqXoFdpKqY
ulR/1lfd8t+3QSFkceNg77akLwm9HpqRPJ3t3FO+ffYTftA5jeMfzy4Okl/Ud639ZIiF24oFEP2p
5BMhADreTNZC6OFg6B7qq/yxYiXh7oJvnYdoRPATFJg/JBVy1EgTt29OlMmIgtCwauAviue/A9HJ
rsaLgz6nSgi/G9vBBCM9DBqqV3XXgf2kvX9hO1DMlaASHcfu1OcktEFnmupxAXXbZUn3Xh+xrG/5
h2tD85Ry6BiiBKwXGQPDo+O76J3qd3fDpANkOdALQzG3jvanbqj80s5iPva89sXFesjhMWlcikj7
S552meKT91DewKBDnMM9ZcbNn8nccuOeHtYUiMsUVm0f8fTuJQP1e2LP3GpimbcLI3u0qpzKWo3i
xH0hjjyQx33JLfoNab3AyGHHgY3suVQi2FWo+XF4w6S0M1R2NTMyA9SCaWbMfVJThhM6V7dM70m6
+1hJvVuHwCl8nr1+tZmcj3Ivv187bKmNeR2I0hvbDanZnUHqKznDyZt+5p1TyCt3qap3gH8svSV6
v6/S3ged4CF0SdTcYwkLAZc128nsZIwyWzLlvcJokNXIithBAJ1Ctu435BAK2dWr3nNRJwNolEbq
+7iyszTiH+8cBh9YDxFRHwJg9MN65cJzBCKTOxziWWF8xZEHRFuOka9niKrwPRR84b3rSC8mnq67
7WZdNvNiDc53/U2OZymJ1buTGGPhwQrPkNyNrR69ekE2ED+/C0VUX/NZG9LNJitwky7D1uslsXr+
5QyY28M+AXz303pQSs84oCyjFvjpc2IBgeuOVL4C1KZ550MKZYoi/shtqK9MdUMnTt7ZjHx8+Z4j
Pc+d3J3akknd+5SA9Uxuh0ZcPg/97JqjXLXm+Z3edo7npHVBIIcWqv5nXn3g6xQ1hTfSkQEnm6sa
YSsJMzXS67ViX8bycW0Rv0K5GYQx5baSgRzGBIdVC0dhTRXNkHAvd0onzNUDtLl7KEKWhEdp4PDW
WUT/PMtz3DY4VZrDXJAn7Q3tk87M84h78QB4HtABj6c5g/f0taNWcW7zJ4hhPKD/8u54/uA/kAf7
QDF8RJjtw/b138Y2t3da3VWEXrb/RudE2GXrA7BDuLEBWm5+g995O+CFWcHDeJbc3ML8gWv06NK9
wtDkuJpL5wlVzPou4jkOZfeE0bO4Bpbc/8eMbTfaRBV3mGc2QXi5qxXDD+ZS6BS8gmROmsZCRHSV
s5IMkzdhuRMgIwb4OCgfNJCD5IWiFRlFhfck3KPlmE33RtoouEDNOPHHU01tx74XdWyyY7cCZNsl
SXr9YYLJtqlidGTaXH1Cf+2wwikcg5RQV601fWEtXCjDDDuXbRuzcoyUg/InaXpQv+l/S2gZB7Yj
i+RVn0TT7BgG7xbn57p8X/eLR8Gd3TpQs6JfjGGUKbdn0LQp6KgmfMf/BDnLbBJJQXsvR84RYBDU
TlFL3pbJ9uTUvOMTrt1tOOda5gQHfeyRO06AOloB3TWazAr83Fl/HPevKDOEo9yHXaPG6Wj9T+GD
WRMt+G+fOWBTb1UV/81EJEgxNLIm6UDSDVdCv8r6XU3y3aySkBx6E9+LD5J3g8FEwDncqs4DQFnk
ElCqmCWMGf0YItDJBI5Kh0K+AuU/PX9KfBoM9eL0gxhyUtdTKqZcJBySu8x+yhvE2ND86Oi7Ta7H
iqzB2kZV6vKn/RivkE/wyBMFz6/SMJYmvue3zD27wOZBAgR1qxGrPY9afodQHSI9Cd7W+hGp2iAR
GODSw7wPV+czx+o+r97rAirzeGaN/C3YTQk02tmhMXL4Owv4lHrjq4awyUELQoP7/Uh6Sr8PJJTU
RmRVrgQ5ty6PoIcXTB1MJkSh+mWSWMg7PPISViDCdwtCsKIp0CSUxGasb2yKFpyuR41O+egxUi5K
2l9YBWqXrdVolDdUxu6CN1wZpcN+fnEHlfEQriOA5RumfrgT6cH9VK3tqM/LJJj4lvDxKXQRC0lC
mzaOP+CPdYXOPtR0HNOkjq3FbK+eHxXp5iJf6KCeYnuezeZqRr4Dd8dD65P+ZZmQ5dPyfqpXKi9A
o69B72ysiDsykpCWT+i4nUMmj+Ic90lH3lk9WGyTvMq7ATFH84JF0nwo11TSzF4p0ix7ZaUj+WZ3
73Jov2ePjMJTtMyRI3gTyQgek6LfEDzZyrAYIvXmuN4gHDDTNML1ByenhRUTFW82j8StOaoAb7Sz
FBCRBjf8v+y7PMCTrQP6fhuWvNIl+l8UN8SwGEnv+zKFyzhs7m1yUv5WkXZbT9cK4DJNNLceiZSI
ws67rdVr7JJxOxiQrrjNMYL7bH8QRu4H/hjga3DEKfxPx5QzuNz+vbLJHSJMcwA1efZrjqLO9sj/
aG5cqKv/GeQK4N+fn8/3s9k+3w88mVpLew/+mAw4/saXjAj+5yYZoGsx0TM9deUfMz3zTVNQtf3q
Uko7c2eq5YhPjA53ek16W7GtHwVdAGxwQXMXHLSZznG4s0zszW+xSI4lBLJnj82Yj8h0hUvk1juX
sc5JYbybsRoiwYcZNAaQ/PqxIpWS3QiM6NO8OmvZ1MoI6N/TXQfr4EzEl2TyM8lQz0Ay95ktjSmf
MIAa+pQ4AGpzoADThG+pCNoASEvex5sx9zCG2xvXk3wkIG6GHc/k2UUupbww7YGRAhDUlk4oyW4z
/fBhSHFpU7tAyyu/jUYxn3I+HvPBTCvUYhJJQcydtt4QnBsH16twxl/Dgcnr8IgbJ2R2UeS9uE42
OJeYgfZiN/O8DOsu4S0HV8CP3RQ0Wa4T+o8m6oJcdPQDEN1hBMjTzCvdNxGoPZCVq38I5EGQsr58
vZtJK7xaQSeHBLX6ro97bsiEVF9d+jNvBpsYY0TrMp3kKB7W0Ca7wy3F8IPgF4+wNl62UzVWJa9H
EzghG7LD6iMWJPF5e5n4PTSmxQpnc8u/hRKIwNxgAwqNC1GGBubUgB+Xr1SZRPNztBhkvMXe2Xsy
kkpPpVI0n59b7KCO2PFoUexSNKeAkLtcxpfHo0379Ozro8Z3vP6PjIWyC9NK1Mu7GjyP6Aek+bHb
UncYnNBK/HJHf5oR6BEvUcprUPpe6ZU0WkoKZZnnR+9v4ufnxw08fcp4OXQY6r+fC75+IMbmrNPg
FRWhgwYAu43N8AUqBLhQ+2GSbacZUiHE3XWoR/BDrYQ29WfC5JEt2kNlbXRNRsuth5a8NIgSQe0y
9roKby84Js3FIW7xlu0FKCZPvnuIwF/qtuwJdD/ra/AC0aa5hzN50y4GTt5hd76sZTzadtpjW4B5
CS7S+Ze63KNDx7/fO64EWs1sTSWh/NYYsHzSLMx45fLmsq8phKM66hqU0JLW99r6xTdYuR7Xe94y
uCBnBy3U9whLB7NnINIJwXG6VLvgCRc95MZgf1T3dCSvdqcwy7Gm/wFWT6ZMMkRQ1rrWyW6zMFvK
fImj+nlBErb/Y4EP/u4owWqMGu23LNAI55cAnPFVyj3TnMBYZZB+uYkIJW15ezePRlL0JxGRkg43
zWufxHOV4VsPRc2yRvqc8XDjeaWVLSFfnsNVfTit0S9zPjGRyHasAOM54qT2zeUUhpM57OxSu0wo
UFpR9lg53lLGX6MAwztrmwavCjETk8mCP44AX9C+DN0HOwzAp6FiiYxIjkFYyfUE0fe/TRuM/BuW
tqJMXyt2grI1ZC3mUEVZ+1yRCiqgl2cJ1pD7+CuR6Rc+ylw5aEENyKITZk3h3ABD2cSXeW/oX5uF
VggcQPCvFtfX0f9Ln1cp58B7wnfKHzfPVEjdM0eiONee5vz8y3PWuIGeiQvQ2pEFA4LuwWLPJwX3
2jw4irivaa6E3HeqUlMZ1XEh5F2Srqs2y85tDbsekqGIYWeIAnGAnoMPqUAIklfZt/YjuRBbxI9Y
HkoKN0Gxyw06tAfk4hegEzSj/GZ6fkw+G1/Z5kmBeZOwEYao0Re/VBC91nKyKkoRRZ3d1DObndZA
nKiWAGSZiemndVcazjxmSlEWwk36DR0lYLkZY8nJf0os8FRpt+8YtdSVDive+MC2vcoG3UcPSzoR
j6fkGlSwTo6xWPyysUZL19F5g9d6Pmhx6dxYEHsSqCuO0sFQPs0qmdNnnLtiMyyiuMJJ/CY0nrde
7LNYX2L+QTNBOoxGYhczQj5oXiags9D0m+3Km+QTjkdUGXQfpz5l2TzGrt+GtA7pjJGmYFfh4pff
aZT1TFwq4RdrxnqzlpSZiNtE/9L4lg8u1iM1bGKZb/TVGExSx4obPAEkEPC2hj/2XB6btP/GXA5I
QUmUrIZiSaOkTpCn75z74qKEB/tjQYTgN9817xqpnwdqTEv7mmCMy87i8vThveID0RP8yDZeVdtS
nJwjzaASqItHDrmbxVL0aTyucNvzLBJnD9yHWIgcHXNk38j4OgFJuppBrfzLH0L5VHe7jmzQD4OU
IQ7TU9e0j/Ax7MgpsSsca21LhTcvY9dZ3DTzw1YMsNTdo/5fZlpRJdyEyLOAEUD6tYhmeR3bxQbV
kRe2UvaNP/t77xAayTGFpOELm7cyzTg4BC5oXQLtrYm+OHbnFhFzCqax7YppOWO4AZ3GKRtJbpGU
8MLAgJs1+DpDdjSVhJaNfGLFhzZAeanWK4arLKwwYOP/vtq7U9kIqklWZ2x4+1tt5TWgYebMlppE
pHtVCefQSoOIgO9s/ZMO77ur3Nq2l+S3gR1cF4tqDWshDdMQtZNH85ag0uciQRaWGNYXT/0QV3NW
aNnN2L6r1JY3vl7KYOgyjz0GPaI9ycR16D06ZBzMVTBUyGK9WyPvSW+ftCB5og5hq/lk2SItdvH7
c3apExrFSbaHq+wCF67tn/4tW22rr/3WA70+rwvlspSLAdinAu2uflZA3f5AUizi1RxH5B6cVVTU
RsOcerrh3NDirvo0lZ/3cB8iAXqAqqGXfo3lcWgV6M2nUxyIzKaJrbzo3+FHz9l40s6utVgjJ65r
kHDg/+xo3Kr2gOsXQL3s7Dth1seM8TEu8VxwtZKG7tzaKsezay/V49PX0Qt5LU+s3ya+BMbiEk8E
JwB/WUrVX60Hz4payX35j7cyHqy5lY2XFKNkhQWcPK1azUL0fbywUwkAIKJaANH369jGiZX3DG/B
SdAawdbvRC3+ZDvcG3YX+J8l73YBjfa7RJo1xt9dFp3krZQiLIlCMec+Hd/dfX0NsfhekOvyk0VV
S93mlng9lxuy7pWy7u6SR/vuHom8rodZIerbeWIwUKSsoXeVV+TDCn+6fLR+82BbKGPWdxl2A/zK
TY8sC45l7GiLqk7TDoMY3ynFTf10ghuBclVgNtZS8nK2aSOyEcZ1TxLvndzf6NLiuqKhkiq1wZbk
cvrgpIw6NT1SaLQwk8YfflFn0DIGSxo5f3ETyrELBS1Ih6YaNnMy5SDfXCbrLY/m959KpqL+opmJ
G8jJ6mpHGkTLCqLEgvwNRIkArDdU/1bVaTmIJsAe/eNcnwMH9azZTB7CY+tKQTLD0Fxl6L+fpNXG
0GLevD2OzG7lW04IpDFx+4782hhS3Z4HIAuTCkxFg1dzwQ6Tb5mMWdFg6mPWLiI2y2UhcNTyLe89
+s/Dx7KTs/Xs/s+KH2drBWANZ0ZN9V49JrK245ryUXefWEMS7niaR8Wev3leApbQWobqjkprYEgM
0BRj8hNIeqbRezv2M5qjH5gIqXNIXgI0Vj+enxofcPeEJ+Z5Y55cHykoWIs5UwK5ddbKvgZOJ2sk
Js5wKP1TmvWe0ejoGvYcflotR0UNhICB9OcoEPLK4byFw1qBi1LGzYai0bazKauA3TicpLTtYr9C
eegoq4sMQ4hl5XjVIrlom6q9VRM/P12MFnMKdgKfVw7u5ZIcgmNRYaKA+Ao6NQ4kpuJ1ZGJWPuhn
tR531oHTO9GRDuu9jpWgQAgR2YcaQITbLWEDWURQU5a+OL5C3G2DDwkhBAhwNW6Bp4s7gea4/HCJ
s/mAmgVcFTsslYS8fk0+4Jl7yAqSe5BQKe+nZZzaFUQSXK/Jt8vC2CgJbitCgxg38WQ1Dnt0wVTC
+xnoc6d2CL5Ih3OkRtguqyBYoFOLQsHPqb3SD3WK5kfxbhDKEEBU8IaUH/t/tQyGVbh81Pqosi5N
zkCal6wF9guRdJLFTD+K2oXhNc9SKZEzDKFvDRvse0RkIzGwDnCD2dbw4twNefUPWX9Qjd1nmdUy
c2wPXYibE4Pj/EP/UcJOgOtkPI2qdjJb7lQFesiv9PebPi3VjmHy9vq/nU4fSY5GuTWmJh2fWUhF
qAThXKg7NBizsyJQIm26KHVEAGMZQvdaXiP4v56duqHJBh4orFpAyuBabMvSJ4D4aH76z8ka1Q01
bpmdDWbf2w7Nd0U5t6XC4sbOhGyodIJQP2oOdDdg7gT7aDceCFE0aDY+w59pNF41T/5ig8KuLqPf
cQ//sYliosWaozawkbxLUreDav10dAtMoqfSNuWxML+egi9nW6U4r4vAUWy7Z7IaFnMo+JHMXmqV
JEGt41jb+j7QXA/l2ZSa8fLWE52CU2YPjLLV8bJVTw19jEo7HK/d7PrRKbSrQqJt3DUAbkfsC6Xu
UbyYK0eC5DnIgo0ybqtE5CM0hOoIGRPBelKzjRHo4FKM1709SHpZHJay+pJbuhHQRcnofTkvd65v
VKYdHqUVOt5TdtmYH9inPdV1aPA4CuEx4qXngGC/Jj1urxQm0YWUWmyD35fijAQM69kqnOrF14uf
vmXpl2gRA+VVKz0xkQGiOwq+ZTdGOeYJELJ/FvSvAwefdSAnrCQx24qgIJFeKaHMhnhBqD4+JPKv
b9a4Wf4LIiWuglxGc5fzE6d1sP4qhr+Obeb6Jbl3a94LYSdhgDiIpKof4cHsNbAnTCpVIDCBkyd7
BKT810fR8ClfxJ72yJbguGAYsxUEKuWR5IbARyQFq7rLBkZNkxld2Px+iEkgYqxFq8uro84VvjY9
jINKymp/hB1xPXyQrnRzvIbB+KUS4YVHmZWQaFExV2gzK5UkKrZR1rBwFBW61VvhIXanOgjzd9Y2
3BNmNL6X0FZa0iSqRlDlP/8q1h2NvGWd6G7mqx/YsoYekfrbhrIytZYp7ljoppNMfiRdbLIK2F/p
Hq58AWhINeftYIyacBmgXc5+g3TkVJqB/oPvrjGdBU52dMiIelycveCFIU3KVdequFxEqheDw/Qk
TkG/Cu6yhDZEXdbIQstaUXZb3Vxcj57j7mTouLpcgSyG3ht4ASwKRAClgmkxcYxHL4eX7XwgwH1+
HoWdJrBraB8e1DFSZ39MGklCMiM2ynEoyLcs4wCBtAdQ/zoMOkg+wjUwFdVkF8mRguDlq8jiBeqZ
9j1o4gFW7TUqUuzwvnZvlchcwXJb0jLC2u2x6WA5JGoKa3jNJL4PeSUN7WSSaAcQf5JiBjEOwaWR
iLw3zWwXw5Hwn9KeQF2j0ex9Iwiv5MdLRVCu7KsjwCY8Cv+O8nar0ptZ/lavdEcvGstYbVkOqtW7
gBeMWhp5IBT6IeCQV5+qrdvyna8du+VougE/wnyK+yHia5WDDukaX8fdJIwh2YmuV3WNZLKjiTDs
/rGsAQ7w+ipMGhdFt7+/5uqYgdysa+j4aPEBV4TcgnCqVONIUUeWJyF/fxSDq3yKKJgQtD1jQpXe
qLD5KjnX1BOx9WSWbxaIrAqElkU81PF75ru5RJ/76PaexZAb0EJ5osXAXk1spKEYY6Rs+72ORAtP
fD8FmHja4jB5sqkKjdldABDYxqnzwpz/061V27bQqV1jljhisJgudrlsEIgc1YjhsFwL518THpX3
i+SpgSRwKdaNQyh65C2OvhfpoKsmBr9K+9ooHU7vUyT4314wtu3FQDhT9t3eZMLauNJC94Cifj16
+4Ij1qh6DRuBbQHvR+Qw3/cxnjVfCgpi9PY+X7kyusb1pEnJ6yIehej87jATbXw1N1oDz8jfFZWZ
B5qNS1BZ0tsjp0Xx2RcXdJBII0cnG6ERlx2VjnCqErC9hlwRa/2YjhQ1zZ+H3yh9xy8fv6EzY767
0XpFbfuH4+fPdnIcO+gh7698OhTlUE+1KY51pLFrW4ZLf63aL6hKNg9ew6aMU/LxcvQmLdAiAKlU
SWO5JeXNDjpu1ooMZxLHfVIc1BhNZQI+DYRir0BCxVWDF+TaAs72SkS6wMZoTEBHwg7B8p/o21wc
Rw9l9hoLpQrqZ+4C0FYUwbubRq382DCzJqexhl8vPYj5EUnWcZqPCAqY6mpCq5uiUk0nGuFtMfqM
2lL5GqVydLN7Zclng1W+lXN4SEplgkWTM7M5E7XGAtF22BeJ1hQM9kNtm0ZqxR1z61A+9oQ8MmQQ
g1keCfkoPnUGiYTaG8gpQ4kqL/yUKF/KF3026UQ7geqf1Wd4tViYflf7mpF7D7ycdyJbsmBcWngf
zikBXyq8OnQ++HTSZJ/Cgl6JYnBHEXHiqOjKQU2E5UCgMogjpa/6utwf4VV0kJJwkvUIL7uL0mmv
hteWbQ1Lu6Wxs52rTf/Wg7JT7U8MdFc24a3AH+QPKlzMpJQ9VtlltCH5d7PwAw8I+pscE0f4z+US
nDZ89G+/ZQnusMYdnOmtKmovc+luu524DVvZkYwauSxpWSNC5c6supUCk3RSegHlGvIC6Jr/Ax4d
FXFx6klkL/eKjb5mKynIWr127nDL/wDv3invchdT+2A6RmJqC0HZcPIp7hX7PpJN1K+sSvaZKNDl
SHsOy/KEfwTLoMdXvC7clwRB+alWb0zQtGm82fNwZyqva/7To8WcQEUgDlTA0v/C40cg9MyEwo49
k+Lvg7tkzeJ7c8R9I4KM6nQOkONBujPQQocROxPZY5VpHDmisLlpDQVLMXQu0PlnMWzJjXZb7MjE
72AdRHX62Zopr7FZ0D8M9/3f94rOgscE3gpKyZjJ7pGAjCA5eR0mmb3mTktK+DxICBhB5g844S9L
r/76yeFBl4JiG+/fHgXisXMP4gqF/ijus9bnSzJF6ECs6PhxPiQfBggFy8zQRcfkBYocX7lzl4aF
1mydGK0thadKxO1u92jbobVPGVliURzm4JJwkfDmOwuM4P2Nw/UXxI1yRNeryzsQe+ddixkqUEZ7
cXeC9lJNPoZrA0l/+CjbjHYO2MYhu/fqicG4SMREl3OwkOLNYwgNTZTe0InuGb069JjZx6lrvkcT
EcmRmVGpojjQTl/wjROMEilBoiViNBpmrCsUGxKNXArBqv2u2ClYLRbzNFtkPxoNBHEp6q9VChU+
dcxxufcXGWfWhq5YpOMAZX7XlFWkwlNCnbq1MwIjQTSLMdMcrO6ToMKmwqrgD6JCAkEy4C8DU1aF
L0Daiq/3L1Fyw+TaXYSU2ZJ5aYaMWZKt/z6GqpdA/1v6Fx5+vmzSeFSWyF+oyZnOvpwf0GDadgQT
PslIQoTAuoMccp3F49j3OvUU2Ix/6bYNIbJvwsTfUdd5Hly/Ab0/7GwAmQyrgGYw53WUqpzP12iJ
QRD+r9sgE1ryaAZwGPZwxBPZjn8x2Q33jMKuYjpIQenMpWX2aga1UjIGday3C2FAr5eZNx2SZktZ
B1yLp9szU4pEM7D8lQEnio2WVK2gvKsrsMaIe4gtHNKh0bRm1GiMuQxvq1jVTOaS+26zWwJgVvJm
t1mucdQWtQR1BuIQPK+zF4SQzIxaASzm2CVXiRRqT0LBP1lyMzCVMSGKp81wevCSMhlQ47wKgpRy
2piyaYew/X7xtLI/jq0f7mKCj2DmgwSLntzNZYPhwvgjlirvsIjXv7WUGopZPMXKuVl/fPA26/no
znuqBOGV98PdVKGuLOxwH3hHDD+s3YiiKpZT3OFZe+VVLIj/Ii5MsChpEO/l1Q6e5i031ryK+xW1
NHa/a1EJsNRVU/FiXFMscskSFrLXUnfqvGSH9ukYl51rO6kCpAY5wB1QqLg805LeYdTtaKp8CDg9
fTYW2c6DW5SGWKCz1QxEEoZCkADTf1/haWjcoi078oPLy98IC+oRGvPGfLCApAB3uaQkU3XG5McO
X2zvnfak9HtRpiXH/qgzVuBab1gsCB9G77yjtHTHZwt/c80/P5nfChyB8wYT7ORYOLLmkcfcctXX
h7VWGd0Opfd2S2kPBWRBE6QRaJk8n7aBhcYUAJyAh5bb18YxZ9zVAbZlNH/Zj4f10KvsSFDXHkgY
bilQ10fk7Jdx3i6uD3iFxj2fRTss7QKQMR2w+Zf+Avm7M4qg/reLTatOAV8o6TAYba5rnuCrlVGT
iapLlgWyh8mV84tfz10ZdwjOszVjbsyMEAQC2qhrcFMtZ6ZGO63oXSmnTrDNj4zOFLPEQPkzPH0p
99Ji1C4rCvDPH065z7Hz/r73lvDz7yioDWFZT3JoigiP+qLxBg1tFWcc8Hf37fn14/SyG9QqPADd
FdpzR+aJqvxxYzn1iPhpjdfgBJWZ2yZsleiiCizTR9AJbayq/59u9I2UpIhSsijUS7BNvhjePgHw
wbfXRMg9vMCn56MZnLYilmfIu8UImMuswojJQbLixZyv2o/uschtlM7LJTtxhVdYXAy+qig/RVID
bmtxQ/sJrnvQ8vnkkSlSDvgB5opnd3GvDQK92JkqjyAgY8SBVQFJonMutRrRLgKRU0NZCBOGzgng
kUGYzOSL0K5bDnzliNFs0jJJw5jV4/8X9inIZNrRJlOb33DWQ0REDnu76UPfnxFjzoG/9rV9O27M
EkVcEUY9jLQ7ZJWC9Q5b+Ba6ytkaVKAnLq1cb+dCEp4gmXjiGGnggdzu5DO/zMSReCjLZfnS5IWR
Bzq7MYiIiVTippfmDys7y0WpzoBUhyVy7OpqvRpkM1PHIqdgBiMWilDe08slFVZjsk6GZeVDfWf+
XjVnyTP/gN65Xpjl+34cLwfUFh/n4+DeHfSoce155VQBZS04RGEeJWQsBoAiFlB0C91eirJ0xl+8
38miFYk0/e9lOSkfa6Ek9tKrAJaXc366FN2AsgwGxiJg64qaPpg+SxRFEgjdEVEAOf0jImPb4qsY
AYcGB0WU5FoTQE3f2oE3M/5HAhNrr7dHyC6zTv+3QqLK4OGrgwg13Y4wmAbyx7THQWcYAW4fYQrf
/I6DROd6bPI3Am1HapiP8kQYyorCSqOTp5aMHgi48SW+L+RWQHLv1PqFr3iyzwcRWcs8B99wXQeV
DiU45CzxhYL4T3NqUGLgU/rrExedME9bHY9hjJX5FqBUYwDF88202VjWEmF+wfITsgB1B5oED5KQ
ECCpivBIS14fGTxtVzBvv1Twom4SA2sdyookg+aYuRAVJt0HCzdzprAZInGTpGhcQLcKq3BzwY8h
iEhz9XXYmz387oKn5v2HPowgLLkPZuBDhwYCaeqnpx7jM1U7EERNeMzMD/Mnz+TE3rPdgszPWjkY
8ZjmpaDpSokhS49mpJeh4T8+QM06rgjkO7NBzFkVJizGPE95vRCVZDwMI6xe9yb327v6/AE3b7/0
Iau5xD2zGrYGikiEuJmt5qf6sDZ80KPuUgztFmhWgTrXe5/PPjwBPD29JKQyBk0CHSVIKFm9QuHs
MZ9VrZsiXI+Uuhm6n3VpsUS4ycm3jPpHvOW9r5ncR94ukrZnJ8g9KYIwwnO0e48fJA+N3qEm7bVQ
jHxTY7huxb4q+CPUNz/eFvs3qpbxzKdyGm+3LFS8GFnDC7a0lFT1s7d1wW1CYwIVzB/8YKljy4fa
BOnGiPH0UVHNlM5pMLFe7BRrDe3+hC0oWxzosMk3VnSW4llmzClYk4UOGZRh0hCTowRlZHMO6Lv0
77F/YLE2FOq3Cgryuttd35EgGvzsxm6C5gy1ypLdBbPQyxFLKP39uKTiY6GIriHUEEqzWxW0pPYh
/LrqXEwkE8dEMhtjQjqQMjrzz58RiJAQU6Hx+3JZpPG0yMZ+V5wStNjhACJajwGE3pkBho28p/FP
7vH7RjzSBkU2Xq89+taheM4BF0ZqT6XM0gVU1Fo07CaH4OZjzGnsp5gnWvzWMBPpePbVTs7q/SOx
tYXF/LzpkEzO4nn+0nvQq4GyrjqI5NMfeBBtqB960RA6lQNibZ4JiF5FufV1sf+POUskO/bgr3NT
TGh3pIrxcWVRTvTNfSJKNXShN8x1CUYlHFviSflKg6az3BBnha7uCDQ5R+YjA2KITzllGvkn4F2Z
eo/YeOKWAFDXEtnWDTGFzPtNNMHQ5ofyScCwdUakbg5PlQo5JVCBb5w0Q6Au+PozpNM0L4ISxH16
o4NYPBqRNrJ09Je3I8y5m6vLaM8Z1qWkM/8EHV6Msxelp1DPJxZZlk9iqo6q1ZSrqwRihedBSUOG
bYN7cve8T9M/1GoackE7Zi2FWLdsJt441+rmMNGPSNDd5940kQNEARyFgax/4LJKaTKsE3EgdFST
U7AUap9JCBfj3k6HfTgkFjC+fBcNIQfoz9tKFlmnRAdrwmL/0i+xRlokedLZlXPYkDZlhzwUu769
cKTZt7pZOP/0BB/yn5BeQFjzOopXMoKmZmOoGQfEtGbGKbpUN0QPqsZSfAneynF0Ckx/sptkJDgp
vdZ2ju2jppApPT91VnK0yMs7pv8uDtN61eyBuMoqLHMRm4tnyBkCxuMOt0yYFrlKgiEhzrQJA6Gr
FFTC92uEIcAf5ZbKUZA37uMYEjxtjENJkhTTJ2El/XIFjstVib4CpGh3466igL6ProwEC+at24Wq
8i9BPljmV3KVMaZ+HQITKMWEt0gvncv0a62ZSF3mfONZAF7c/vgfrLuG/ZTloamdZwdMH6Dnn/OI
iEBaIUhzAkYVjzm/IWoIEO4l74GKwowS+BrIP5Np6CJSLdrhirGJKSjFMuHvvfljG2Wav5Lxyv0g
IXaME3ZBjoMTrxeXJUia0xG1QdSbNcvHQTYpVO1JxtZ2+K+YX9hcG/9eoiOqilJlhY07nuqEmOhu
tFR+KlnNwjqKxTJv6RzsY0fpv2hnzNyJnzLT412ejbRkFNRd0zQYH9q+L6Lr8PIxZrfg4Wu82lLk
4X8fLNBUJ3TVNX/Qk+iY9E8vlPY5o7yAtvZQIuuw4a0VaYAsq/S7muRNy+zK5V552IZ5edWJy0fG
6Y736UcDuTQBnl+Wa8CJcN2TFr/tBFnpnFxqoraTUjGfjTuWY+MIHwgkIyVLpQ8GRtZu1R/JlXy1
9julAoTvMEu2dR7qo2aydYQ3xtaCkp5+DOmiGuSxm2iyHicDAzMmwKcP8U/Ugo1sBigqEo0Am1B9
8dkt9HxM8yaNXIkPq7RQ/zt76WPY2J+sEjB+gzcF7pYI3AUitHC/vKppi8FImlv/szrEWxlrJl0z
RVnagD3rKLXRRVmcVx4tFD4hCjj47P39izGyp9fkJrpMstlmiyV7GaeFKKWUVoJPh5mMcJ8kb4vM
wFrypK3lJP1eIyj348AhiYuZhH7NuqVu1/Lx/IgmvpXKh+GOmcbJ6UU83ZRlJy4wsCOOLrXeN98b
E7gP32ZW5z42rDw+6Cm2thpKB76FvAaVcdc+tn8boiISrpZnwlsJ96d1GQrGnpqef5qLfFpOoGnZ
aGSPTsEJC0AfGWUuG+gtHYKCusDYivUOYpofEvUJB0TyFXCDvgNMDVnVbIBWcy4D0vky0dDcFJya
xRx5lLD9oihUwzE/uZ0o8rf78UMO1AH/SHoeeJ9IZmdpl+xt/X6p6uL+3gWXieLCQqj73FkQS8K3
6wfKVPko+mMKazPx+rbwt+L1N31KOqcPnwPWRA251PJU56k5zVaz/eDs2jUYES++5DjTmF2UpEUx
odVoco74RqdkvAHgjoYVxPXQZcfkSAIaJiic4C+9hmB1DAjlxDAeLWjDE0pKylt+fVDYZbGg0Dh5
2Xd6Fe7yOPd3/D2xZRpF0DZVdcmZjkPYx9XiVbS2FyibtQ8D2TCf10pNTHKedg8FCoKj/zyPqf78
Vv7bTO2xpxunke7zljfP34fTV0In1eABSc+808pcCryd95EMC/md5Jpi8tcUbYyLTROq1fvhbhxV
umaoWD7KHCQvRMuPDSuyuI5vg2WF5Ejy92B8gLvHS97g2J4+Gh5gtaWCVyH68rBmO7/GEF6zN20F
gotVfNSWmH9oTMfB846pAXIJod91e+MmbE36SmVweaFM5tjr6zTc2M5V2id82WCLpcNoa657vSDz
GjXfYMnhdhgwA/6DiqgncwRtdjcOwoadLLthTEw5YVj8IVA8h256ufZKD17J+NP9m1dmVN85C9ap
vueoXNF1phT61ZR7GBwIDYx2Gk8qgLeH5tCgxkjD494ZPxlNsg8YLv5ODM5UE0lDmLGLOm+ngEQN
yDf40TlkF5n/4MZDLaoqhc7P8YnqE0Rydx1r1weqFZMQkm52yWn3K0G6tSVCyZs1yo/MH5Ov/bMU
IFDGECudsUXE/+SOGzwCABXASeehLAP4aKW5HYnxpTJTBDe8HtbQupSG6m+KN3egEf+flzMN47ev
1wOGHA2CvpychuddingSAj5QXX9RDxc9cPuvI0mmjT/syKCUPvGmTVyWJ25Mtem6URbCsjqCgI7K
AZQJqaSymfFW8/gU+q2PsaEecsYm7/6SXz54eFSjcEQPpkFU2San7E8BMi/Ka7kRdULs84YoAHf9
1SF8P6ftP1wpITCNyUt1J8GZ4Zp2glHsxrTL3n/jqxMcmKunVnHcQjhIP9uJxG8AxOLHassmxSiU
x66u94J3AYucq1ZDmG0dpec9waLx/PZRM9lC1mLrYBbbl/YK0UfO3CZBeBdYk5jQj2YzuYQ8vy6r
KYW+MIZgg1JsZDRNHh/KG1a77xEHe/VNnYhj3310pXS5u7yBidUBEDuou0dTX5gG/UHGZ9gMEuc+
mXsQkm/jewwB7NQ0LxQQ/Ju5PmzH+PcGY8EwpoXOB3LPATYHRpW2z8T8/KNS6I4SrAsTJ7G1u8YW
VoW2M4cZNAq0hcH6fd0y3huAWqakiii/qN6G33koifLlsWzGwOoewqJJnUaVGYa3PauXoZV9C59H
g+A/iNRUl/UQiQHw7zcBfjF/K6jYQlG7z/nKkuVzO/3oWpn60rUqrHa+N5pRCXpsGtgs5ucPLhtM
9jlAjjoBvpV5ntErCGkkZiilQxs//rCkaBwoOleEpzHCRXmSkuT2Cfk1LqbyWbdhG3mQhf4zj15w
J1gDVWf1gyTeBUXLJkRxaboscx4Yznz7udZSkMnhd3pbx/mSmizFaqwNFSWJ2JHz3LLtO5J8yT9X
P5+q8OnTycsgjyn2EuI+Vb6lal2lx0XNpi4ZLB0n+OxlfXW5TZ/6IqDBQkiCHixFSb2NUR5bCW5f
Ov79iBvHKvRkjQpTBzfnKk6yOmCryHHxe0BoRMvpW99rfSR6ltiSxHW7fbXGoZdfH1G71GDknaTA
crenZEqR/nAuFLJp/+4Niztgvnhs11+xMu17fOqzJtLYFYZWTe1T8pJPFSwVkOy0JxsuV7fQdnqN
h33ppsnZEmK307a8JGKVfmSHUXso4flr6Q3XndG9P/POLgLOdBp46Zx+a1W3Ecu4yy3VmStvSd8X
rpbf1X0xi5mvCuUBPlzFf1C8eILDn2BBDM7DMLSLdBi0E+PMM/8IZMfvGaqzzI4mUzX198M40eif
BxltQtqFOV63kiTc/eYc0Q+ZXSIdvBEK0lLQPmly/czA1VhSJ3xhHUlWeK0CWiFSZM6j14YeEwF3
+MoPkfUFKhul9mWMUUrwH0HtpoRe1wiI2l9cnnTCmtEM6+7kvZesG+cuA39D8XZkOPL2J4oS0nGR
Nd524Gw36AB337pnt93HUXUnKk2S3EaXoGvE/aWVmiFyCD5ID8c7wqA3k7wdZ8MUfKLFA84pq2wb
D6qE/rCOAQ2S1PLzt9qXzkPwKG1cJtldgOhiPvsAPK6hVqvTjkhnb0VSfNzzxJSQCaJOv4nSlQ0J
2esCKclnEJALvDMrnQYAtleNvtGU4sKGaVxBSaoAeHWyzfrsDtFbbSu3npq+rBzsu2gr36EQyqun
tCuZfr92HQxAPo0TvgwfFYc1szjZjjd8v5kh3ADfJr6wU2C64tFUXkdDufRZ8p7tFDeAVPrw8VLH
OVcTAbJsm1U5m1SVe0wl4mLrZZcy814t1Rvh4zvG9/bTHrdzfNolR2rP0p+L8z3XGZChBpcQftOp
mjfjAy6vGq4NrQ8XFOeWIkS7hm0RLzlZpPsbKd4mjjDY/hHL5tkOfn1pk/DovBg4cNHiTRt1MTmM
yv1jbLevfdhtACurdWbBlhGpqAmxPBo68c8w1kipYEAl2hyShzSKnuMHpRedZKNK81RrIXryrY/n
GhiFram44ezzTIE6ybzyi5zwh8nUrVNNwUMNFelZCebVAk6AbKB3wcBZzrzL03anoykhrlK55oY+
E+gI+CRF8OisTa9AOV56nTXp0k2YzGS5KKCZ/70+WPFKLKA7b2H6jQr9AyFVHU2Fsm63hzQUlYeZ
9VAqrhnx+2xB35kiSKvbp0En3SUIXeg3v3XdBWEmk0wJcEcVu2nt29thaeYxjc/JI+Bzvk5Hn8rs
uf0uFMhALHDpoknMdTNyqMQXJLqq1vvnJnMy0hRJB3w/WZBmkGqnXs+mmQ6r6NsxVeh/Hk8vKvUu
9Ng1kJli1rCotQoTeXWolIDg2iQyd/X3BuehNSZbg7tYVslMp3vfM1L1N/2HUqgCUuLjjToewx6F
C3Y3e5bzVujLvViHsrBRoIh7jzOreLTZK0SmggFotqNsijIICecEjtkNr9dvxMf/urgjjtipLDTV
maCd2bzlPg44716vdNKgsZDS1wom44jETSKzfIjISktbS0NZ8toy8J+2hXoQcHh2xr4ORxgq7P8j
R4+Y6jBg3laKOBV6Uwufgfk1Md1iEBbfbnRhCP6gG6KPSt94nK1VtA6Tq/Z0uKFSNWNIVF/7Wyx4
f64MMc0j1owGfldEFsHi1Nffusz1zfHnRk534m2+BqaE85cwxxy4RB8ReplTT3FTuJm+00cZRSSN
qC0Ggfb4EpzGUb1bfx+EMODnCzYDhfI02Ty5nirO6P4aHRfkV05IObRYUdyWhMk6Qu9jpLNLsUtP
cx48fvGECTm5VjXS56o3leCDejFgd0uQBh5i0/BqovDJzIvKcQfL38OHm8TSZ3IXRi6FW7+zOEj4
i3/d6LBpTBKvRU5W5d8jfD/0EwKOglXPG4y+5ooR5tnSTgqzJVTuQveX9SwMHsW+soZXwyw0C3JO
vfTJjov1BxdwtBWsEI3y8EqxE8+1fUyt0hCnY1corYnJXRIbpuYXUtOP+eZ0klv7GgwQzQyNVfnE
/sIi2Ll42pXnTMkAzhbJTSJlm021Z0Ntr5ewahQzZmMMEfs48yE0RIWIkEEwxevQw5mjXd9S8Si6
OO7Su4q//EnAOfguMoMuKJEjIOJHbudCQxmCvxMCgoA2R03YeZWG1vRoVjopUCzrOxou76g9/hmk
/OWerFFKm6Rz7ILgBrQ3Sm+eQDMiXMlXCrg4GUE0Vi6qVIuBTpZ51Sn8Y9jdd2moIXKokqE2CeeZ
PbSLYLIEgKfUDkrZeGnEDhw8xGK6arB+TuNwgRXQ/r8TAMt3rD4PSr8cAVV9XKzvWm/JUwh99UaN
jWGotjiy0+k+o72jqNj76ivqjG0rbmqRhigugLOVfmcWVov3sRePZ4x+mTvEXVHB8fPfs3EclGN7
ZSOzurX9rlvMSdTb1UkDgsIIcgqDlcen3EQpj5+FR4Z2taMwIwJqfz5IXMZ+5x8qcWUb2u8m4wl1
+8JHJyKVOliAMUw+9/TFe7I42nP0CcX/mu4Deu+jcAXtaUkg230U/J20L8T7BHQFR7/xOl86zD3U
GWoOICmbrqfKYi/tm+Vgacf2usk/sduM63U2oLYJ6QaTbcNWh5VWVk3Gm2oDCilVq5Got2ZVT+rX
KWl9xXf1EyogpWxXGyKajAIdTjSuTtKH4WKezfPQ9CAusq9CHaYRcrCD/99Jv6VgrX9T6yq70BEa
u89I1kULRiPtsUD8uzGOdxD1s2OXvzzF9eYwmxOPrRpVLpJzhyTqdhxZ62SlzgF1t5ndwk17X2Vc
w4DVXmR4yvpm74vUVYekagx1j5SkSSS4wbpLp+UhWKSAVidSYXZJzvMXa79tFxQclLD6SyCSTy+H
hkUQvDACszv0B67thuDFHUtPG7hDmO0s2LtBmxPZQlU+LFJW1mqTQapjIWOeIhTRWmKnSaizqngz
cVaQhZW2NnKWpPdDKPQt5Sz5QjovsLJxP2WJ0ML4JaZNFkDC3WoGTVJ+YQuIs1zfs/GIQPSBAivs
6SDjAFo2gnrtmcF0Gh70am3ICfP2miPa725nArCWEZd0yeg2fgWk6GDCDTHB4H+jtblC5yq68RFi
r+4AVTOSIZfmvDbsnOmQLamyH7suLLBiKaee0HL0lcHHKw1Wm7eK9cIroF4frckAQG+Ghl40WDnE
ASDgnd1RZq4DbE7iLQ/MWeEpA7W2jrxk/Z87L5OltfgMl7//OYV6DAv+yWa9XcP0DW9l/H6BxfZ2
GnZkbTDhNIxg/BXuTkZwLtbIhe0UCjGqKhAOGxOOFR7TTmjOiNjJkBwMhnzVZiO9GjNZBl4wYOpm
32daQuOlKd/bbthHvTgRtK3x+jGJqnY5Iqtjo15o1WR7YjYWjT/fv0k+EWxSiqKZb4dhh8tcZHJk
HQzLb5JVKWSomBDFU3yeY9qnKMkxwgjg+uXFqg9AZeL/0EQptEy5tF79E/NVeeX82I6Ko0InZHFM
1hgSURELkQgK4daD26t0Qt7mml+hmLpOOlQDOO4BHhXAQUxb5ngngLwyB3T3ostJHRFMGbCD5Bzm
IvxNrOwA5hZKIwXsoA/gQ7eNjL7x+JJM4vW3JrQBJYvwrANEkufC4OUgYvcvrOlGJFn5VbnZhiNz
HnxjdB1MZy+IFhiYEgC12h+IcrHb/R1BSNR5P0VznXGog7ZyGgL3hX+BwjFUHZ0HaQq/WapVZroU
wTVuAyOT+JxClYi/T0pu5Ssibl5xcbALjCdpz+XkSHNLmFb1Tucd/Nz0STilADMIS6roNh0HsWri
pyz8okEHflAh9AFCFQHi4g5aaBAdFbDMbbh2+fuPndd5jTmILnnKl7HruT8yNJ89SYo+5BCg8Rt1
38/4HWn99Me+rL9IEFTLdhZFI0GDOJd/E1pyDtd7ltNMEIqXuZl3fiJatJCwpQxYHsSg6pYlfnY/
CG98SUZ+PQWquSf2aBgAJts6jo90kSlBSNQlQjiq4CG4yw9J7q4U46AKlH4fX7X/mk9q2phgoMLU
mu9WiPQionHeLiD1kDD2f0EUQisM064ERoOXyN9cqrDJNTZAEcgrnZ5uVz7uk1tj6gODdFLRg0BW
hKzT2T268La7mlFCjIwlJlboVAuz1YHspisDcrJxoIuM/mPKsN7DX60Smjq6gjUFHjMgnodLrSdj
wXdoURtok8djhWxzTCffFKF8SZ4x0uUv15Y7YODh7TMAujr9q7QntGk8BKuDfv2zqeLOHzMTKIpH
4oMlqUQGGXKDARZSl67Ru87FHfvR0eIVGpOsCv8gyO0nVgXEOgNOgoCf4jKRNjjIfssgYlzoaTIm
URJx/UDL96WSIx1jtgzG768jrlkwVdbdczSWZEkaeE0E3icHkGo5FLT+5RiPjl7+NbzNtqNA1uOZ
ARlk6is0APjQvaJnLHYs1CX1DkeODeqWIX5KmUsiZvB2sTJ3XdI2ScR93hd3cuE/a3OJooNSNwJD
JXtrVxKXLQcYQdN+svYaJo/AH4f6DsDgaTeZPFgu8sPMVVDA5RvCbK3Jfrdwo8at8MqqhT1490PU
QurAFqBBi/ZHF7AFkafjATcNN6CDjqo8ld4xJRclyC3xqUbMhxkEO1Ks/P7PJlKn/4lZw8An5uOg
jAbRDxGFsXWO949h5WzkBa5EUp/v3RqVwKa00qPpKCvO9kD+7BZ2kJLp1b24RbPuadPtXWGkuA/X
cG6uCW+nAWK1ul18r3kXYAkSJgre2sTfVGUYC10LjmPpKOpFzj+GqhrCnTeTp1P3O+Fm0R831uhL
gqC4PNj4Y1QSkT8QKOkOwvJhBNTbRie7+go9eSFLE5cl+ZdJmpcVZZu3ycVKTKvJF+qZBw6GzA/F
Wikif4qZYCQwWNyttiQRa+oX5Ib1Cc0d1UyxGWYknPU9UaVrBy37x/O9RDwpazvtMNKPexq23PoM
8sGEw0aiE9s1mrFr/1Eqsid0LNkh/3z7GlBxRYeKgbf037BRTCXlADkQkKjB/3MlMPBSU5VoKblm
V6GAffyMHLzg1h4vCvSXigbRE4cd9An1PkHSsqJhVDC90UFxUI82XtKgKAbI160Bf6RhRo9fEsQ7
aSvrgVqfl3x5OPwI5yqQrhGEFf17H/LnIaJ8EkI/ZpOcBb2W20d0ed/TPlv1aWUMtGZOGVB0w0AV
2GpsqINkq1kA2iDU8ruzwQ5jeGRQJZU5g2a6/S4EONm7w5kmKlyR4lsF7jy27tK8M189fz2XWKbm
RkJpQJQTpP5B6glnR0Z6E1yAwoFGqT8Y7zewaw2eW9q7nxudmcANqKPVvIBmaFOMYa3RF8s5NtGU
EQQ6aSrBkPN3wdKlmjVCH+afzAc/gqnO/iMS50bkJ1Kq3xfuE+HLbNuRwIO1eES6FX44aj2ddl2Y
csLvFeu+fLfGIoL7/kh55Tk0/xMac87AaBcwvKjNqDPssI7AxWDAI0MfCvVAputKe99yBcyxS71G
7VhQnL8G17LxhrIN+Ze0WEYsKN5J6drh0g4jN9sIY+Rks8lB0W6AWKfKcLSfgUj6VeDqwVxq9mBG
0yevxloeXJx+OSUhrNCmNSshiAhpC5xj+gkrGF0XrBXgGFo2kPnAwoFcPDLAo9yJ8j7XhcneQVHv
+12EiBHKvdjtkbbL3iFblguq/t6SMWjwyt4uqerh/BJ+5C9R7guG8s3rb1hNzvTUyYlF4eklJBzW
+HL0rHaSu0EF2sEqBSWlt4kJ+BGfj3oVOYQ7/WsgfrHqZP+3U62okPVauJ/xe5hh3cTRJsoyAusk
PB9c1I/X7LKTAeJrlhKfUyXkaYWIJiapybWyUh8t9CeCn4zvhu5sAlwc6TZHG1iKsH/tbQNBWwl2
iJJ6ivDb7k04Ma3hG/5TZECMZ0lZ+hp//iHbS68yLJdcNhDElim3JYzCFO2/qFIEBNcj8BGHQ4kS
pJaKxp55jWRvFgroGBQkLtqZ9eWUuD/UpgciSHYCc1EU295DAZYCdurO4XNVPSrHTx/XMEuAk9AZ
+jhXHzoSSh/7HCrHbsYd7sDhNzCcgllyaCYZez163eOQ3EcTQJx37aZtUg1YVWD9UAmc9JO+i49T
OTPlFpQk7P7MZiMnslmAW5n44v1uz7BRCG1ua4G0ZDNRggGygJ+oC6kDts7Nr5z0TsQ9mZGZr95j
Z4RwPSBIfag9yTBrmmTUoHCy/6xGrMIdNMJ+1xiGgEMLJ90YoLmah563DichPZlrLYQb38x2E1I1
quDFd+xnwfnkb7opNbB8CX3EGzAVv1JKdkU/qx5jZx37OhFib1vGkEka0ddZGnE5htA0WCM34xJQ
0NPzdyOG+9s7cxMYRB8pRdGkLBHbL1NQXriShJPPelyB5CFR9Y8fx98Ph+OOaCNWBINnSBjqRAWt
rNtiJ9OGuGE0DY0MMK2p3kB2/BRYfyXbRCLKoV4tpfgyEpF72hoK45ZrbDe0PS3LBcc4ALKAGWPD
m5hx9fm5PyEocnExGdLj7Fju3SxhV3cv35P+7zvt3I/kpM1pGzLUxk8Cljthr9AK9OKFllDcVa+S
rMuxgPArmtRj1qhnIDfl1p2nINvM1wNYg03JRouPEnW02klvdiX0Pjc+K9vTNoL+MexN0XHqGM4f
EdD1WOIP8KE+RauCTgyRopsKzu6j136yMJqtE0d8VpCsD+6MISrqWzS2+FFycCJ/Bo+MV9t4J+Iv
lArIhLU4GKI344R7YONXtJ9djUY/AnCeymv0eHMaL8IR+k//S78BtHvGcRr4mQiNV0/QOMi/qxKh
vXISQdZWBzq4E3UhcxsDirKavml38yYrebghOY14UkabYO7QjNKTk0GVNhqlWP4zDY+/bN5DOJFH
0ThUV5755F3rWlsRhC6ryLGDNcowz6UVs3UTcg4V0Sfq1CzV8Kh0c2jD/n1BTVAdpG6bhLMtjlDB
GL8gJDHrz77PJtC0JnKEQWKzfZ4gpuoKiyW5RzLh1EY59PWpNbuDrNNm7wYZ6y5fcDn7IfDWG4JM
wWA4xJuHgJFg34TdRnVQzag9lfEA3pqQbzLqq67CeplV8m0XsiJMwU2OuFw+PDwRpy757UbVd7uE
p5QdB/Xc9F3nx8wxsmfVq0UhlJYBuuH9SfWoOwA96lrc9t13ubMnxP4pvdr6w3D8PwMYHVvhlyOt
qynfGANSzd2Ohbz1zQaP4j+RcssiRwLIi3PRsUdw3VOL0NNhSjlngjosHYvyyrtq6wxnB9x+yvAw
dD3TxeATvc79Mlg6j0q/WWJtZUaWtgu44g6CdKFka0bMFisL6Dc4UvuLYWy3LvQl7IXgMrNUSuZx
PxVSYP9dKjzkNj5Hcfx80LbKtCrsDbbeBLzCIrv8LmSpKc3Jt8qplKh7Jf+UIw7P5wS01Yw7d3Qp
mfYLVyoVJc4mYgpVFSqHi1l6+oHv3MvQm/sOHq+5U4FdPYJC1OOep2zlkkiv1bbmQ/ZIrMr164/a
aD3imTiQbp1t721nb3PSZQG1N7ktxM+iZYmU7odlnmJPUnPSZ67OUUgi7V9RBwCb8SaUhOXOeg5+
XSnm5YZa7nuTjWeuU8MVKixsn+3pFHmXUwoehaekKbiiEXt5IJ4K35BN369A59b4Z7TH84nZw5QW
zo/PqsF0XYMvSz2OZ5EBW3Wmh+vIkezvQ/dWuTy3zBpi3D0sirTtPOdfhSs/LuC5MiALthrXcGC1
/eiZtLp7IgRiTxWyFbtDQeXSWICm2lnSr8UDvH0mijPBexfmaiWPajwUjRzD3naDLgwQ/j1/J/O3
8jlrDInamdrq7eQaG+JCCQPJ7Xx8HwWp6wqJ7USh9SHzkF3Kf1l5eoiQeMuw3HMnm70G7Xi3iGUR
1u3CIQ0wVALj/r4Yv2VKotR88yz2zX4SQwo7QCADk0CsTHBdwgFYgjnjaCtucKaD2wcn3GKrkL68
7Fk06G5dS3/9k6wvPeVymr8ga6HCrlCveI2Dby8+f7/kggapOlCU1iwsKhmRiNyLPHkbgLPl9zaa
P0uNLBymETF2q6Pw9yXGgAYd6Da4kj0gzuCPjUDpRfq9ela6f7vngUcBkstzL3vUdEeKOPGpnmlK
zx7h8fjOoJzXxMsd7kpsbYgAsRzSCWOuUihr7Kdb7Jexjzrn7GAZX833TsUT/joJN40eKXfbVTME
Fx5KSIhskQMX1EDv08Z+sKbGPgaeLui0briJLO7O9YtyIkxVyUbpY6hZvC/EMRTz1/S1V9lYLYXh
vbXxDFcXhXAsYk4Uj/ipMTHyT2Q6Wh1vQMQsIv1TyxAjtKlB/y7IPwfIXcbgyv7RPk0uVZCYIVPa
+iVCvX8f95+Ce6wNozbZrZOLd5xbnEbTH35qWzoVshV/hiodthLu4v4QpE6GoppudbTYH2JnzlCH
prpqlbofJZhFrqEgQQePycfdcJfxlue4kXNw5GuYSXOt2rn1EetRi6Hv1lUH0XxFrfRQyssW/N8v
k2ohh3hdXw7zk7ojIY17oaqXC1Q6P6gtJUdVjr4T2817CXYhDDWA0OLT9tGW5DItRhlwTRHCM0TI
NbREg2E4vsk+Sx+Qu73UOo8XI3IqL87Usla7jMZvPnR819ka9Nbg7FaO3VGC6BYuVq7UrUbfDAkS
pFFpc0scCnU0fXrLokhwzplCT1PulWDBnISLjoXeZw0K2rEiJUivtJW85iWb5h5JLfDnQFv/FfBn
etUQpaDbLwz7OcPO7zDa+ntpGh0+AbmH9vbRQh+0W0Ut8a6gJP13cWEOiKCVv3HU5tYKyFgA8Me/
WVGON9uwrEztrWKdueR940pcyZx1gkVND0DuhZAXFkIKknSL81axpOYtcuEgFP5LsGRKXLgsBb9T
w4ngK4BZHfXfoK9ssKtmvjdfiX8KXPQ2O40qSaYRSht0ED6AH1EjLkEHwVtCoQ0dULcyBq1U8rSG
SP0b5k0ftzKrfcA4tDOcW9/ZQh4PSQ5wswMR9tuSiE6G1M8OmpzXqgKIgzfTQIvNYtQptdUt8VBO
JxyhSNcNs2GGUwIuHRORKHwK2qi8OHv1ldX3Su+O9YHUzzfgGVFm/j/TurKkp0yGTZXj+7Y/PLft
rNrPzosgcx8xPdmGNSv6LZz2EdpzYNgHOvhgOUo+ss3KgVhqdfn/OuF0bJQTQqlZ8YLa7OSkKgcm
RrDEMfBygnJQgIct3MenQtW2+dT9KR2KYmpAIYl4oE+IINUkKWcMnPfiRnazqhb/U4RzSMqvWxjA
vxGi1U/Taj59M6tvFC8RV6y1/8yCmLhd/Uz7ba1JkceBY4CvUYsTe+73Ay0Mt75p/yMVB29XbZx+
/xa+dl+1KGMKVplV+2ra7A+C5tvl2GJ3Xc7Qam22Zzqz08wSF+jWp990eC/5/fZaMo20eHu5xI8a
7//OkIIJssJvo/bLggClA/9sTvV1sYx8BsCLF1v41CXRLFHqOz020r/h6ByWkmA9kUftr714B5Rf
+/3kfFilwUjsn5KCAwTNX5JUt5CvmZb1LOlAEQmlUZQO8+tn1EZ4jU75YeQjYMuAWhesVcaEorht
78M+kdufHRIk4pvKwcKoILf4h8PQBfv10XS42sKVdGm9ZuuPNwheuwpm+7IbH++6GYQG0ixiFOi+
GFCI5Ohyt2ur5y/ftCVYKi6svWSRQeqxYf8pjC7pboui/hFbjAWMbzZh4hGTOO/D7Ni+V1DCggZa
bH49hqU6+Jx7fu4kcrjsv5v/A7aSntyoA1S0gLK5MdTlSD7CjFGbVCoLUVUtVc0GsQ5WcmJKC3EN
iuuT+5FnaINPNDODrDEO34psL7dIoz88biR/9tSzU0N3eVOiAUIuVh9eRm/0gNIS/WIq4O1fTeAJ
bpLuCp8Qixp9+dZdv3AHboTKqm9z5DJ8+VfRK0xCEty0TAVhaJSTe2EPJqZQ+r/BFp9AdQMbTFU7
dZ5NWpI3gsy20DtK1SZbdFxvzMAsRmTeR2FqDD3YdwgHUPM24T1rJ7Y5hfdbMPLicJ/PCR2Qu8fL
OlbNZoWIuJhQUPRweCjmyLude6q/tISueSdmLc7A3rkE3kIGD910UzLF/skrwMztz3RsctGl4kdR
ADrR/aOQgG2cS9iya1vTIrvlbp5TpcBgBJwEqBEUOpWzG086grwjnJj7aDlQDdm5T1ezumUEdskF
Rgh47KJhQNwFlR+bDF0Yi8EV8Dw1KYuDbgr+e8a4lf0QO8AzWp/jzKauAP61iJzYG6FVRUvhji//
8Am62aafROObDiDfkUY40bimcBA2n4HVDT2+tFp/v5yFzTCO+aDOptPS5J1S87QZmpq0DUv7i+H2
ftGkUXrgvqJrg+3yiNd5XAiTxwLDgt+g0ALTZx5Pd3FV/S9YNqaB7xBrUSyicYRiaNnO/+a7obmG
xNc119CmrVIWO6A8iapvnVhIYAoT2FsXdGZveydzYquAaXZPCRJFubBT6GbNF46G2nLKWI9x40zp
0EfzAMrMXKDtkkwqhwr/TN54ma2kqG8q8MRV7j6fAifA2yHFhGXVrU6TXN7B+z5u9GGAN0ysAF69
lmTDLJ3wuiUhySiP6JWYlaH5S3qNusCQxHGM6anUv1FEFmGQ499wZXhHH9TveSKvOfrFhj5kB3D3
ATrRXS/LqbKd/zgrrE67vxS+cpZDFSIJjrjaEsVZasCfCAw8Vfa08nEACUmLxho6iL8gWmWrKsSX
jZskSNbiwohR8HCcqNnzlI6W2cVAPx0YhB6VCOYrVjxfa01rIH5AhH2aqxNwvdgRl8q3/hj/3m41
vCS7NLfEJ2lJ34jRJB78ZIhNQhCS9CRhCYYtVa17+VYQxNnawc7waJRlpXXGkJCEHH6oILB6MTYg
/brUIcWySSY+0sag3FblVTjUJQhrVqKr0jipBYstThQsf1HRVRn6MApTh/TX2FrSzsqQup+8YEIj
TSPmU3Bn7UnDtTYuPBnVG6DVd2fRxTy2Mkt184578X4zZIA7VbD0FTAMeq0yFhrS/xKTiSyOvKkt
gIclXtoL2sERBTnutaTEbTKXazZ38HA6PxoAO1ZiW5waEKVXVt4JFaKJg/w5c8be4jojXduLePvM
RGt9g8lfhB35YunyamRu9tkqEecvQFRen1hFYEPHnINxjqtbJgwpHfch7rrluFxxvS/Kw8VEGTNM
cJNxsJUE12K/y/R6yuFkSVqDyIDToTiXDNyHMUp+Xb2V7lUnF53nMbxL5Ho9JmVUi/WNYVW3nZ0w
LIbq89bigNE4DqMaa2G+p8o+t0r2z4fyWDSJY2cDnU6uslXJSqJPn1WYXYsqB+NJGcmO6KgzAXHd
ADewC7XAZt/kAolNdqy5ftsnLbdEYNeVpBeDntTsRkmJzzl2MN02I6V7iZYF1Zkg20r6K6V0nich
awNeIQ5nazwYmR9x+di32vGomi46YmWvdG+nVBb+TjMZQBSBE4bSrAWXhs1tLyGatWcZTUQaZEJd
fdqErxJPD5zYi/Da6NrwuSKGrnY9CmBzkW/tzHYCkaQ8T7zy2O+9a882b+6HOyf2e/GBZKIm43WO
ZKgSjN06MGI9ieeqlx3HQROYfB+hIEYEUgBfruS8P8gaMteFFzgp3sI2OR2LuFDUnDT6ii6qSVhL
3IvUoyVQrh+uCs4+1FmtaOZwUb3fpkaC7i+shOKayYqLgzNpMx1ktrwdfhn0wjhdlQHzU6xrBmgd
DRhEMH8L6NNq8vbOwKVCKcsS+LJTr64I/ojt/VxBZSDvonZ88FEJumPRaKzMylJAs2RMlQA8NQsq
p2OfTkyDQsN6D7/uju9ow7RA61bxFlkOL6nGd7FA6+82LhZoiwpTngxsWOQHRtDCqEiwtUFXM16y
aq0Jlwk/cf2eFKC6FPgR6Tg0gVcJlO5UHu8Y8LL9ec+baw4XrARZ7H6vqH92f/s9EBmhJ8X0uGPO
OlrNObpp/f6i/yiP/4fBPq8qOpnu6jpduruP6VqcLLAb+LJugzNprNGF+OeUjKzAGeCq/icquLEQ
DPZ/NTHID/TkmKBZucjqff5EDu9DnwZngZgrwxyfiJZbXtUAt0D04BodExfn/xvJq6p27cOC+Cf0
AB90BVZAoB24ob5W7IP70MuWJ0CFcpmjFzGyB46RGP8zO6jhvHxXRIQlIzGLr6k6cIMaAMt/gppS
1qFw2O05ywyiWmc9MU8Wvqst0R18XdDPk3/gBqpO8AszNeYqTvsaVy+mmqBfzs2OcaumBBiqSKD8
CQiuUkinOgJUpcl3KQcSZEY4jjQ+dNNOFniChDv00bM6Dhiqub6nVm35tavL62wcKYKxvOXDNiIr
iJyCQBQf1+EppzDNebYHoq9l/5CVYoBXskQVqgvVrIGFjSI91CZ79Ld5+TiAhlC3D9mtAI4yP+6h
2Uqd60z6RvlOvgdTZzy75pMllr93NXulC2eOJ6/gqJBLg6jbWNv0SesznGPJtYogTkIDYuw7fEzU
sE2E6te19fROYAH83m7MX7NRoxm33awTVryS68Bw6Z7szmrOxjoixteIWnL3Pp7OUY95NMfJmZ/E
kZmvIF7xKyBB2S6WvSIk0ygRrWiuCk41zQvjK9YxgLuFraUqyNXbjHmiXz3OKnD12briE3FZG2b+
YK95XPFKz7e42814lLh0k8kKKgC0o2vrytDwU0LNyI1aMTpYQqa6C21t8YsEI7UWB7DHInvzNnmr
pzNvM6Zdfv29Ycq0LiBpZFTf24ekux9MliMM//jXQl47PzbemxCOZvtEW1Gsz3f1/7XCQXRIu9aF
u51NMUM9auq9LnDAN12+Nzq1h7qfxiJAjqYBWl9d0WJ8Y06MZEOrkJel7Xdmjo0GPNfuzSFq/tIU
1ov67bv95d4vrOTSsXJArVr+fCXSGBLFQ+DaHlr3FMoXzQqNoZKIoFcjYqGiIN/iD+0EJ+tBR5Qy
j2VATiL59ppTs8Na85xItFZk+bLmQjcAk3eBxCAkQ+CgSnWTTWM7PtuNLB5PDMuHXqFyKiEfyxsJ
3HarYCRLUh7zXhBwDyUN+29b4xI9BnSUMCrLBJoF+PwrWu978dKuA5MKE02icHD0bjiM8Q7/xyrL
+W/R2h8ywaG/3P+EQkS6zhsKeAKwDBLk+EHtSMftJ5RJcGFhlPJpmKbHpoOzdCLFRJ8/PNag1uIU
4T7jiYNFH4RdONHg9Ct4Rn2qECN4alcQ0Srq0VO0FJcMs7T3DhN0GtYnJADGJf2veHfqH80n+6wB
aU/pU8FdhEg9CXLCSUJTtqjICph11fb5QhXcXNEoOJHYsqia1JIwQZSBwYYLOnMCxa4/iRD3FHFq
5iLuFhVdW/xLEQ0JSfVd05D15TJzH2rhPXDquvw43i7hW+P8LP4xrpo3ag11ShfFrh0jVea/NsTc
zQZ1u+8op22ZJkG3AfatTixNGCJI17TPSJ8WbJTbmqNxZ7t//J4B/hH38gXhqkdD53o+AZj22XKJ
oYqUK3V6nsY6/pZXPq85NNbM+zg8yFPaFfPXV9zgSSCkP0EP20+JZYat/OF6b94QhnMPG7bO43zL
1tv30aWA8Q6hfxL3Qtn0n79Y2ZNOf/vsOImR77EEO9UoTI3sSr8cGOuFdHkjvzORx1nu3cfpuXuH
qUYNPF5/JH+HYiJneR/HT1gQ9tuZaEy1fOw2YFa3xezhui/z1LkJw5Qh1R8YOKRS+iFmJwBzC2A7
k7sZ4ouRNtnGyTE3FHcyAYDb7gSA5NA28rToHDbVl2lg0HoIPnFkUy2grqy7INFLNY6pBPnOLpla
0DpO+trPbp2EV2sUPV+PBLaTnqzgSklErqyIWwJJn6WCurXXSEY3lLagwjJiEhuYFyW7O4xbqqrv
3DdAr+qkBKkzIoNy7QG2xzqO1cJ+tYcdT2ll2Bm6s2aMhvLoZJ2ofLUwmfnmZwaU4n4jI/MbOPDa
6QjluFgaRh1ndyxzE6Okwb8hAF0pqyZ3VCK7urZBwC5/+cIB5VaUxjodXlhI6JcnKqg6Sa2WZ4WY
i86kgmdNMnnuIxzms45UpGEPseAQwj0AKAqQ7i4aXeYdBcL7YGAuOuhyGaohTtfIMtPcoWQA6H3g
nRGIVBo2OM8tIohamCIrmRqERnDFGYrpnEYRNVN2pp+Mi7+h/WCzRVyT/zqW6hG0mKyl0l17S6ok
/GjoR9fnj/DHZiRXqgzYr/XLmXHn0ph4v1dTq2BcBf2JoSWpb1R+p4UXHrpqFoed7GEyx/kbHa7/
Fk06ud1LBSYVk8PzYGMTBsxfx/MEFzSyfG25vUnMSWth04eXFcGUGlVnq0BuwkV33FLxC7UKRDGr
VE1miYVoDEefZsCKJXSwbQ6qhVWqJiFQaR4INC7z/rFT22/+hteivMyLG9JxaWvjVVPKuAPlyRlz
GVtPjuWmxNa4gjckkjS2uFuZma6u5if6DFNzWO55BSuI/U0+sdBiLW0lBURmp9I+A19YPFTeuUWX
/LjDJyUiYVm+LqXQx85b/hqBVhwd/zSrvdb+2eaElCnyzDvhfKZppvqOGBG7/HJmrFnkkOMr/h7r
BCgh1NgjoFC9h3zvQVD8S534Rb8NEhl262Hv59QlfqN4QM9OFMzkhsultY4gUFDeNwyJOH9cjrVY
lliJWedo81Y8wnlsMt0ESktB2EatZD59KssMRHQ4imAhGfbNwPk51n+cKDO7UdnwkPm3cGTiEOkE
H9yBJHmSXu7anVcPijKSyWWalOUxaxSzfBV0FeP/P6TPV4qIu2xnJDNLQ7LPpB8EoW9vSdQ6Ucty
2rC0BwMWnNI01CV3vO9QlwjgcwF7bfQ27okdpAw85YXgk9uLFp/AHHhOA32uXmadBDFjKefXNnih
HOPqkBvNBMl9r4O6bipzdJVYVRXGEZQVDQxBEiWiORUKRhtbYS+x9gtl6DDpFjOVcO0tHi1uSFXi
4vQrULVjxtdlU9370V7m8u6G2qNoEv4XRg8Hu33gjEJVWxWv6L4YmRZk2bN/+XeYL4fC+/f0q6gA
ul/TJR5KjBAeNUVXRFmlZX6/K4nDUaTUN2wgP0AMjvGx8Q4qMxu4LFkO1Xjnixq77WnPpXPUSqOh
D2l6UEFkl5lNS483LsNcb6JI3IYN/Re/oGaktwBbLeFdG04JXOyPC3iinY4MAGTFd40m8ZfkmvC/
5NIP0GkV8ctc+4cGmKmHUi0hKF3sQC9km1HX56HSmyBGKiMHDUxE1wJUd2Kcnue28Pw4EXUR1QIr
mzv90YkKeIaANSytVMM4KaI54ovisIA3BzQKQV+TjieAzg3z6n6KBxf6i2/3jIfrRKIU8VQK7QaF
vF9mUQ+HMMX+v/TiHAcbgGuBXfJnn/2+GllEy+nTDlDSPjUXAHWz5QiTKe71/86YC+LT4jfI3Z/B
0GwauhuvQBOPsVTD/dLUBLRxGFAkcfxbYHAd4fJPzbEPVrqUasp52WrYh8I6CeRlzQGVVL4gfJaX
c+9X/YrKpQxpvi59Qix3sq9g/kHgKMPrwSBQJtKVICmMHWXo1Gz/SaoI3a3OuuA3frSIRBubTz3h
5fRJohRTpPL1zGlOk924bNNXiUMpaPx3RWYUaQb64q9IgQVn9lLaucB+aa1q6WZAgGzDzittNlo5
aHwnEBHBR0x21qk6rVzCsE8Llrss3Gyf6MQ+aO+FJKDUmb6VYRo+nEYXVoYJttTRaHCGQ5N1YfjB
/yPy5ZpkSpVPdz2k4ukhxyFZaN9+qZ6DQ2rMlGOLlq0HrEeAAc1Oa3VdI7uQeQnbieX9cgRuEvxX
9NXcsMk4M51R6iJjliclz5qGeXxkqwV6Ks83+XLDHQwmFHgDvVAjVZKK7/dYKOqNBbeUETH+fxiK
QkJ9kNdz7+py+qMAbZD+3Y3xdzRKLN1tCZPd+a3m6h8VCSMjl1vDcl4T0Yz9b9UImW4BTq5FPNWN
gGm/QV0y+eI0rvGRfnseVXBTth6f46qYjn7JCoOPlT0MH9F37op5rlDdd1A4Z48CTnaWeTpee/0V
7+Cr/tO0iUZ/SxgGmmfK0z+nocPR5560VY4J+fCxKXyBUop5ju2SOGYcsO3qoI0VkTw3GJqfagZV
39tgpJm3XMAlV6/LVAeWuMI3GRsUAM6sRPuNS0L5mWQIdfcwevmUY+28CqzRi55YN+TzATvGBhMi
GNx71C1EiIg9uxGRTrnLQoF2W373xHs4ubMcyAG3b5z92ljyy52D889aoRvwoJExMMmb/o1NjmqS
Re/D+IneyIeI8bOOKHkVNA+hqFcviY87NYOpmgnCxv30nkcmRlCJygWvPkieS8dgF9In4iIchfRM
YrXo9CR8cwuEggujkI4rh3ujQioxrwOzOe+oGQssPrGtqsEhMLji7CIV12Uss/XrxhP7GBHjQyEg
hEcIsgn06LV5qR0a20Xb/zm80zOjIlv96YELbIFLwbLGnksHIJvMmXbr5yATcuD28Aei1cqPA2za
tJgsGV+w5PzaFv+hueYNV7dka7tm7lndXhfjk/3WcJUfMpI0NdDYBxwGFWgCJPBMna6ChUxQJ7lz
rELKZJZ/elm5Y3yMugUoq+3rB8O0sifbGprji59NmwSd4tHOSICiMMU5X49BbH+03sdJZJBql+8T
lWKqrI/OWY/Pw22nT1zcfObvnyobTNdil54FsO+3kbRBOIYG73h5t6i8wDc4FoVb4JTtEnCWps+U
1F2GI2EMhxgwoAFs4XrB3P2uAjd+xu85jqiGAehpqTiAPXTByXVT43nVn0N/QWgRQMfkOjXIiNu5
QRnYTlx/j5/pp/ZJrWaILm9iJWmu93nkB3GXmxC5Lu4196ra0jBs0LslFNBFOJ6Ik6BbB7seAhxT
SJ4d1BF8j7GD3vmxXnUiSqQTUeiW4bL+a4Ui+DRsnlu5zX5cEXfEG7k7soEn+zDqEmGwDRtvwny2
mB43maT4bAsvNsxo7BUTdiRxlIUdCufV5ASz/rNlCpLj02kl1NMxxklK89TNYByb8AwWJnb+X/Ko
Usp9mBYsMxmgDyJIEERO198S/F9R8TGqXoQ0jZKiEMtsasbXJ+0GKePTpi01d2apw3i81ST2RDi4
N9DzC5YhUh/P4v7ig7wMQEtvhUbMj0V8J0Zi8F2iOfAV91DT7C82LlJ1pReQ0Rm1WpQNwGc/Y+yx
mUDLKq9GUSW/mt14YOgae0Bq9avac7/Ul0mFV79mukDXjcJtXxoFLEyKLXwrVopYoDbXE2BVL5MD
L1h6Gh6ebSzi4BjhO9wcUBNCZjHlubeDFxjBg1Akcl/rOCYloHBjfT86e0jK8wTWsX5A3KXs5I+m
2OnHmaPj3xhIhiSv5tS8TKiojlT2JZrxXnG+sZMm0wX9KXiy5N52s0uZbwdRi5PFYTVx4XtSgbWM
YKRm+qn42REi65XRkmYyF1r1GTDvfIiRrsKGXVg02jVEQoteFgNjM833IZjb7VYFJtQ4aAvhgS52
ITiqR7og5SN4bnMAVxgDN+IkdPkGbYzbfNNtXm8DJ3m26iZXBcN4CNnhxAGqURbAbIxuEEnHAPBT
bBtr6PdZiLme0gL3dpu5SogRkcAt83rL2RjKbpBnADENii+AfDV1//YcnATAYV0XjP+3A5AqMk1C
N7bXNpV/05RD55tTcFVN7AV61QqvOL6zU7zFl3Z30YTP0vUw4F40rCG+ZaZo8p+rZT3vhbrWcNJA
nsXKM72dZDY36cxVaaKA9q6uALI+hCuSwJ5h5TAryT/5z7IS1ZYSdW+fYQ8L/WDXZrIE5VkxikN9
OPMTRQ5QIKQdzkr4TFCNLl8EtPrSIJfwV0Sy9ztUweQA0/97bEsJJ6ej0KoYuZMuJIRa+9PaCGqb
p1iFSmT3ip1fQRvH1VI0PunoyDRJh7WBbdlfmP5wprAuGA+iYpNe70sOETrqA2lnJl65R0JAI02Z
q6HlmyYeBaIxu6ssnwQ9fIEZAurKf198npeMML7RZ1a4tDorTpFPZSxxEAM+KoGJZMlq/sNhJM84
DFalYg/cQ92dUw4ZBv/Ka5gZOlXhcUnusgcWDj9H5S6iPTPlwA+ghJRyPnwIkVQuinrewjcKAXdg
eIW7dOFh7sqjIppJEsnCsKiUFjFRyeGnw+nnhlV8FpG06WQ8CXU6x71u6sjNHWSRcw6RWHQ4227J
xpC6qA3MhBYGCCDvMHJGsPa7OGIIYKK7KumAgeP+EbHSdWZv+s/3AgN0MLX8lPFiWnMq4U/roqnx
5zZhJEBnOn3j+bxzk0mj0wDsHDe7giYpSjSVkCYiikiozLLZ23S4EnNZD07gjEQ+yTk1B90zW3TN
tH5mUxbtL35RJY1x+zLlBZGGPVMsVEGvYrOBSShaieUVNxlkwFuyd/oXlQE8EHBU3NNsi2Dtb6vF
pT4uQvRoL5nWMovbNTWuTjLRriJdHcwBp8Dv/b/RGo5ZxUd2ipGnBpQxZDKi28slEJ0EORTO0Lkz
IuAM/8nwmuQBxt5bCZ78iIpWRur6Rv+BEHq93ZhZUoR1CW2zxXHrdyS0MQ7ONzUCf5yOUfFZ8BUy
srHbSVMAv5F/Svd5ASvd1LxRHUkhYecmoAhvlVlRikZ8vSQXTWN3h/0S+ZiEi+ojZtOv+FIy4egu
K9tyLj+7BGIWqml4/QUFZQsU3SlnrVqRbNAPT9NpzY0sXaPnPps8fXa3lc3Js6Ec2ASa7W2s631H
NQRz0SfvRoOXjX3MT2x70aCXePJtCeRTEZNrv0U6kcVa++pawLgqqhg8tmyuJ44lk+0LresG45K1
cR3XsOe4d9xNcLCkxzVjIPhEU2+nT3PWEf+sCRKoodlUN+lTCgbxepVc4dfoNaGytaLnWbTCLrXj
AVw64D92wjYjOb+H3gkmD61f5/10b1JyLiLyddf+Ak3PM/ZVtk+fqh3BM1DtO2tN4XU2FD/bYiwV
Py0MW0+jivMNBS9OUZJqddFoH4O8js1UZJ2U3QTs2uY7DgDVAFwrodHmFLha6M++n4KoQURm7ys5
za+p9+YClW+q14OOcUyU28rhIGrkvA997ZM4gkouhaftQQTjsfkhEX/XIT4XRRaOFuema93+rfd9
gzUo1n4q59Mk6g3GoeD3PTMhKuHOyrzN8lqpJ3gWVzBKQ0KVHB7guFiDs8/PdB4zO6PLgdV9208C
fOxoAu2cgsWu8XwQPIpnmLss0qwPI5BLIksCbcyAUulmzs3kpENFEON4ndr/mVVgK2FvgASmEmfr
F0oxC771fEBtLCnwUkj8Si5inz3njtmd+S92K0AoR3QDkzhIF5Zs1hTbmHV/5fz+Htf7GytxcuTi
DSfF36blNJtkRM8xSu38YQ2ItiN4xfZBH8+e2svcPIcvLbyYOgglEVoWZITl02wVjnAps8Tb6Y5X
o5ZzBiGUOy8ICUVB13at5sZpRhuY0n4TAZN83MAOJrAdHBJLXEn2wCmqWHwMw28vZ8VXq0JcDQQq
cy17aBBml2oUeQ9hQGHaaBXwM8a2GfkvDDErC2eM2VGDx77CZxWagbOTctqswA1rr8y1SQkOY3Li
rLkv/sQ1dcs5T5TfNMF8D0x3KdZojmOTd2PXbOvwHnBZqbtmi2qEbRTlsCMlfiQTMIY2WEGU1Osh
BnM8l65yRqTcFyitdTNPKMwVFety2Lh87O8uX3tnsVZwF1y+Qnbg6DxPXyXN9k54pZ4c1t9TjrGW
bL+chkI0FQaIOGIat9I5h2SCryFQBRqqLgbnUWbsjC7lUORQPjOwzjG1ambm+LRGMUMfyG+EQMRR
w9WlllvHpLqKXgwO47oOBYhZpmUHt5SsBNAo+1DrlVtfmuHhtGWeOlexJ1VjXiaCZCvA/dF+n9pg
nhSpAJk6RCp4NvXKORIjYmL1O61vllV1yOeNW9X/fvTXbsBNscNyFP9P+uc/+YVMCm2PNZ/A7/Qw
jiGmK49V+VSEaHYvu146vBbwIMxhDXC8niwIaoltjnlWGaijdKsCI36v4YkP2Ndt51gldpPPxhki
M/0/VETWKDcnbIQ1FPrXrH4/lzmeoK2GJkeYDKGSyI4dc96KN3KHWcvLiplhtBmkqpLswvqbIlkG
UJUhM/yxizAn3TIxdjUKDF0uy5Cam6gfLsqUhqOzCfEYeXseYGJsk8gcYAMe/ltcqzSyTq4m2PjB
+QlKFbPXIEJPN9ZXYjxw073EN1++PMclYU978NFVLbhvqeCIOmw05A6YPGR8au/y+fwlfqLuFbmh
zAxSR3Qf4pxHJhWVUbysNmo0hpoNZEyEb7+YExnd4gqCgiNwdwCNku+/AIcMPd5y1zCVsrrKsPLm
mMVTp6y9l7cuqmHujv/J5VgkgPKg7pyxbJYYOnWctrUzAu+qVRCJC4e4OcUa/Wdxwll7fraJGL1V
jmTb6XI23nhD2Hh2d7MQ7eYKtqv3VaksvrwAGLsg7nVNCiPWvTY4OXfPay6gwzAqbZSQt/ke0ENX
PkS8p8pYZys5KSAXt/Y/QnW2ZbqmHBCOkUqIvLhWz03SEXSc5KVPnnmGUQbfIC4F7E5OPL+MDp/r
iE3KmHUm4tvtV6UX8kLXs/70IjHJI0+7le3i2QWXsRGtyxqA+Pq8WYr2MJIJ4noE/Qr7fR8fs2EE
wp1WTTEVS1AmGD+xHwm4BKoYjOAWKVEyhBvx9TbrSA6fgEPmUe855vep27vUAgfQl571CU3HNLWj
X5Oj5mYCQYsOC+qE/qPExpXKdFPU/DUuiHmzJGaIn4ueY9UlKjhKRW/0YEysI1nCu33GB+bBpTTZ
1Fw/6/d8zhzdx4PH6V5j5pDN6m6FvCHVWyu4IjPTTWm0uqH7PkCa0jnTyT6RPoCg6v9FwaUiAv/g
SlKPtG/rNmpzuBtg5vvXas+oLi3USbBJTljLr2IlIcwnHRTl/xCkg6usw9xsJcsTNHCsuee7ubj9
qxJVSEjVtwfiUibGcjUGonTp/xxOtKAG4gXpG6kpnNPCrqZdL8fnZ9c3rLNiPFQHVgtOO7X+I8q9
e8wmAarMxPwGitOC725YCFkJt/hqEHiSLfFzrqZz5EAmGLg6ru6GvPzvOqMbvcIIlWEvTzRTbRap
yCnz6ctwzVGSJergWhD9/gMjShZN+Ge9wuXQb67PpDNwBXA6JLf/P2714GMq9ilzHvTTT0Api5/i
ns4myMIwR+FOrcNnOkV6u1UpE12wnJIvD9/7YdbRFYhzsZnSICaksI7Z8QlD34btO+St2bG1fm5u
ZRIQ+U/0WS9Ph88nF3gfZ19E+UkWw1sgAXzDToMB8P3+d2ZtdkUNHLrNk8UHjm8ToaKjvuMheAbT
zBvsP+ypAUSqCjYvqo3vG5o7+uiiPNx1dCERrM/FkCLCSNWVSV1EpocXhFpRJ23S/BPM/g6YCbNS
U8SOLYQxVisqHZVTCWJfQNWFL1J5xo7Abnyr352H3wuxQ73InplpHv0vefBxgmTehmv9Zpx79iso
X4ajdFbsR3ZdkMXbmypRIrah/KwABYqn2eBDAnP+xXk1S/fTDqIo6dnalNhMxqYJALK+t6urkIM9
UF9EEFfSIX4L3G7a5HxfxeG7WI3v1PlzKNZg0CBCKKN1eSTEvxLqpMmCfBG3ec74Kiaozi77GUH2
DFDxgiHyRZ6AG7cg+Yruf/m7pQb8EDufYDJHSLCL67XQQ4ec3WLc5nvkuC/m9eXeicrTSp3sl1L6
sjJ/wEwzG5b6+HUuZC+RMN6gULk3FI2DgPakvJ1BjVPp7Gh7kvWJQXjEf6HGgk+sjF8t2xzFltYO
8MG6jGi93eM7lFjMbTVhW2B1wyCrWYulp0QF+6rhZfz6VsSCJWJ260p+kjiniF4zIplMRGDGy4A3
uXvfOXLi8BRt30S3Zboi6VzSVjCiTVBomPUbRu7/vtcLLvaB8kzImC/Jn3A3FSkHgXgT1O2sMInm
G7tuc82wzizAy6Va/BeJZ0PKHLskO14XL8zFs6p6CqWJZsoneVTsl+RqtW7PLrgH2P1MxpwwgJTH
rkEEY5FYc1MrkxHNLOQu4wMv56DFGaH1B+dKKQi5EBRgUQav9pUN+ygqXp4RuEhGg9bmL/26rC2l
ghhccFAC4gzWfyRrddzH1QQbJpNHjtpzrJkyTqciwspNki2FLl1y3PhWtMXv4JWxxKqS3j9WxONR
SWYrBgNnU/ojY4956E7wIV+mALu9sGXYp2WYhz1q9aPWrOKJ/sqomj8YLVeR21b4FQw9oY5OZd4L
Ukr3uIdmLhuka77EuLL+u7fizzCA77kIx40bFS7U7Inwpj8gjSd8v2bGPTDZyasFKK61WSFaiQLB
vJWSOlqTR1aaqCyrN1fqHhmO5OvOIaqXpqOwVsQhOadwmbQJ/d+pVPnPtcOeFzz5PzC/pwBPNj05
xCoPpoXf1M8ryeCZj+z4U88/ceFMs7OiJHcd1T84RgPvMwGsYnz0oybR7r3GLob8hy4HBXMomvt5
mR0a8TlqBD4EAcFujj/RXqwkNr6FaQXb9Gt7Mbpl8CFzCEQPu/6IU8OGAkI6TCbSs34egcX0ThB4
8sd4/RiIsmZkxFqI1E6/aZ9VB+8PKON8qubihPBgUj5y6zjLuiS793WPNI2h5oc/w4NZ9+UBjd7Q
4x6YqVafJyPfDnYtUh+cAeOn43Sg7rx3M+Hr1oXSw82hGd12fdxbWf8jU9MAWqltIhvXfoVSurqM
lGmYFlhmJjK7WP3IZyWTpiesZYkup7Jn8dyJrJN4RJVIko0aZNxnWik0VT1yt/uY84j6qVQ/akpq
67F+sB5XRrR1lw3B4qF13xdJpkGBCoKY6gHhiTwi57Vnx2OftiC6E+q8RPZvY8DS+Dy5XEmFAw52
Gqp09ahrFpI4Jd577pGzNZRnu78Nh8rnHPTGj+KjFJclxVISguSWvjwpNjI/sOHMMYkMONFCFb1Q
sKGfzeZzlkUnJmiBX18mYardxne6DyR5p5mrtmEUtmSGpsNbPUkw/v2TkXvsxj9+4yYD9E7ZvYB+
2dOJkSC/jRTE/QTPTr0V3JIKp+rMlgZDMgMHbkuhlLWFZ2FP8N9dpE1qBN8tlz/nLDhcqCEO7MKS
HaH1tF1Y6o71PNk2o1dYSAJj23gFlnOsD2vfYzcnLErWplqrP3Ghf8NwUWioei4DqHr/f8WYClCg
Pt1FjQI55OlReuDIINuEvThEL7QqIUB2gHdsypoTOtjWHTh4a4V2QTtmZqtslG2Guw7XKsL6FNAW
gNHc4DN1r8+nBGbKvD4HT3gy4hmO6pAt2m7Z/symrgI7bz01y7+nFEhbAcPnmLwg2pNXBcyOplkJ
dszHoS04ihO070mD4aj1ZxC/v5jNEgdaFRyfGczgdlMwSwJEePTCAzR3xpj6BqUs1F7yGR2Xx+ud
lSBGMkd4VwRI4QwBnY2ebeM76yafECeEm3WcmnjXcnfdPDInmznnmTjT82Hpi0qd7e8A/9+TY/I3
y0o584tAvHFtS/wCbgc2EBlOJyhPXFkpOXwupuU3NCPnH0F/Pv/4zaoPiFgjHo1AlEuM44LAHgrL
W+dGJzWhJnb4hbj7pVlFWLVjH+L4f8I0tJSpHY7eDhfp6TX9cYlmmC49DUtPPJGHqBndXFawSSBe
6EPM0zFH1cAihjBD5riCX44BebpaRS1gF3cF15QLSc4bMC0H3z59IBS9iXuMw7rKmRb//7bv4Hal
SN1w5N1LgGGdCjeUZAHvPaEwG/4qUJUzzB+K6koWDeIWtAYdZ7CzsUF4H0OEhJNk3K1IokF/+1y4
Q/QXdC1vFknDzyBw7SCB7ETM0GQMr44tYpfngf0yWjePWOJ4DAqzPyUUsL1tqBfXcc8azBkMRIlR
2dViJJXyz7076Cj78UsQhYLoPyQ2bjIoXEMkmkpc+b0sHaBkS+Q12jIAEoeOX+bNYHChG1voqic1
Kng42ivH4/ykt98nflRH35s7AM3OzHgkwtSGqkI4FwQsZAHyHyMyl66LNmZC73LyscGAd6pviW0g
fgpdSXcKO+pl5ciGbzR2sZQFptH9HLIDLM1KyLM72LkSf+tcQno0s7hf/v4ltq6Okv7M69CoYx77
Smw60g5c3qk3OeJVf3IR0j3HILcAbRVP9tDr4u5Autiue3gr0KevrGUNJ8RN8+nuvasNnQwBr8Jq
5z2P046e/xNB27TTCkFAHohF1O9vsbPdXrndcEtK3/103BPiQXvBYgLSFbnqvWlDE5HdeU3rXm73
JkmuYM2blQ3oY3+Z8LagO7KjeO9pkUQ8mrDBYuZeosQY8eDQOw1LaEhGv7W17Nsbg1Uzc8Z0yePe
iw4jl9TKkjYfW5OTOYeHCeAGXEaxGzFW8qTEZvT+mLwbtLDqKrNiLn79hoHJeqtpEeKV+OzDFpqn
1FBdXFsw1IMqwdmh2vw8iVKtyRzFR6GnznsqNL1CVodZp1FS620+4u5eMZBnxOyx7FdJoQzkiPeD
84zX7W3iwdumPn8cVIwTVbNCkU83cf8MTyDR5asEyS8P8zfbR5Sa8re8IWVdIw5JBMlzfgE4UVto
bpf6efFJZU0NqAHTWCJ+DiSUfxcW+SbwBJaqWH4aqORHhsYBE/F3XcehgVh7gWx+jKzQB55YuN+M
eQt/JcVmeJKUXBcOUdUoeAc7JT2dUOHNqldOAx95jc1aD+KAXgoG8NhOjqGnKPbzNKkNnUOka+UL
ArcsZNDU1gf6X+Rd7wK65+x1lwfT0p+zPno9OrdSMK/GsSAQUI4Ck/J69Y6784/08O8/h4W1tVAE
4ke7wD3Ud9rGKQ9duagntMkt+atcP1Ptk8T7ISR6exDNJUoZnynXNtIAzrYf+oDknMrSbDhGaDV2
JpYLLRNNnOeUVmXu44iYCDePwuItw5uxMtduZwLRzoFRe9kasTUsfVqgITWI+FrP/6OTocS+lHl7
/Jcn0AnNhEMOBNqZ81MEDgAiWjyKU6cvYtUbxPZSg9zckf1w+cnZ6gzlflBIZ/bd8xAZkTq5TEjq
nYo+3/wDW3ZPOXrtSJpT6CK0qIPm3afSTe48vNy7ERQDg3OqZanJNettW1hDKABkVJS19QzE54hq
4hgu1Saf0EcIXaNsn5iMvaoKGId+y1rjXfJawnqltS3VsvI4uX1g+dAKzpe1B4jDUg2Qu4/QcOWp
bA3yhKDWNzABNmyRqNACe20wIhmSSi2EQ1lpsLnDiAaXnmB8K4B7Gfnp+7T9TNx2RWHrs9PKineD
26E+mb3E/oxhw3I13eRf6zTTPqHXkUcPBHSvWysFnqX0nndudDtwzAwskU+GNYT5nsk2yU0zN89v
n9/Asg5o91NSsO7U6dB3Conir2MEA9r4WmeMp5JpPZKlDZ9sQIzCk117xRvCQsTQqvMGj9bStQnq
9EeI0u7UbMYTFanRZVDGmww5UEZnBpvURoz3BWE2dDxghP1IRxXsflVPz8UNaImqaR0oQjT+uqUo
6AX+0Wdd47cqRESVsS+dQ0oPHH+/jmg7TymGx/UivIVtq6JCKa3kF24hVp0uuvKF9cGaxHCZU9yz
19Gfa4vhzPxASIoV9SbsUHX9qEiLfPCZ6wQsyr4M87heDgBOh9sp0cFep2UPB54J3tOdSYeWbVut
zoLF5rnSugrHcboPSSuQ3dQ4n2FcwGKucO8j055N0KOPhyPaR0zi0qXDY3AuDYk5QQX3DgA0vEez
aCo8UiK1iT7dkAvJeKodHpjj2PXdu/P/dbye3dWHRPBDqdEJy8bNBPBGHHNWleKUZo9DF5C0sHOl
svauxwrt4Cjq4gtIz7PwqowosNcPebWpDE5ub1ySBm1kRWUQUDrctbxiOfG14JWbvY+lhR6Vu80a
ThaDDIKhBNG3PF1beJYFJdATvtNmvr055y+DBSUMI7ygS5aE+dZ94MuS7ohqTJJbSl9DHEaEvItH
CaF8lKeBh14MNWfHTpS2L9Ejtj/M98m4k5gGhtAwtkJrFwEq/tg3iwmOz5JSfui99FgONPiJlLFu
3MxWxPsgtTgc9z9luwZMmroKAgT6XV6/tVHTQFSYel5oL7iOu8MaDa0GT/Fc9msYplpB7quz/obR
KN1PSJoNgSzxU7HiHaOFTEDAkA4I8GQeIJOPn3UdYDTu8WPJVKc0muKvWuiVgSNhdPUAugJKXcTt
VnmLR+D/FvJ2VUqoiAkYIYREYLGJbFBTEC9JqfP22/vUkyeaQb6FfSPLAu5HrakXLaxpBqskq/2z
YQ3en5wI/bYqSHVpLHZ7yRM05VqRf+BCdvAf+fk7JWrNedFZKb4Dhqb7M9M2MJManzQDgh+B1CbA
wAMwRbBiNJrMuQV78xlDvgkSCtBijvTHmzn9evkVch0N76tEU0JUcXOjBPyOzy7UFngFx2JTxNJA
OWMTfWS8Vzn5+AoragTYkfFpW6K5fkRegSA5ZDeQsamB3BXn1ItBjNoNsYJTOL6f28bnn+HcdMTD
gLBRz3xP8M+LeiuW5k/5byNec3Clmdq4UEfimPL4iqIy7FQ3b2qIcgaT+55T2mmqEFqoOgESc9/H
wBnRH4VDQ2J8unDHW+2DayGy1st3/B1Sgl1ogsHa9z+slCkPC844z7V3Cub26yWs8w9DY35jyz8A
NOjnRVgEh/slDshRuzQx6IJPnpHoJdjY2bsppia5Cjvzp2jrh/X8QzPr7Mv4PLLjbgVzRSohNLV8
wYTDiJUqgmezZIDg1SZNqcNwDwgoIWqFJV+rii9n4g8uDloLW9J3wrxXMXhq95Z90+Ne6JWUEQB6
Lq5KCQsEEBLdZC4YF9nP3MA3MXw6kMAwdQ8zE6FUfeZxgXVIMOnlJpDBltwygu8wl06xVbePM7/N
E9M2V/3YMpz5ekNYD7cSx4NZ4Hf+wCsddRKgIe215bHmLToh/TxYPDo4qIyzB3pZH8qBV2KiXPRo
tH2gFMSfnAdh89p7n9BdKUeyj1vgmXU2Vi9QMgRaqNEJVnrZnOgsti7aayxPLKmI7vYjKHYxRUWQ
5ENNNPSASR6l+tjYkxHGTCINkXCgpVoVenL6fgca0KH4Tj1ef5zR7urKM4MwEZn5ugeA2ysM8Dq0
jOFPkBCV7uSx2OyInZBtfMWRZ4Nc5u4S8lkRgF1vQze1VbmK1yKdlFKORz4PbEROa1krYmU5ZNIh
Jo1y2vh5ZMHp4s+gI9Fd5zwolLf10IDhZDj/oKvXzITaGGbpEyHTlPn24mL6AK9kMPsCzhm08BEQ
wzLTeL0hKh6qtW/d6EI/BNeLx/OfeIE4RkXUvCz29eaaPpIXCJsJxoNdL2SBoUO0zlPO98RYvu6H
b73x1oi5SrDnGj/B3G7Imu8uKIrQvJw13od6jLPs55BOIiH1cW/44FUmhWaV2pb/dFhTyDUzaT2X
TfDq5uEMV4o1FmVZq2wb/MssT+bkf+60HWDB/nHvwa1nruLhnHtYKtikZoNQnmoHH3ucwai04eqi
j0i5MgEao0/vK/jJf2633WJVQelqhsEfJJqajX7hcS0HcqksqEi1nwHd7RAhCPMEvzhYuE77f942
iXW82rjzAwy9eQbJ8+B+6+xuW0NOVfQdy/aghh6+n1WSp2P04t2MKOHf7hc/Bo3OACANBsgUo7oI
6Ig2kpVDJt2hMzup2X663RI/0/aWTW1T0AvPpJBcd3Kr37K7p3TTiPtWMvm1eBP1cblLztxASVpu
SVl9f+/Pw9KyfuSHhIvYfmSKHvPVsMixsEOc73FENOG/SFWiSudRtp0fv6pk5C0UgUjh+NUMyWwI
8PP2evUUWSh17OP2KMPcIVWADXqwI6LThuuR7RjsyKfBVsk6oGG1nrjkOmbgpAACZ4RMCLxPlfnE
eJDzbkvkNmPES4B9eOBod1YZOC4FWu9nq7fhVCJVpr2F27nG8i4c2VbUPlTw9FY8dHGSqhYblFKS
8N64fwJXhhI4cvFW14DGBNrkj7L5tBLnoKqLp0fOGJReRfEa8Wd8fidQ/QWlsdIB5Sro3BEQ5Z4h
weOaWkrEcJ6zL4oMUQkxgtS1UltX09f3AzNQ7QiiAd22XopALGCR0YUke+5O+ODnTJ0muBxdKXt9
qeB9fCttS2blF5+aWXNZJ4xn8JBVHeDbYd/EY5zejaKSJujnIrTvNxQbigSnaZ88drRijyAsZKTu
cHnEf8eS+AtM9guXl3uNc01tkUWr0uLqZp6/OTd+/nZHL9rALjJoVMDrQUUNfR8x/u5bAzsCRWHt
SjgYpX4BzeHjcgCTAVdsAvtllV+9Ii8lY9zCfHbkK+S4EMa4kdcFK5pIi7FDAmqLppgCY009Va0t
dNiL9MR8G0dIePD73W41AHBpAxxbtRP+PiNXrxK1slXNf/TUpyfvBW0LWhsGRH9H5kbIcc9fU5Le
ZhGxTg34haigtSY22zCSM5RAoparQJfjnPFaMI1qp3r9UqZDfsDqQ9OqYx2EbbYh4h4OdT7Zz5os
acKzoykIwycvITb4jG8pdOZj3jodgKBSLgnF/8OFa8icUnj8kgZfgPOQ3ziiYJKMu+0TzQtBQLRs
puOMHrjsUXEnd8htS5C58LgaSYn0qDNp8msF5AFOZmqtYd9l7ANyXFS1eO2EQPRswHVrrQY8NtSZ
N4qpxmuMnQvoVN5aCQn38qhwre1hlVp+0UPH0awmQ07KZlmUHafTXq8DHzLwkngRtmLUzQiu2imE
31W4Vng4DtaIYwQ71nq7S+nend0cVk5WeEHZo2K4S6+YJVLpgSQEcaeWgXf1gdkqnPF5ISnzm62n
dwTR1Z7mdAJ95PEYhfHeURPorad5ZQkFFlyTDQq9mJOMl51u4MejCN29ldtItQfclTBzPwsta18U
Mu9zIy/ADcvjQGTyW7SuWKQPyG2w4tnbyd2W8UjAuD+WmnHMMu1sWJ06ir6MSPrtMDtXjs0zBSpO
q1X+gCzRHqZVXePciCHPrN9GgpxtiF2BJHKBWxCpSJj6ZKBe5nGzVUbmlugaHvCQgfSUK2T9eabQ
5Qjw3Wflr/0MuGXGDz5QVwI/kiLhLJe15SQ3UEkwlVmg8tPjor0oU4UVm+x5Z7U1MoveGQcAGwyv
3cehIEHZWRksXxsn6UagXB/B0lYL92urf0O4LNhgbaWSnuJ79lEHkUZ6F4cdZtvE9aCSJSZaHywc
LMVnYAgZrJkodTHzchlbf0XGDI7UWjr2Ci65cBTY+Zl6fs/auXmgEqZOLZwM/1Do4b84vSkjSr+P
FHYokM7EMSQQStqb+BHkjby5aTh7UTu/bVWaifA1nVGSeC3jzzs+I6LIkdQ9knaof0YPMb7Vf40h
DahS3BoWJ4olk+MJyIjy7Z6nHhdra/pWHXD4G03+PUQoe3th0D9jqqrpYNaEbFxyxDaOK+BbYnJ7
qORdzhEbIq0WRy4LyymZR8w/KeoqXfiT0ooH5quWNfxZAS+VOGSUXzsQZZ5CaMMZO8dbooSJyvUo
hd5o+X9lqQi5i6AFHaLzrwLvhursJa6Lhb8JdvkvsjawVrAurb9jUGG5Oj1HWGRKFowoc3SFe1GJ
8URQo5U3aKbbY5FLBJ9M7eIjKoS1zpGRLmF5/vprb1895u36HFh6rCaQg+DEOjA1BnRrHuJCBj7j
gbAJ7Xmcsb4amkX0PRF2+9NJ5TNqxi9rKnWXwokqg/37ZSWeqmnheztvfs4Ia+CKbOgRLtB4cDiH
9lD8GRrou2WJN4pnYVsj1lACWxYNzb0yskXX+aJ2tcJ3abrl6Dyl3Pl+/wjnyLZX7y1SVokDbXR0
2FcIbB0nbaJIQzTpQFVr0YRwtkXccRUkxe9Is50YPALqXTLZ4x2SjqPDFOjhAaxJc8zjpso9uSDC
BcmZxj8ikXZEMEJo45xF7NWG5Mq1olYutZMdiqh6TG0ztHX6Sqk9ol9oWRAhT2psjQdU0ZTv+x3H
Z1ialb6dNRp93nJLyRsQw5EBOTPWUSl7js/3VmEh19gl+QfrXkIimmXAphyZ/MfO2xpt+PLlZHnd
m4s/acvg0VbRPCjfBwJqOE2WjLoRMj231KN2uwXoQoDd/rxHq7zz4mdGXmPe3pEKEjqdQh1t8h/w
HasOQgyFG7ta/QlzHeFibMleyZc+JJkoTQkKxcfKZl1H2Pe+Bn4YMh2o2xO5I8tqx9E1JpdBcURU
XAtuvcaArZjJCRLKozKAUvSBRhhKR7brx8gTbMfLNUuh9UFE4noVjnu4QV51Jtoxn5uqNuzFjfGp
cPlDNTjz0J77dzV/ABfVgncpud31rCt2zV3pbupD7V1HBaAdhsMV+7OY4cKMBB0nR/mtb0Buwll9
rDHsvIk5Cn6OPji6+zp8Z7Uepa4umBLbgWZfCSbk/uGmo/mcs7VyCjKBwtDaN+MdquHxBeif3Szc
XbqMk+jHdi0qidloUKlDKQCBNQDM2X2HKRp/4ih+xwdVgLhDHpXQI443/wObZ4dWhwTpC8IS9WEK
jM8Y6oSYUpySkuQm9qOdnAf8DdCevLyyZ3b5UoFQAEdz9PrvSP4ubvx8EuNhxsNGkn2afTNYLZgB
Zpo9vWUBJrrZm5bPU+zhgF33jRJKIVOCTtgqDVzYS1iTpdoY1jWoD7bICqFMVCqoixzu9gXeI+Mv
PB1VDSQRyCot1JzMAq6ukx094/W/sCJJE4F6Wh4Zb4AB2SNyvS436FSXvupmcveB1bYjkXSCAGoN
NN+TUJigWiQdFqfsNAT8l6DsdhOU4kZU9jPZuMvGKgvBEAmaCyH8fI7e9ajkkAjceoLCO4l1VmGp
vI2snxNjsJTqsZBjklUD+N4ZcgS/osbvicrTP4x44lipPjqlPfiwmk/M8D27ow3fRHkWy0C3CdhW
aoBBW5LH7dPaCzoC8EJFr6AOhgwIqfKRyvuuZ4f5h+alhO63ISIY3ORkI7x2vDrVj+aLivxSF+RK
mN58UTCaK9UPK7JtgKTtNfMYAcdcJDu8rXPLgrOIe6CiVeD6qWLsfGbp+jZ9EeBBgz0FAxfoZP3M
2DORGWKthK420WjZ7G+7GBA9Wv+Bcregrovgge7oAdpNjIEVoZz+8srxxPdRQWLGE5bPSsrwu0jT
CkjJGv4ZtdVC9ZxeZB60W9uNvppxs6AhuMHIVpohaJM5esGPIJkl9FX3agzFcTxTLkDmBGILRdNj
3IdK3WR48MspWXnpGlYzNJNRPlixg/UTwGVb8oP8KQJIa+nixAww/htIouB1mCMe3KRiDD7h4dMi
DFItvPj2o8cTFSQdzz7FfhJy3FE4/J5f8zkO9tD6nlokkUBUTGO68KsqdfL2xrxGRHaTlw0l2olN
IYbiZtsTvCVJLZEcHtnEhyzihXoiLbx3wdH3t0/4u6oNs9qQwylwdG2AZA5r0voHz/Xv4msRV6/N
Qk1VOXrXjCTSVYRwdRYDVs9tzrTmc6G1qOhIolqxbdNa0PTefDGTbu+1vWbLBk1mGoqLpNgrkrS1
4jivmnuKVUvawxIh9vB2EZnKJAWjIkWTrbn9zEKXpEQlyR17G5xdKNoJ0y5ly5+E67WSvVJaXAJL
bkSz5YtW/7nUdyPiP2m+uS6momMNbDvWbQA/Wzqpf4d8g0o1ydm/vFWMUUEnvyK0Qyd5MktW9PJd
OgcwFmVLKXK6MdO6wn5AkMyZgnJIHCpk5L1aFkfq+I6I74H1YjjBTOmQ4TPwwn4Ajy0S3Jsy7Uum
6TK4cQQYvN9+NdUK9jEoz2m4fe9/7s+aElJGwQMMNrKoxJm84Cd8fimrSzpdOhsn7aqzIR154cz6
8PeJFLGv57uj/wUrufzDis/WGBS4FLe5i/4NSUCtXbMPRKYtjYHXpjEHVRavN/Lm0B+liYzWaHuO
Vdn7n+4xKMfAtFAYTyTny6S/BuClO+tkMI9azWF3aqhy8U0jVr+dhb1BeOzQ3yE6zi5paAJkDvin
nl9YBZ5C9WSXY7f6TL4rerSOLT6ycBu9LpRqms88uWjA/Cv3XsHraYIlUgyCgwCdvaWX7MCpM0hi
LkvjWtWssrwyPqZPqoxkxC5bEa4+G7QD0SJrjtPbO6N95Nn/3XSQW5sw6cNWk3+GS9Z9o3IdaUAg
6k7W1gSwx2rer+0Ex/B49T3HvDXwscv7LypVheXM7Ft9YHlbcy0y2O3zkudozFGBaAYMs5geRnUx
hyh2FSEAUuo93pqSpXoNFeUPXWcOtjM7sY/+8EWh91Sun6Ql1sn3H/A4EhN11haC1aCw+xzQlcXe
+OeyHNxNmzZZond4PU8xfflMnqyrxFIiR8jOPUs0yOIUHtEHxsDy6X6nYKIgPtnMp59bWe2DEDYv
OCFph+Iygf1VLZSLjb4JQTFcw7A2hspvDNH9VoGWbsRFLMnMjL3AnnXwt1S1sC9If0co3VFVy5zu
5C2ZcAYLETA3QmZ3elNv0sAJfJ9gHRYnTvEsJS4tyge6ODYLhkF6fbFkznrsqOfBTPT3nE1YU8Xc
x4H7GAiFh1B8cBD4qLSOW73qN97FhsmjKudsS5vXvgzQdKn6FcbgdzJG+S2zYXccE4+HrxKw9BfA
/xaSrR4EUX+AVLVblekLehU2S9c8cvc1tVSHElp8Pei7SdELWq+bpYTZqPMmCO090Z7cz2kMGfI2
kIXe8mOaMEA4nP0CxfZy0bO9U8uR1d3gtNemwejKgAgn3ZM7wmzJ7ZyPQnA2Z2f7tNa6IWA9bs+9
k1IslvbGDjuLBpRLDH49MY6eeScl+McupY7suP7dAvLCPuqX8n0mrwVo+Pcrnbuf3PlgUWbT2Hyl
AoE2xV14FQEQQs5dxNzxeMkfB2A6uPrvr+A9crzxCzmx2EPGKJhAy/AAfxmytziCEn9E6YX9I36z
OfmAw7ERERSYN8yXybaSrPPWTTKT7quigjsihmDWyoZMbZz7W0+AfAeYYQ/6BrhfMVthHR4NMGj2
lw7KlFefew4YURyteVf1xP+xmFX0PJCwZlaXqmwkShY8IUX4vdZGQO6rfvJedI8GfV4YXup+Qk2r
lCQyI2bSMOaa4PfS5qA1ZYlaINxCJySq+SD0yya9M+gbyLpurUfcBbHxugwOqOBFrCAtRnYLWr/9
SS6vU9diTD9yJUugMn24kk/m63kyj6DfmCkuzXqx6S1umLJMEDuoEHf3V5jZNYp7Vng+YzMk04Q0
fWARtl+DAFwBz87r4B5JDvFslpskToYNCKIts73ZvDFBIxBHFp0WJznJaSDrQMP8oYfCAowa8ZPU
CmSz1JOaxU7G6cGGzkkAsvImwRiwYiU+ZcKTRcKlDBQt5iUAgBmkZw2gDn3WyjKm7RnZFoGAKRA9
6Xmt3Zap8eal03yuUYMFZoM1oQ6xaRHBJ9hRN9KGRnTKXijucmKYUaSxnC4C2fmoRxo7bUPnOcAj
Qfqu7Za0M4QUyZC8173lfAklb80B6zg+NbBkXMgBdiQhwLN2Ntiln8D5QBvpLlVfiAqrJK0ChgTE
CJeSnQvWdUtWIK1Lx2UJivoXmvUE5YNmXwBwOW3fvXBKtObBqG/pBLp1hC95WkltoX2vMdhXiSjq
/MUAdynljXj/ATMd2nLewCVclr106/E/pIdkvh/oPSkr0TJ5yPlLdOwPWj7PLPCwKlOx2mCLqrZt
HjPWJIiUbBIjjHfFxQDoMo3vNCt/eIA+UNAzQJc1EPOknMV7xQ6pkX/IYLuPa1dSA0j0tchTv8LZ
ydhi4cSKrYegJaalV4xEIktfGtNBvR9kpjXLO+uUCh5FX3yJOwEPXQ/K4SpnASXRSoazXe9YaEkB
Uw30OQ2cDrhSXT04DhnN282CaxOey8PsgrBqZLUSDfqYaqgC3pXU+XFU145O6igrZd4SFGNGItLz
oahDenFJ45l18sG+dTXLYnj1o5ApX+fbf4FmbOIJUKgG3XCHGRPpaIo07VTWvTH3JF3atIR8gCf3
YK5f++sF3ToeFf393eB+dnfZAYPZX+GGwSvzYnxf+oF/9HPkON2Itr/Cq+tj150BoYOA0miCpwJi
kTLOqBm4V3Bvsp+rajQbWaJacpO1clfgd636mgEs0R7iRKkzvs2+I2wwEEAqr8Q71ZZ7DI+asV5F
3vUfzV9o0QQat0iDsIzVjun308w92+taBF8wHHnJJKBJpf9lAIUPZl2f6Ht+040XnEqZ2828m9IO
o80F94FOW27PN34l5jixqTesq+wpSJqbWH/H/ECRkFiAiWA4/vmL8dYiM/nVfby6xad3R7K8uKrm
9JsC4NnDaB3zI2T+H8s/4cqwqAMbA717ba96vKIRE32odEPeMycrD+hRLIdpY29sstJiY6jaK6ax
ZVLPI8dPhdubJlKoSwrx06b7wJ5Oc7tVF7Tzj7g7ByLNkJCLD02Q4MlnaJKVvklk4nPctt3o96X3
J/Ubrwmtfinw0D8y8pYSvJSiLKvTX5mYFxcx92TtgxmqtBZRezizbUTJNxLX58aIOxHdAMp6RZ/k
GHvI8PsH/3UDeYFVQwj9sFUr4fHQC4x1h2fJcLybHR3Gypie5+d+xajv2JtWF4svCAfz0Ds8OYGw
vD2eLDX1ODO1xlOl06FHd4HrbIoCE+Urah2DZfcs188JNtYYpzh9JyE4nqqBcu5W32oJd+kGkXHe
yqjTIir1xfLXX/yI0lFCYQrjEMHOoM6rsFn5cW4rBQ/Pqfo3stfqeu6CKrFwhv6lho6hm+Qfl24l
gPaPe6KrIHIt3jTIYfKBCIQR4TeliCFmaqFpyMJcvwacM3Es/aaES8jsj+XrjR7XFNLf1+ruf0kW
B3ufEh2mmP5cgFRVmqWcI8pdszLIj8yR88s4zvrd+OiJbVJj9NvpA341AgZRMvQPTrCjHACccoaw
4rBBNB4lwEtWu9/tyCjTzBv7Gd0QVO62Y3beKUO0H0ig1sn7JIMa3qF3n5IeYsb5tLYK9c+R1QHF
ihIco2XK682qrFi77r0aY0ZEcsG7vZucQnZwE8VX2+YXdioajeGSiMbVm9W+4SPSpPWucJZy+SvN
sf71ps2ZU8D0CL9QAY+1qaOb57kqweQxJJIemu5Zy6O51Zf8a6ISTeqRD96bzE+si6rTk/fzDtSj
HwaE24WHzJylwtkRVPKpKRzH2sOcsEmHPmWUullVeOP+MPUYDmfgcvP2BAH0iy3plr7QDEf1ZrK/
kMZ2Df+LEjeZ3oTPxzvQ+V9XKSTpUSihSjfyrvjsiGQ8bB/Kh0e3gEyYzJ3jv3Ek+TSn1Q3Qu7IJ
wuUUG6NfeRhTb571CpBBeLAFexYnG2n5PIw5/V4aDSNDmpilUZnsTQEjkX3lJcUphFTjPaeFZ1LS
orm/uOHsY9PqpVKPJ4rpiL1ts7VmbGAGe8BqcuNY+tlBPIlsVKQJaEKhMzYhmof44qmMTA70MXCY
uAyvdRcicAH3w4Hi8oD7JS2lX3XumddMSR4CTeHXIAGOTEWZ1wxUbuCHmw21iHghMrEGIUN/6Xet
Wp4Q3tj/1T8rOaPOhnBnEJwjsyyWQiHcTWhuvikrbjdZ5MnYL2HZ0GQafMD+OsGG9LXhh6pTaUnF
bGa8w3TesIg7lWc6WklZCxWiUJKZFMm3P4vUpnCd+PZnxkY6EopA+p16pX9RlKJozrGc+YZnDDi2
RhdhfNlYDm7UJ8weQzhs2zE4IrKUo6xMWd2bRynLT9+th6pVKSPBIWdPp7FIN8013A6IWyN10p9G
QUYN55/aB0abIGeyXOmvs7NIZbn+uviPcY8cyqTtPffzI6MBaUojE9A2VdGDM4onqHOg6bw7YvuE
oJj7RIEwLDxgL+nIKS/kYIICv1MaQxRlywnwh7n7aR7nGtlrG91zfW3O7VwtnpBiTsZOETfAa2d6
QygBfai9BySzJINL6vEJ9NrDI+u8zlT5HM9UJJlf1X2qA/fb5pNrqv+KwQTvWrzjZu/n28W4PdPw
eRuqws14XYoIL/b92+b+ymkHvANH+9FHhQTwBkWjSKPKZekB7CSPvwMoxtL55n2TLP48ytFS0gKa
2TeAZceWRRTXRV6+LQEgZXuBeV4crQ9KgEUilggIBwdNC03KZGMxL4bAMyQOpLNhwevduJmS9Rhc
shRHWktUy3TxDEpZ9z8smP9ilU42PcNZHEC/DqT9IYXYfRR+TJyqQrp2hxKrwF5xe+BauzUQ+Ia+
lRwpZYQfibdW2V1TANtAiBLX6a0Z0dY5OQOSgn3zzvNTEJQHls3jcX3ehqXV30dfbR/LyGtuGPT9
Hvtn00E/N7xuIXZCGwaM0hjwBSjiswYjK1nG00m4z2uI4nxdKXgRcy/1EKPDXS/cheHlJjxdoAWa
XA2jtBrFqmdqM7HFkb8zM4nrtXaKse1J2geeTtVumJZ0b0T4tLMHkfxJvZho1ixNnXCpwf//374w
DUGoJVo8rWeqVtKbX4pAtyOMNJP4U3jRZp25rFq6UdbwiUy+Gcyo+hCnQtgTpO2clmrRJ/ZKW0cy
2ANMNcDPazhc2rLzJyEkaYkflJxllxv0z2iXBxbaep+M7eyltiZ4kbzcdqEZRoaOpTLgKpyXPMB2
UXaYv1cgFdjJQzvvuKGv4/V4Kq+mQGpTZF/uV/dJdngu2dSLYwH1EfQsu/83nsnIB+IdnGwh1TLM
8IawfpFiPzMLx2B2mb87FwPevdqjksHG5tbN6M6zQ0P1x4HYMUD9FToyod/jIO2Btrpq+dgz4ic5
nqal01CuRHiJXy6hTE2Jc+oEWUanBeAAhA90aB7jPkj1ItYuaoVVmvq6q01RZtdiVtBpFbewAOKf
0xg9S4ESSS/XlXIpRr+EtrjWBE+65TRJ5NocJEu9+W1E86ERV5GiO2I7o0k+pYiAtqgPjfOo2YV5
1kjJI6VtLOdMnjW85raT7yN8JWZNwTgEQ3gC3lYrZeU/HxC0aUJNWyv4qqd6gXgf2JPaoPiYvCSp
4NHDXUGmi0LEzRPAgP3Nc90lKMJ+HPw0S+xNdLnnovGbAMpv3EQwJdiWhFnsUTb/H8t/LIS9GrIr
MT9YepzwzkxRNmH+zgUCBqlckNSRH3E7qnzeZYdNB4c1TQ5XFwtrS/FsgKVeM//R5G4mNaXcCLMp
q3SBCeB+22bnZw6hPyx58RXXFf8kvNA6VUzC/SJ2IZav0qmHNdwelPFjORH5lv/NtPQN+FBvaTMb
bEhxfwxdGRVYLWb0Nhrq3snwvHhfhwQj65RA5j3lTockDnxJkNyblv/I6eM9e2hsBtUo4LgAbLo7
iT79bP0EIHnEVLOtuJ96q3E4igNcgMCNoZ99Q5LkN1OOalmcBoM8vDLzRxrrc55hz9sbHBxzN+cx
bEUr9KXrCGXTwK+slaEgJ9qEvdH7A5M3g37ewVmVHlgEWZHsBcgyuvhgAmQJT0XBk5UeEv9uUx5h
C5GXnMSIU+bo2I/SZto3RTAIWTlGhQyObPZvpS5xw7y/2Fps7XR2arw8Eh80MSzE6sCIEzYezWHV
/sEz1M38zgN26FUm6pdShxxQywCzb0ZLUYr7F4Pz7msdekf+dTDN2CdQUgnmUwQH/FisQsC1IjOa
o20elgbQCeZ1CjbdlRomFwrLgQOWWj1y+iFTLdPBVnD6Q6qRBg+q2vn6jpvTbYMyxDqSa0aIy3nG
nX0TEAcFHfY+CeebAO6aj9DSaUo6gW2tOH+uHXtk/LvN0RUbPe5MQQgEugKcLoWVD4eyOsgqdzqk
sFCiNucBx2ytrWtV7YXMsqT43tjXWlO9UqKCtROFI3NMU1R7s2yg8+H4Hf9oSZfJ+EhWuPlyVXOP
uwSnVkp2TD9DfaGrDbfQBCchjFUrD7IvgQZJXBlXXBPHBdDYShqq/16GGs+5Evts7N/Vpaf9GJhJ
Iaxw4JBU9WPfSelVjyeNZ6Nk47A45R2OBdxw5L5SeWq1k/TiFtmxcAxfibfYuEquuqZPiK18rAgE
f87r8/dbVfNfcmJQh3b0+7zgg/mEIqn9+TaRhd3pr6bMfl6HbKefRbf1Z9g5lMR0iS8VF0hn1wNU
ce/kZqsKAH3SVHplGkiKbLkrxH2MA9yYgjrt1kjdXwIfcUAvRHqQ8SZCuW/WeUG0nocCbIxCoIJe
GGVUjCDDRWuBqDfK1zkl85HN+S83+9KW8wR9+2QXsjZ6o4Ax3/SOzueYt+7UeSSjiz+GK0jc/YG8
QF1PtXXHsUQHAwxWrjrLXEIzHGn5x8bTtfEesIliKgrOjUIlZkxbCHo9EwMAS0GEWs9gLngzFVUv
i3UFk+riBmfjx1AsViu/fBO60vHyqiLNPlq0aGjGaIJeuwF5wjIHImSw/85DG6vRJH8b7VSSL+mv
APwh5naTBu0QKjxEU64mWSotTPMo0AJYSidHakbfw8QMUxenIEHDflEjBlxitf46j6UTkVIux5U4
HiDv4nKOyn3ceb33enFbPSHjYGzudCv3Xrwnhx/JabLdgB074O3KEsxDkTgCJqBRA/XiP1qiQv9h
414AiogkYUA95tETHpP9fWlLwFHQbsQjSA+od1zk7Rb0Hmyyy5E7/bSFr7UBhCJG0kN2sclaavQp
86ocvfRqi+V/0WGS7KfVLbO88AvivYvJG2cy4wcBhYJ/3Rk0lGzhsbzc9MbxLvLTiU9+cTRtBmwd
D+oFwgBctVZAKHJM5l/e1Hol6UsttF7PGTWDnHQIQJO+c1blqBiugjKxjb7s8uZCQGVkvk5AYrlC
RVK6HxWDzaWpM9nXMgMUZzQ/ZmuCJtjG41zhl/TAtTHCVgmJMXYyMTTGcktijVkENUfauxTjT3K6
szD8niZmtiidcYAzn8EHsnAiNT2ECp3GAPHn3fdRj8BvK1jcdLiiC9XFG2ie03BKg1hN70kFlUKx
8CnxlVqmRoExKXP1k+tq1a4fbZ3BqDvbOa5CiiKyIvEd9szzdR6IjlSZ3T1sCTzQPS/8ME0JMjsB
ogCBMEn3lbDHINBcRvnCYaqbbIlbW9VeOWBOsxCLtlKNY0vWWmQyMJ1QzEucQN86wkuQieFT/p4N
v9Nuoyia5P5S6L8Y/Ow3X5bIqA8shWFz10DWJGCkgecV3rFDQoJZ7kLTWwDYWganN/G8IIKk8TrV
bDC57MdyWtX/POj/imcjbwuHGhMTtflLnwQjnBBTXmWyFUJ+6di8pvERlPVb83dmh5CCQRFZEW3x
eKozusrllgjUlwnBIevWC1RmDC74Dnu4UgH4f+qW4WQyPEm2NB90wOZGuzJM6moR9dN5ko3Rd+/n
BgkLhe7lZNg3ms5LYykGwJzLd2CqUL47Q3Wr4I6FeUQqQBDWIvaysZtb4MJCp5we90Y5UdjeoiNY
uPhJpt+2pTFK98T4wJuclF3lDcj+l9Q7kR6sfiIiY3mvLxrhRpcgcn0dVXLJ3X5uc5NTg8arip1I
T6ViFeeYjDX6d6AE8NJNrpMb6Ae2EJnjCaduTCcLo1vsaVtVMHjjvF7mspyIU2ma9Hpz2HIlOB8d
ezqdOeyRxJhfsfNzU5R1lR6N/ypNm0lzVzF36DxE5u39fdwfOQnIhpTspQ/CYbGaysKbq9ZbiNRK
Iod1MTZCn+IWp7XMy8FevLXydlkRthjSTDSKYljGEqUbMvQYRBbaJVHUzSUol/ySzxpjQUUBrvQ7
XAbB8kgF5UO6UJzaYs8jGXiQX6Lkj9Thuqs1eMtO5hwJtoxgw5QCyhqUtL4BoktmtyO38vcXn70i
sWr09syWf0GFqMW3avgpsT0Uor7j0y9Rr5jFaVchu2KJsiWG6XaDo+zQvS19jEENuXlFLZo/FxTX
dAr7rNmH/Avxm2HEbHOC78duak+YutsDtPEdI95RLZMxmisxsKD/BQUM5rLy5KUUSfXZHiKiMoSk
yl59SsnPbYqShpKJFL5ABWhZMl1ujW+ON/zMJXhK6eJeCvSVLJiiQ/vmTuFsYHBNsQ2IfafqTn7a
xYntFuz/G0eFmBY+7l9YIb/OG53RM7hgeKgcnfGi3pOuEM5In1t6PfwiDazk5w3DoluVV+qt8IRJ
dG4w2NhAopn8lNvXKDxqZ4wOfEaE5X9Inlw8Lghk0jByF7ra4kDz2yUOc18MDtdaGvY0VD6Z6XoP
wvTErXA1PenS29gJqTOn7ht+nPnMd/vX8RjPe6J26SIoPZXdctHIjBRpX2no3U5w3XBu5l8tiDW/
TZSFFCXJbkmR7kGMJ4+u621AJQ0ujCSptNjwxWU0XIMwdgDANFPLbou+0rdE4byaTxxPcfLjp1ij
dcrXhYIvlPn/S76AvMWPfZwf/g5UR0VYQqNgdIXwJ0NgIC6iJgiiWjXL4MZVTxVTG5urv0T0sB2A
QvKr32uP5ROe58ocuHtXorXYxE+J+pP36igz6aiqKXFWi4/XDtjlj2PwbJcQ5PryPifVsI49Kj0E
DhSMaq7dtt2eYueLZDAbM8fnUyypk1GxzTZJ4DHZwYSdAe15EgcX/qd2VOPYJDF2atQbTeRnHwqw
KL+CK+RrGAnc5D+ONK2ha4H4scYPj87l7KpY7N+IhYSJra73Exe2881q4glBcBVSgAVX068g5I6A
G9av4tFKPkagiDmuCBFwKFTEC4OuReA12gjGVSaThBMWYRiu5j8kI6TbGp4Ot3sVwS0L1VXKIqwU
sbOcrmPoqBhmvmsztCxekONcrcL45XpL4fAMo8oacYJoUWx04OKNsOPG1VWjeGZpRM/lbRbG5cMZ
nlnn2JafLv4ljyLH6KmVQX3QKKFItw/tcVbcdV8UH2zTJ+YwiJN6YS5ifVOPdKRkfrR7/5Kykm16
ZE+cOEcTjMfmb98TRqBEdAYcBH4j0HyiEpW13lT25tYXyjQoiYsnnMLLkeCTYpirnOO6sOKf4UTM
0EcZieDLhD0Z56ywtitAlAXZhOAm8GZ1+2I4g7KNyQl58OwLDZgI6p8KY3NPPiweTJ/fs80V1PC4
Dp2oXAF/GWmvGOdq4MIyoU6K8Y6z5AEQ2wxhUbPxFWTD1EbFq9/GvHah/jellFzbAwxKGY8mt2ar
esSYoV/0heilse0seJEehLuKQ/TREgvTodeiia46w/rZFFKad1dpdgQE8EZJDjf+H1PxuD8b8QQv
hNpx7M7rkimJwOnPEVQCVwH2ntiDXQCECrpZ46gii3heZt1pma7b7Raq3eLzrhmHYAAkcOrrIPJa
eHnlnvyYCIAuy11WFVrprh5cXbgt/0Dt2xk9QfpClWLqTE1/dM2EUIzEZ6QV+hRKNcNEa40PC0gQ
qEOunrBEYwE8egI6RIpUP5PRgbr1M/LRM+xbXajiXkKcfkglP4PvjO3Kbtdf9uC9jqU9lrqR3Zm5
cBnsDrlY2ntaeuc9nc3tHXQ83Nq/btiRBbBZi4eX3sMW2Njit6drDPKMw6JelR6PiBBjsAEpIByU
5cZQCUCNVqHrRfS1bztl1EQlIa868VRtB4BNg9T5TfE170R/4/twIOHuH8XduJDJ5UwHo1sSxgdz
9RzT3fnV9w1nAutRErjVjiQdmMJJdd5wBHT4yRv0pWZhdIJ1Ahstjfprhro20VbwEbRLuld3+Smp
RJ8IAZdg9Xcj4pvZDKKIQYrAKDmQUxaZqBpgHHFulMQ8OwRcb2T63X5NajLrRhP0aeeDOryj00xR
bS62YAullpF75tJNBYPWxdLIekKQfv7CW74pINCr4hsSqGIPX8zcodo/0Q0HoVly1TDdUQR7k8rV
+5smiNaq0OISnl48Nxn7Tu9UIld9eC8uWztE2mfd4y9mBx1NXOI79MQ0IRAlYvnzsl4d25iGbI/1
j9mc5j7z2VxvaLKVlin6ziEmpB/M4dc7dUgehNSTR/SQd1qvOHQ3nOOsngLDSdKJ+kKeBLCZ3bVF
k2ajAXTWn4IN0GY0Wt+7xUG6mTKlbGakJ99RxwAKBp22RGIguAZFpIQhs/Ycj6vEUwASlOXUpP02
G+UVoyr1KNcrTb29bfkdrMjQYmVrkUNdYz/0YcTOcNhwzDMVX50Ci3CaH/7nMRDNNUSzkgcpUTHW
E+LaOF/8/LEeDGpaAT0ZdQM3IVPT9aKpoJG+svYkrGtAPkgUVX0B3HLWi6DJCvd11PFMIaJ+zVZ/
AbtJ8sJe5n72VchA2326fe7ozmE8Zpyq4dD1llrkF5Mv8Ak6lrJXc2CHgNwVws3Uqrv7tGz1kad1
yELMjBlzh8fJv/UXZCUIGTQF3vnZkGjai4y+FL6aibmK7tpHwl2QggqMrXf2uMX0BDgYGXBclHAi
QZ4XFOaNy3aKL9IApmP3O/2I5Ednl8njM7bUZN0adJ+zPG7+qcEjgOqcwDiClm/mjP8hB/Vit3TR
rvORFcwgzfqi8dJcq2AT567i5ZXUxjBlmPOe875Q+mCUUfvsrhsUm5WoqCSKBLqncr6P1/W5u4oV
22JuugNA5YvVmOjBorqS8qe6kqL2NUS7KcroU1A7zPYu4DyaVgALzE5uuo+0sG+AWh7n51Np/VCF
OEpLJHsLFeLAvuTtCsOEdQ0UGYOD6pwFHyoa5ibYeAyfot4BdhxpgwxHiz7SG1Zg3QByq/gMkCEh
PO9mIoMiL8+B+yiHa+PIfiasu2cIpkxjwxD7rEnDc+jebbflNT3sCDRcZb4q0zEaTPDHs5rzq+gC
HaKC3bNb9svIY6OMsGWJOhZ/2szvZa15fr+GuZcINHQgiYKQPKxmrJd1hhBAFaC2zhy3CgiZBfyg
dKjO0+WvKXvxq/7trJ0KnfknowIrqAJjCzuxtMtbbUrj7gBht+Eft6Sdcg688JQqdQjwVw/7m3JI
3TxOh4q3lTY3RaKG53Kg1XcQ6s+YbxGZY+q1DdxI6fc+K/4oYH0h8aFdfKJFWtbnynguJYg/mW3X
5zu90Sxtx4+pGKZROkG+pTpy+a3kuBIWO+xmmDGO9Ap6/mC14I+0oyh9Rsp0hcohSyEuPUqewWD9
Lr+mCDxO5JE7GETB1/sd10TiDvRfXhHr2TRDhlJOxnl8v3F4eYUYZgvItq1cqE2kUiAhsfyEXp8V
Z8euho18t1HY9ppltXSiavTyK4ln4l+RbdCTZkLzAjLH3gW81+K5OcAoAjwFK7G08+1N1eddVbtd
zCiL1a0LpsYbUODZ1LqQjwBsX40KwY/AQNGTuKRCQL9VddN4MDBLiuyAOSnA39iZifFVU0DATuuK
Ou28yca7+afq/HguLj/RjtFwQyBNmSv/B8jy2epgGgWwLbu7WaE1vKxjC5NcQ92rNGZETcjXErvi
AX/4eDoqB1tQGuJ99WK1dceiW3iFTBDZap5qythSR4jsTLFom5AOAu4FtbMTM4mGQx0Hd5DkTnDL
O8fKpF3DjBOX+xc/ls1hOcRP+xXGIXgHwfRpIsnRUUpPPRaydMOtiIAuo+8TwfvRF30y7gy0KquY
aA4N0q59/lcIBpNZ9LJPQWnCav5LmmziFkQXBU9G6mZ0+WBT/tyLi11SOl3Oo2l/g2WHKVMhQX9V
FDdSW4E+JiEAy3UTwEbKqb1ukRAn4y+DvhqqWeOYHC2EuyHx5Kmv/ZdRKLx1aePEu5rbY/QARuWB
H8osxQC7geRWGL/GlRnzuI2zKrEHvRn5b5KzMpG6d/L8sT8StzG7Sh+wg1Oj03I4Wu4aKWohfg2W
fzTJivZjBSowrvrHsxMSR58alInyOmgwhaEF/YBqFL8OzZTYRMEnN8yNSUiNfL40ukWwI/X6wP3w
YJ0OrRUF6tDXdKfDC3DIzJGIYAsP1IvPrMPIEA9m24IRPER0ePAKTChUiaOtm3n8YuUH3Mr1hDfv
pH4KmkKa3lUYsT9QrWzl92htvx/buDD2uK8ky707UxQQtlx+Hr5f2/ndSDNvxUKdHCyOgNenDXd/
sAIETFAe1OpxBOrRBo2AlmUG8imH/5amA/e4VIM8DgXJ+god8yb3skPoHAsj2cJIHJ/ZoWizo9ZE
+BM84IJbVchRP463RSx6qbvWlPJlCEN5B87uOSVL8ZXTaejy+JP+vndoDsC2NGIUaCbSF7tA6WC/
wRHIdTADBKtuF5CPWkYZUsWHH36d1Y9gzHJmL+6ijJP/sryPSiEfEqFKHJYN3U+3XW2sIy2Pz1Pf
Z9d5UH/6kLtE41k/TpZJ2r4Yf3Q70Ncwn6lhNmHJ2YG6WvIiQJqKeql5Vw1/KerbJWftKY05XGVA
jWLKSZzQIszAuU0bhkRrUT30Moc7IRrsIiHfNpFXYwWhmWN8UioOOuAu8o8QcBaXRRb3AuqGTIK6
YxQKs66IsfBmBfezYx0PczM/0NyKbNGWISQTmtRj45P7oXHV1FN8IBOGw/IhxMJSJGsK7F7kJVDu
Wq60Hjvj2linMbTj/CGTaUYa7zkH6Di+didlR1LwYGACDc1n8yKj+FJkcimdup3uNBZ+3pH2Z+cW
fXKBMYAbueoTbSn0uXZiSUT2RxfYsNMzPHrj7mteEbMWx6i/lKRLrTpc17/5ZC62DbNxG+jTTL4r
j/hZve7BZJFgAyPIUN3OJpl5qMwF+2XYH8mRbxXRD8v+2v5yv8dnH8fVYPPaK4PanyIzsi2mWbc5
Qpg93DCswZIBBSzcZcLAn6V4FtrbRfQgjXE6ey9GqEeNJO1Uos9jF/4lZaQIk6TJpJ2hRlfKBcUI
z5ZDOsMsKLd2OT8v8jEpgkLJy4I1L+atTyARHlq7SJiwqqqJsAdyBK2WrYc8/Gby+FnOecQkpSUU
BSAZw5rNeDo2f1Rd7/g70gvooAwJzd9vrHhFwtp30e87FUX56eZ6jFKP2cT+ERKAm8r+4qwVHvLi
k1wpgHV/TGH2kVzdD9cGlVDdfYIG/+35bmnF+VYPkyVLn3cChYWRo+CxR8qgPCHzLI9Z0CXj5Emh
itnUdxAQ3B4e1Q7uG0iq0X03WTiMXxnG0vPmppnCG6FRGjDcx53rpPkE2mnRUAv1jO1Ar7d1Ykwq
pbOoEQv6En1FYw7JQxroBy81DJ69EevLTOZJGOuXe/tGpjpMnZlZ9GybDgCOFjkQKQ8CxW9GvGOp
wsWjdBpgxDHaoArOe7RgArGliDwlIZXpj+0/1d5buE43y8kchOSf2hP8y8wMy3UOjMQgInS6FO+w
U+nP7MaHo1YDItnaFDzkVDVeGLU/3ttV5Mc7Wez12yjsm/HiZP0GWPVnSuf5r0OG1gWt/4YtozNs
+Z9AcQG7/Lv45tk2nmfiaKXafU/ZfS1rMJdIyIahkt3YcAcfx5s9jv2sJFUCcpfCmFyOTuIrdPRb
qaJYpDYbwk0edRIv284n7AM2575Vgh7ii+Cuia6as8zHd691TD2wb2pugP9muTPx1U0H8fjyECr0
OBwisvAxp3hlAONjIPPPa357CwTHkKiV020LH+lscwQGNrmXLB4hAnhOan8QdrhKLiLBfqTzQhrN
B5NFTm7iJdZ3ebIXvQre2BgETeJcnQSDEAdnMgKxD9I9N/bZ2KioSCAcTqs1wUCOcVD57nwnubxN
S8LRNP1OxqjSiLWhF/S0sYK9E9bsn39vao+BiRP1HYND8TXZo4t7uQqALusyETr+W+kphXzbpZrZ
vxj27G+XMTZezJbizspl14Q7pRmgmL1F9Tizf9H52hvKcStn82zyf0F1k0ipiJyFKfaC2ACDWUUw
LInNFL4K4bKf+UzS1+R3kBUKamSQe0IPjjuKNGho5ExUBGsaraB+leni2gcbjNlw/eGF6wjfilgj
AGua+4EFX0yxXmIg2UFnX26RRym3S2oAnlugNv1ausfnVAJb+HCVVlMvp01sKRk91dUGa5dfsIZk
FedB5pDfymet42/SS87xuQv+iqmr3eG8pwV7dKgEbs4xskAe3ttTfJKt7rmQYOdwjAtYoET4qQX8
dMv9ILXGsmAiwbkiWn/tqwkCK2TM9XZwLto055dQ0nf1MJ8/L3E2c6+nVlm9M/wR2FHEg3p2xPGR
3aIM6GR9cr2vVmIr541N5gq+83ktsd7wpm5opoWYKKbXNi4av7D6jBAbFWp1EbkmxeWLb1BCf6BU
scAh4Srsf8ZgveRm1uQJgnCKLY2LHEltuDsBzfZRrLjyjykl6Mjh/dk04kPNt7BUEuNQ8o/VTpiB
NoaLC8lzWVKHdFDW0mB0XVMqKBNnYwRzHZwEIV1goOLq7RLEVeTyQq0AEQa1gOpNlxdcoV8qw5z5
4Pk0J6Vb5pcP95XefvBKqs4cLNBF7/Tg2V3vfWMLwAd8C8UhrxFssDN5t1iCXqh6EJlHuHfQjU6p
tfn7V9TIspFaSvYh3o+vSBsijI/SU8gNk5NjGVUq7Vt0WfK4eTBRFYSr9Soibzg8+v6xhmWy2gyE
CqD1gTIADtVTbR+r1eq+EO8L4aiIw3/HpWdkLSL4lZhqFpjajVOv+xAdLWmKZoo3YEM1E3Z0gsfd
b0QDXIi+IVVnnP9M91wXdL/zTfw3p2Opu8R/Q34arnDJJSQQhmKuHlSB8iulAKzhE7uEmo46hQ/I
iCcSTmoj5BH4oF7GeL+CBuXHlA0FjXdhgB2bCPVsQHbPore8OJeR3JlWX4UDpAWeaEuNwHhSLKiu
itAWNLOD0C3dDMs8HCxyuQOcwPlZ40Vm4EWFWojaIQ6s0Dg0GFjBgGuk7AMdMzQTIFdA9zu6Fxoz
GFtC+SLFXJMBkMMfwumuF/yxpohpMJk6nYuCUtluwLK96K300zlMJDxW71GAf0kUPxani+M0njf7
v3Brja8O8XAyDMaeki0wHV+qXzNdqjOKsNkdGfsYVs/Ui/Ci7v4NhB+c30s/5Jnz/yH8mZ3MbTFW
flGCY3FkQKqhQJHNEiL51Xzec0z2KQbBxMmMV5jB5G36AtffF3pywRgS5Az4Mr7wLxQn0dAP9lMt
IyBLhVpOeAB7QSVad1WootA++lKc/FiiGLbI1xqGp+JZk6+u7z/WkYmph1W6GDD7Zvn6XxZGC/Wh
LxuYLh7BkMFZxaFboKgm8W1mSZVSsMohzU1FU/kpQLV5yDBX7CvgsO/hYZ1JcLDLPp7JkwG618+T
M/crb7Ojb3k/y14vH4A83brIuVaxul34JWskqrGL/Cs+Teq3XnGNC6PxMIwoHvcE7azyhvpCngi5
Z1H4UMW/Q774JViuhIsMg8G4ss3A9hNknR2rI28PzMU16iOCeJamm1kGyaCPenIrK2OP1WbUqxkj
kAjM8sd/LL585xfACYldTNpdAV0jrnGFSdOjO4yF4kCQDNM4nlZmSOmzPWYfoV6tSxIhFf8ZzbO8
U1efpgwR/S5E3dh6XXzST+5PkOqwCoAEmegNPYYKZzvdYl0BOPS7eLuaeutO68M5hc/79egu2iUf
neXToSi9LAfSdPWC9N9UaL88tjGxPApcJ7S+jnM45X1gVJPhGrkKKvL3t3GjAtG0JfFRwShzaF8M
RINgl5wD1dqnvIozKTixIOtyXcX3y0LCOmlXZ55y1jboXbe8+dFKAtLtbrMyzVSdRBggkWh9USgi
g2FV+hkyyG8YIQZAnxhB2IpluVNVRs59Xy/fp3JFk23v6nE4YdXvRd8wi9xjH1AbW4ISEOehNluY
hXbupbpfvFExi5aCVPvyY2eXx/WOQGNZhrOFs61BhF7U+kaT5lWQ/O+oWh2cD+wbVvLlpQ1hKfZQ
ybV66kDRWmei98X2E5/TNm5+ebFBZ2LvihmwyrhfvlArFejE2XyU9kf3uVUHxVK6+rFGdA14zVHr
qSBpE5sxU4mQGnr8z184zo1lX/IXtb9mSl6gCQNYGPRwgPAK9O55vUcvyo4PEaZtIXedD4CBH1qE
ncUKwFwI3imZWlsfmS6obQnYwo/Fh+vSIh744RidrZybJBOP52Ok361enI7do1RVpNfWeboAdjtc
6Fzf2C5q8ZiLR7eK0E3dxCzH09vNiFIGKc8RFx6kVFjnjlO23LzTTZiP8szBfRQfjaOe4afVUj3e
mJJcsuoDXcNUNNDq6m/Y3gtH9/XL3iT0W1ccpQtqPVUJghEHAwI3Aqn1SL8/wM01Z0TAihCYq4MY
36JZgeipdT6Bno0EP0PZM78svwRI5xjtTpl1OHZ9qczY0JKe4zMTRLFQO6q5l/M0mHZhu/zEPofQ
m029bMB+kkuZsE6ilNDvsrWlVJBskO/vM2KuPM0GVNZNuCm++xKFD9I/jtVw5WicA08UZwtXxS0i
QqE+cAbSCPoMMkIhmtC8nWe3mb7teS1xhkuuhh99W6bhXT94d9+oiL26upQcFIxQJv15LYPWDsX4
S1WdII7sLv68q6nFX5GMfYO22u8nCmJxvPEf2Nw4+VEWPneU+8wNJAJUnFsXUQXx11sA36MN3wE3
20Grp2XnxPSAjUKomGGdSBqZPMKRnPvUrubYEOTMHuCr0MSNVnr8YHlOGbno562p0B4Rmn0f5zw+
4hJp9DaGxCo2zbAw38FyIYJk4OaTSPfdJJ9SqyJU87fdoeC3MfQlMstwL93qtu5w9dpgXP0y98Q3
k2bbTl4+4Na9Dq68ZUN1YgsnCrwflDn2E0/k5KgrziTQU3VdyZxIiBPI08gIq0bFrZpnVrQPCM9K
xDtsXAZ57f+6e6e/s29QbLXEkKLhasdAtrwklkKcMi53eiQK6bsdPqQtzGtXjxXR4mOjbmLn6IwK
MByRsWXnlwEol3IcBYEzOixssFKTVTHP/vU+1M8e//vRbHoc940DyWX/BSGg2KVbHsPencq9uYXW
C0GcRQBKiEux7uNWfnXvflI376kGScltmnJH4uLOt0Z9lK3NVOyrngHM5ccJN2AHIgimK6ZDHmXU
rm7kRHLvM37g9ewtKg7K2HOv5rXq+sUx+7CfRyHLorqa8GeK2GGQUPa8KG6zuRNE9G6dym3BV7/b
Hi6RVb0S24AKQF1IjHP4EZhAUEJwwky4t+eaZl6N3Kb0VrzAakpAbJKurc+vpcVFJqKXM+12kRqR
hCZPTRPRxRpzTPwayfaIoW2gbXp3NUTVMucc2DH/SNfRId3+ya/Y9y9Vrli0y67Il5ocn77OZH99
LPrJrYAi+73HCoGz/gTgk8AwQzp+Gr45iqYhlHq0NzVeM4euYlLXib65DfpYiQEg+V+euliqXA//
M+2P/q9tOfDK0pIBL//Hs/u5kFA0NKprZz/nCHLcQK1C0GG6jLukQKIt9SL+4z3i42QfYLgCUNbQ
WVAeZLdrklwSES9HZnucrkxTNU6zZXlN0O/hQQMAaZxoNk4sFr5y9wqM5UCAwr5tS1qfy0p3YI48
SORnIGT49DvhD//cqkAWlhnk3KwgYd3sbQkscFFgs19Yy6BXSvC/yEY4XunO2IVdQgc8kzQsPNfr
Q/oDqqyJeDaTjF/X370Xtvs6bfl6P3Es3YXIT7mF8xdlZEAq/fRU4984nkGFQcYX/jA4J2+bYfP0
DTIBLaIDwh7ruf8Ety6xKF6j2Cqw6NJvrVKF/o5AXvQ19ddNCL5WPFE21VNbXpUKtVHwIVicrmUP
bfBhDYW4xf3hj16NcAqu1aXiQNQIVIwhzkGUWjCY7BhTQUsFy6IaN+wRL0EprIwK4Y6EZ3+s/Cmk
u0vQuLeKqgdl8v5hRHaaQyeY/QuMeR90i+604+YGbSUHrA2Y4Zlf3OT+WTvXoZAT1s3t+HlNf6TV
Ql59ZjCWWqGSPY6Cxh38mnlYQZBwFKfOoE99gG7tXUwI7Yrma5cnf9mxNMheCsmk7gpAzW4qPZ4B
jIk5iFM84/ZnedOOMldLezW6uxyKJ3FZBHPw54pBsBwuDXQMf7622o3bzKEF8TE9qN1wA+bm2d2A
SsX+/uqpdpE2P0y5NK66HVjgy3rh89AqpEz1OVdc8+MKr6yhjIjpGAIcIH4DrDekXuTGYFghvLsE
qrifGPnxjLaZGnTCIz7yAYqZjye+/t7r+fbh4XuixFnW3k52h+x3H1KNopY7PGlXqeP70QOzCmAL
xmo1dUDYrwJ66oOfYhgkIB7xTPFTOnO+cFniySepCqx/TODGZrAyhaR11XXh6/V9MbwXJapgn6M1
0V2XmQURjSqHCawhloMsLLy8yRXOwmi4BnCDW1gvIORPD+T9tECMmmjIz44TFajDNvF653U5KcAw
hAWFqoFaePtizUMSnNlRLOkBSI6BliHdUiV8f2xsv44QjYLfoWKP1cNoM2rTUOPPv/n95BnEJ1aG
C8T9DrNnLhDj1tQxCUBzuznTDh4IDg9SBwLipmI/NZITL89IJb/76ZGti76Q0CFZxsGIhaERVhmQ
+ynvY8xXwk6pAsFBF3NfodTz06RgylAMseaVC/dnB6fpezkONJOxfs2A6jLyaMLacl3P7IaQJLMJ
QDkIhzVCvjEJHJjOJgCz3SaeP5/yvvn2kLzqrBIRKh9I4OVz6sZh9C5QijaChAJcX409EnDjuiV5
D4raRqMFy4Sqp5S6iUC+vJKxdusvNYsT+NMgcQXPHyvM2osfYSKPP5dOXbH7YZ6Cq+IJ+w0/HtKA
HRNJMnn0I4goV+HlLafLC8BOXjxEtcC/WDHbRQcGlaT4ukFQOT/Yl7DdtFydS8R09dPPKWHGO/cB
hVmJc7ryLY3/jrPa/3FSUED/kIsdHQi+kvQD283GkXflm/oybEvqg57XETk8SeKjFxAiNNn3C07J
FjLD4GJwq/YOJe/Fttk4/e8IEROHWk5MiHnyJmzq993Y1nEuVjq/G9uKlxO2HcRISUz/I9aevRvi
+HYYA9rbzYCX74v9I4jbQpqzc7t7LZSN773PDLG6SfhGFUaPrGL/HQEe5J8LUQFYVtoI1NadTHHh
A3wFMSGgdpEme64Pg3N+CGWaFUx9Rd6AwJc37Km/VaFscQOk3vFuyUgiNJr9LLPqDg+27H89eenT
SWslAwnyB5SOc2AU3D76oLUh4VTbaPtQ0fZU4OX/skDjpQnacdOyBCjwyZYlJ77bYEFFlCT7blql
HkYY4F4S4fp1odoAGBwbSBKlTCCIv/kl/2oFi3ZcL74ks1X7FYa3J0EOr+YMjcFXdBjnQxrdd/Qa
dIzqgYEfxxWXMTITDe1UYb9IV+9u5fH7WhFWwRKQfsCzRmDIgNxOhBQLhNsrGc1ncz/XteAjdcmm
/Gx53PkvCgUZTlOmTddGKy3N/R+TdBofV8mfdCHSZfIX86gGtnVeWpNdsB8HaU0BmMhHylHhouFY
EyU2yv+BldSeLkqnG0rxwN/ptoTD2QXVx0UmE0ZkXDbPjnU9LGYETgBKZ1OV0ktrdTzZvPKt4zdu
Q+lx81N3gmwpPwWPx7LyIkfc1fbJYHl7oD9fmFn09u7/o5HXJW0mY2ncF+HWcWKRuefqYX8ZfTv7
oLWVadwq46EDfJxQkmIhQn6YVzUTxUWqdspvz4fa4EE4zVrlbFEzEcOq92zshBBBi5sb4ikliwtL
/ILqaKY1UeDik9Y8l+e/f2lu385sEzfI+jEmUZa7WcfGN6Lzy9ujItgG/pbdl1a2tSfRrRqad+ka
KRcTQbQy9P5YGI11xxVQ+xuxHRMISk8A7pA70sepi234ltpyBALDIuU5wkGdhM26xNbjC0Y4MBnK
+dVjvGXcFr7508fdPzBPpqmmSbO5wIIHbW9TZwIrUm/31fqYb7DsXUhfwsTk+lz8u2R9Apz+mwII
YEunTd0KG5N6PlrFIcl3YS9oroWFpf2vBeQZxVDbZwno2kAAZTnsCTU0GQ8Bp9BTgvjV3mKnvEVL
VDi0+NLB0IR6LFdEPXfh+/c7bRm1BeWwzowQkJ9Kvy4C6GJtMMUxzWLA2uwm4G2R2bmv3UqNO3ne
nEjZNdclZQGN/b3arWwjUKbLJtVKPRE6KXfxbynrQ3BAPHmQEWgYhLnxAm5lYxOXMFdhcB7kajxs
5EKV436Bw2/UWPENZPFmP256CR6LZw/1IquweWsOlX5LhL5mlWbu/x5Z/Bb4Xwjuw+3DpLrFJyCo
K3f3atWf3O8HOVrQE19Z4xzg1KTNcTJx1VyqrD3tjB/+tjjzLTxE5akoK86x+eVXGVSdqsO/m3CE
UYDPynXDW6MtNq93cZj2loPUwg1vGZr57aMkteju8NvtuaPy8e8NeZo/LQoywg+lUUBHqCpgHie+
PpXOby61qsojO64r/sDFEY1Gi/tczrHMTCJQ9p0Rix4QErUyhnCulMbBr4CqwfEdcx1GC/n4dXjP
fBoHG6GCEHj402/IEWS/OMdMWBKGXxN0BfwK4JFWrVWjp0Wtaa5IXCtmCCuQNm2hBF4mj+G5Da2f
9rq8hlYr4EYgYz3oKOOOrVC+SlJNmGuG0y1pQ6Yk6YFQTZrkOinqCbNsys3qiJEOvyTkwYNsjL+S
BT8xrkHGgWiBacW2caba9fsHvi3stM+NHVRXchuyuadku7iSPGYRmnYymQ0uJTJOez9/fRPOBpln
ljAGw/nlo/G051QqZgt+Vx9XAI1gujQE3saxuanNJrCwDny6dQlJRRSAEp0589zkCB/C9s8YtZb6
oEm6lV28JheUwNM7xtJPVZl8J9yaVOQy/DuxGhDq4HTiWGXz/2x9dLDAiWBFlzlL7J6ki8mq2fRO
JOjrXAf2cydTKJ8Q7C5H8iUSAZNOIm964DWxeWZtrdDnObusAsILiskScr1sOgXcGysfC4Qwv4ZY
wFx1nVOh2z4+d0XY+St+udnmUH2HsK31yE+rZsRipEFYQqIU2fTEj86s4RyUiS4crCqKbDt2XWx/
Be0EE+bsuaXWSmGt7JHHi87qfU2Bdbc3JxIC1NtzN9Y7rrUx8+PKjAr/MaezvXJo/tVAZGTUTZIc
QZffviVyVTamjmli3SLYS6xla9vs5pD1YNe0PB0jRhaTA9zCVRuBifZtPcqOy7B7m1KHrR+mOIyb
Q5KQVbB5o5OHIxYpuI5ZSNP29ELSfDLS7OXnwBecamg7XJjBL/h+YgRUN5xc8C41S/0O+y7UqwvB
lQlzgZZ6DChwb6csnTxQIl8mrZ6cHloRMr9fUIthVqIs34+pA8QTF/XaM/xD3r5rXYzvMon2kOpv
taBmBZJUC65tzEmgLHwsXvdoaGx0NWr3tAWWZVz6aNxxANA0WshJLEJhGcTrq/HbkkfLvpGTIAS2
qNaC6QVZy6sFMPS0ptPBHUr7reQVzZZTNUj0hgeFOWF/k9mj3STkPH8Jx7KPZKvJwxs9kJQXh19D
z/22534PR5D6DyAH8mz3Ea091IQnby3V2YPJgU0FWAFUUU0Tr3z3i2x82wE+nlopRDj4HTF5xxF+
rusx8jn/7Yvbe6gQOpfwnyK+ZF6kKsHAKs/ULwGgUkaI6qTM6II+CQotzGZuedGKjTRLb+fYVQij
h0XFnQEWeAsbRV5Y0VFA9zstlqZkE7e9jEzoh6iffTJSbKExxzMG+HsprS+0w/rMS2h0R2HVxrqy
3eVdqNn8pYanNQ9xAk9MKOtJOhR4jYtwMhwIWkgL/8rOVH5zTB7TCOcG8Q5+V4+62gtrMu8q2tey
ZBZpEhwi24paF9uOBlq4lK8ulcYGJVZFuTWHlMMC48FaUoxNz7C8dhExPf0Txp92126Vt+8lwvRs
hoLlpRDT5mX8/l2bjl648RNF5MSLZzhFD5XAu07npxN4zXB+IqHkXJBsIpgNPFsS703thlYVZzFu
v6R8k6lmjS9HmSaQex/JWmvHeSMf6vHZyzQagL/iv3Nb5RRB8Cg42MPR2sLJk+Jk5wi/WUBfH+XE
s6XEz2Dwv3t/I2sPHznNQwq2ms3axh2xKBRYe++mXzO4ZSTsMj+cw+EehSEKALns77lvLSh/UAuW
MP5HwT4OndrbEpL4sabD3pHOG2V3MHK3OZ2jdPExdQzrkSHPRHcawiThFrgpuSucR5Atzcf1vN8T
1l3eAA8hZ+QM+NjE3frEk2rHKUmdMwzswXUwVAfLi1pWESvsG98biXYszDedXetlNGZ8kMjZG4iC
GD6ojK+QE6P/0vrZmo1LVsOmK2EwLRJa7yZ8Vw5TFh+acdzcxwX8E22+k6pU6NnpPQnq1yCnje2e
lzUiko3YcnW4PtkDgFwmazg5Dbm3dEwUaaN3wtVBkDnnutiMIHX/yEKJex0C7TuDGZv9tWm+TQTD
eqVd2x+/w/hlBcx/kpoVl53jN1YHVMAZ6SdadgkPbYna3UN6A8RBX8rLB7g7QMaaj2EWZvJSxaqS
db7b7XmtcH/hiDO4hgeaYIHRzoywVpna1ZJk0j8dukNm06rSOTl7Ak5ClrXwUrwPM9JZIq5Q4PX1
1njOj0Nc2Wjb+OfgJX8hNVLA4HkufZHf+48XBLJst7ipFuVjySrMHHLMJvozAGy1o3fuLrY0YDoh
FXo2gi3JZp/noguCTYlE9BoRU6jAa5rUvKJEC/kgz0xu1gRUPNdo/8UTVMsYr9lCcA95cV0esygk
EENdS2TVSQQmRjeLd75LAeh8GyZEqUgrurhO1Y/o02vqs3a1u0wH5Uq6O6uXg4E9NRqsp7aHw6j+
CB/6SKho36p4Q8V9U/BQtBTC/9gz8hXyJQg9rERL3qN6Cb7YA5XvlSzEUpBwBpc0kSwz7aidfjqD
RurXOga9DY4ohWtvXVGkDkUk3Jj+PexdcZs3vR4YrOK7vepfuFGLzUxnRhK/X7QjrLXAAGsykjUi
B19hbbg4Rz1NNTCTIagtUZRf88yf5bOuozhyshQLzb7MdYxFaaFPVcFsQAw6GlriNFK/CuNHpCTP
/QAqoCMVZ5g+NEu4Rl4q6hkEupmnskgYAUKDujXOTGG9QThk1uRJXoAYKqkH1qmT5Vme0EFCZS31
nFxpfsTcYINInYvqOV3UnHCJWXz+G/VR4EEf3L1JlyOAf3hkkFuUmNhJXxo+zoaoFLPOHJAgy0L7
gamcm4o2SS7AEOxT4JxcGns2htBWDKELwaY05Sl8csSg4nCt8j6wAd8fTd3hVGR0DGh1oHQjydAZ
nMUY0SMoYyXIRziFWMyC6gpRhmqPPl8LUpaDPw4mSzJ+QGuEXwzXKO7x0ivaNpFdOtlAJsoyF/ds
35KswY/O3fDMels7yZOfxWWynk02UYNtf3ZZyuqOFe0lWbXNID7ThBsp69zDWzpNAM/t1q5FT7OI
4PVtgKfPJ+EhrWVwrkh52G/W4YCaCNZa/ajEZdZRTC1d3+kndObbdGkKtDUbTkATp4XxPtGWxDw9
mnYzpUeI+IA29fr6/5MgrRpMnsIW5BcChQTdFPIRuSdg8rrG/IA1RMl26r+z0CC6yfsVFH0vISej
ENZxdU/Jgx1j0OqhyFDD+8B7pkW1PGzOyUbYNY7JCJhZ7pZT37FdundWBiA6uCWG3nh0x1LhEE8n
QZZt3a/I4DQbVACiq3rEQcLeT1OPxekxsFke8vW701GVlV4aVVXNakK2TPAhiJRiKMkmb/vIo9JW
eEwweHVTch/RPlbesFVNxkEFz9ihLJamIsS6o6KGNV7R9U8MjEpJ9nZ/XyKUxfhQrpLEtsCqqdIH
MEbv1RnvehPJYrYa9HRAhIW9LqcAATMqP4xqOzNaR+mrPvwkSrfp4OiyhLclImtZuK47mGi8nxIr
/Vix7rJQaZLCZUh0C71IohfD2ClcmHItmKR36ndJcxQJWhga15UaM+NiEXtvXEAXZSLk6HTocWsa
JuYSWVqrJlRzZQMQ3+spUg4Sskxu4DHWeZ0MangdUCr6vMn12EclmcsI4ZNpqg0m4GS5SN4RMcFb
CauOTh81Z/lJ4ez8NizQXr6ERH4xaHKHPOJFIjX1kSUYx6sfCgfJjnPcPuZ3lq0X+YozXe8SX27+
62LZ5/TZOUpWXW01ufGF1WeERKu0r5BJ2ja8z1QXqFZNur/qdAFgWYyZej7K2iJAE5a6wYwkwTuK
KF8OVWR7PfLB7rzLpnCG3VpoQgmhk5xKZjQI9w8XchahywfvxN1Xyo/etW4oiCJlaCuFFv3cOJ82
jpyT/9lGc5XFgXoRiJqKR5R7df3pG/ea4iieuiTVOUsAtixKJKbF95DQPMNVZEInPAUZlNVHFxgp
TNkIG+1VLGyZPI1VoDa1lcBg2svdfMCzVUC+j7sePQNwY18EdXBa4eAnOnk3E+qcD9UvIA6PYgtv
PQ7nAT7mKfHCdUWruBOb3S/+RcKyy5zO8IE9PAReBvzzih807k8vDfHYgO3/atpqNEiDTTmkXaEo
m6+bTwdeRHIWGnGd02mvjuQHCTfHOhURaNuYTmtwkNJ/shGWszSnO37I1cTI3dBzBsp03nynUJmN
4qvbvAfARuPwF6JF6wI+yE/DTrMu6uZ8wKJnjHOYUMNMFdDaclHHM0lCcA2avRAAL7BKKL0KqosR
KMwHQuZrLomWRQOQ1wQTSDPbjRLQgN+6v8wcb9wz0wNnysLCpRrWCKzeotMpLKkZnb3lXa0EoOnr
X31SxzYzS5d5a+WRkbm9r4zPMuOvYez4m+TvsUvFTPZgC7qXhrmPtEOzxxXAGYTG8UZBuM87C9fG
Ht6Hwl7SXbLgwmNLCg4u59TO6L/I4pAF98WKdrkT13j3hEdXAXgiW21+8f+DwHu06aDPM4krEgaD
CfDxNStMotfBctuMkUDV2JHGSkOIpZTQwFnolB50sV6/SgNotB8+P0dD9DNRkrJ8CdEVKewqeuyb
el+d9Kvyu9mltWaNsNOXAKL1ooI0Pbv+SdyDni/jQ3lhCIWDDmsxGN+NTUaEbaTMAB8ryE0Z9riu
NK8jJDqisnibcy/BT6IAl8uuOfVNgKyo47BNL1s/ydJG90kcwZtl1Fd+6peIqrSNFHFCqKwUzu8p
aTIhPl/xFt6A9zO5o0KHNbv5ZOuS98uGV1OCpUQFuq27pwYgt8vi46hAaNnHB6UmCVdXMsEEIxVA
c/M6/Pn+blVp/0QdcujmTXLgBlObGA/Q6lnCtsWiIMN6052LFuji/EwRDSNT96OzujHfIOLRWMsT
+29s2a0YZ85NHusuDAS2rWF9HZw3+J17MXDNV9qv3fe8tD6CiwIk/VdpUGN0rEuI/eol3VBAqSvH
hzz+2l1t9/xv89S1Ntvkp7iupMkfFZQr6kbqCTIfa+f8OPAhVa0vCuwaPgvFKbNN1WQDRDhZqa8K
YjiYD1qU4184lJRdixT3Cqa8Qour2X9zW8CQdRDj0o2k0V2pxd4VYb9YP9e8W42QCJ/s4o16SOFl
npeZsLn9LzxdnWDETuOo5ZINIQ9A8q5ubSRMVpYQZoPzrwiGDwczgLlTjJIJ9WXMh1MUJ4VD2dHC
WYl/6QnXyUkl/oE0+OzIvnS2xVOBICiDga3aY8q2Zpi1j9IUOehMOEynJbH1V8HdHPxVbO/YBDyP
398VGTE9HMcYYZMbaGUnQkDJXUU4E8s6DN0SSUiHlXsB9etR0ncQIpyo+tDCNu4+i+vwqvzT7E0f
nSMPZX0hOuq76z9vdM6YgomLmOcQ3jTTowK9O6ggI+e5Sodvw8vBFJYs5HatRpWhwbfPlG88aQAu
dHwFxm1G5uKuYNcrpGXp42vqaPuvQfWUepnTuweIYVxzoId4ceVP/3OLnr7SFcXjEGL8hZnEXi87
T+f950XBDaDPc5uT4viO04DK1nf0uPlsWBDl6qzPu/PhNxPlRE0KPDznXxWF4grtyaMUjJyqfIEk
yPoQtduyLn7H8QKx/AnrF7LPsPp8hsvPIf4masZd9kWYAvCK/VKdwDPYgerRM2HB2mOLEVj0QyhD
pL/8uvvF91jy3gEfB+CSFdpOxb3KVzmCKdxHU+mstuUhfU1t8gWKhWOC4vXmxvW0axuyRUUg67Sl
Uxvgomx62KQV4ipSAhfChxKKnQDlfDfCWUFS5gLIG0npnlBCRyaPzpLcrzR7c0WrQ4kyRRs0ZH2p
0sELWu8P+0G2Wuy5MmOU/+qxebm06YzGC1dgDfng9pgZKnffM8qz578WaYKUhOXD4pH8R5pUxV8h
1zQVslZYBVZVKJtn74qbBHBVzfAHRUq2JQWh0pSvGQ7trkj4+iJpi3+Rw18/cNpvVjFSJ69LYir0
+p4uV+8KVFUWHS/LjG4zC9FiZhdVO8IEHZvyRoYdmNZtd38Wr3qRqg7dzOgq2bkQB4ip3rTm8gAt
hxnTTZtSCCPH0SLgY3Xovih4iauaDYC0xRKQ5ATFP33Awmp0Ej/EvUrieM4XMlqJ8sYIqdpV9s1Z
+U0oBkrk/ki2WF/EVjKmIf7uskGnyIu2l6PZyDlK+l7HSt2rxunRR4KxBlWvahBFemhi+KEnyKKX
/ulRAZs/Rl2Q/xiPBODBeWnREULibboj98cpA4DuXytcOf9oL5YyN40Fdf0AQ5DiTzAfG23wvKCL
528F9FzuIheZK2So7PJtkjCXd8KWKWDnm3X95XjlY9al0oZSdGkD2VH4LAmHbPOFaaOw6KyHc6X2
Mc30SV75Q4vwSjwfXuQNS3kWx0sPox33OBFN4SZgtd32GJF6TTJSn2YzpzZjHRIGdo8Dgg49bMn9
Hphs4qX6gLixA81KppFBA05NPkOq8L6Qi5xhwnnKE7J7FEjJKPKE2bbY+JD23sJwl0lXFMk7wmog
8/ENVCnu92VpWkHp9m1tAZ5jIHwkPWc/MNqpg/821i71gk4QnTipi6twLgxHEUG8N2GOkZuvgVdz
EhBpm/R/Qu4bDpxvxoj7BQdJp8Jzns8s38fcAbvs9RAu1w0JNoV5FWxRSuBhYvalDmVKMxmtwRU8
G42amw78WWyr4sYQh+p8zgyVmnkDbrZM+pIkWTEMIxPj6bvpP0pJ6tKLT2FSh/sjNhj2AtRvtwq2
+QbCG0cisMA3SMyyCIFIWZfsceDSaKLvbYilqOprMOFuDkTHNk2G/QZPvPOPCwoqioALRfQW/Dg8
oD6R1p47qIMcxQYGXa+sxdV0O0Cdvr5Nl2cKE390Eskk5bFkEFaD5pmDks0UZTb/WnLHIyOsphFI
e6tInQQbLdi+EM8A2ZXiKyw+e0zGm3Al7AlMNjWNK//YSCmNEDKSFZO8KCKm6WP/7wj7nSvMWjTL
CsIRjrF9eOu42xcWv0Vp3AZK45cCdJZ3s/2VItKgKJ7/H1pAZtmG9jH3HPb13KsbZi9TK9RoyU6F
98VaZYQVOj6nv1YW+qFhdN4gr+/BwNj7CCGes9HaFdsN7zn87j5lqDq+nRXL8Tf3I2vHDSLM0jtn
myzQ3/g3+CiAk4sSBaZuDsjAyjRPaUTWjl2RUcZQ4SbdjUGH+9knYDNEwGmDw8wp5l7sSyRAnT3b
yBsCUXZ5QNXCTMcxSdhP0bElEhdxpCQqf/KvtxvE3CaM2YpFpppgoutct9kH+vNO5e/idqyP2tXR
4UEGmM1imBQZoTOiozn+W0m1aeXQg46JuZIOBNRjf1WjDg+JQ4wq0W2hnzAz9bQJr4cTBJ0YTGgf
iVeMQ/iY1eFrPCfek9SYJGxRBOuvb2f/N5f2xszXHFMac5gSZOwIsu8ddq1wa2TEcMPKqPGZtDnZ
0N0QUwjMe46AwVeAwEiy1vdPEhDT9HUeRnVjhtsMAdmHGphplcwkhL/NdKaGLE1t5+GScCRewDPk
CjgnBEBJg7qh9PfuGjsKaXeO0LQEK5rZM6nwOKF4/KvUqt7ZHxMJyoz6VMB1y/dRUyO9qYMp/LZD
zHzxpTzpLdL3W8TK2mHHaJ0knn82xos8/Jkh9DsDMZ9618/JIg/WNFNvyY1PORxnYXkncABN3deQ
of/bjTJmL5CELq2sRds5u2ZU49ntiJQ60EID3+0LTYLUvSZtZK3hAJ4AvH4BeUkVjgpAWNZRJjao
96nxXaR9/aYNNUigWkVNa7YfKoHZUucwwnoGk1bZv8iw54xSNOPWQiD5ew6xeKeBDXN2OjaN1oDl
5qMrweJd9fY1N5r+HyZQnjEBXEmV+fhrFBdSuLljjNvjWJLo1urhn1lgXatubLNAgC/3ThBghW/X
kD8RBVJ3F3nj2Br8iMkJHa5I4DLJF4Z0GAzN2Pb6JAhTjEK1RWckERnO58FTSlzRigq713lvEoqs
Mo4mykb4o0igtyEHVYYRVCQ1Z+rk2IvwlBEyDjt8PYd/XrF7i3ummFatmwEWY5a5e5a0UdB/RDq1
wbHdedNolKVO/orrHFBYoG/aBqaoxN/k8H1uM4lMQNYRE/yXlBbLJvI94nTXcFUp7QuWN8g2paVr
0ZciS/uG/odoA8Xv5qepDWKNxWl6PX4+OSoic8gL1N1fAlhnXWXmuCf/WhNzkTxTqP0LwEayIpVD
1GjYXS06SHWquPhc8MaW7gure8qC9e471TIH5kh+sOYw7QSyopFLwgQkNcIL6ouZLRBzFIHpYlBN
9oc2OPh90UfCW2t/MrJjI7LwmKfkks3DwJCg1HxAGnSgScDw7aXjlGDw6jlNFv1n26aq//qF1Wzq
KHkrU5JMZmGRFToQ8k+MC3s7a+X7imiDdyyRTSFXaP35E3Wg++k/BHsdyilV/uzJOkP9BeJ0QlKn
PTkTcg1fce99vtkxfprvx+KiFFDvBrBSFqmSMnW+VvOxXQ5TByXRKsmLahssOmCd/MkOrAXArH8a
HRnLNmeWxm7/4v/mDdQmZsF5wIfZSJ4DhPAbHJwNHWot49P+zmo95/QORlXv6PHjEpTfNs0B4T5o
43N6a1IjkiwnH8XQjKYq0XSNIRo66l3CUj1J8U5iWhda6KfKen1zKN3tBfMw7VOlWKmWerSmKxdR
E1hHbIBQsdv+sBywDnNo6v4e705r46FaLTzU0T9+zS+e2rI4MsYplfW1pxk0f5dw+As0Rkwrm6BA
iJ70xu/O+Xow043GpR5txDigFQq3rgdn5wAHMsQLjVoUIeHHIUBslI7nN/6xXP+uQhffkehHvttP
NU6FTPj/GBthPZN4bowQqpa/wV7xQ8MbPSScjKXL0jScKeIuzq27ZUWsIh9E97C7su6ygni6L/RA
tlFMul1zAc3WaRiLn8MCVC6IgEwqpHZS2tTm/1b2HKZzHwlUVEww70TsZgbqdvTSkxR+ahqixWi2
MLxQ/o79P4vh9SkUbmi17albdj8qYzZhotre9pwj8voUhp3PUGbEZSFWE55vGCYP7aCbF/1ue8SB
HEUdscVO/Up6o1IGssEIDU6mdV6Xxm3xVqKfqRzfb/IkWt4RVt2RTEZdduS3DtmDycy+K5L1RhBp
R4/RSciQ3F4CQRMlakecnnlhNJEdiu0d5UBukhL70Z+61LG6fIkh23CYxrhCoUUmBJ7tmY02PVE1
l28frGuJQWJJtRNIGEXRqsw6IaPtjUViv62pFppfKTnpqU03/1ZDQHpRTStwL1+oypKlbkmyllqR
wBVRWh6dP14fFHba6e01q+PVxBryaWqdl9yPFp7lbP2OT/eNZsQQKloF/tqJXW9upaUPzbYlUHvf
ab/0HPax/ODiCqrYSMzSLKEaGnUKf50zX9YpwulPRXbV3dsuEHEnMvnvdc3W0r4R7uulCT8D2xqv
83B/A0Q6Z/PqvF9Izm6xUT9qusH/bRRkVhHbqYpUZ6xArNGA/PUj7b34SNnVGOKThBk/vQMw5ga8
HCLl061u475YEyEdGj1fq8PF7m6rgyB2K5movKJGXHuewNSWsgEunmRO2WrTVdtuOYpdFM80BKeU
7IQiJ4nfThVSRTkmANQsYnxGQNyBP5TywoZM9/DKXAcDGMn5c4IQkDiMOvK+DM9JemZzk7j539hW
G1J1LYsGujBWJv6YLYrKNXCmpM9iA3Ul15r/iA+qgtwAqLdepuPhNO9ePVAAeD06qjsD5JemVR/Z
TP+1O5052r+LRDIWLSzxWYKi0l/UHzAvxyV+LnqlGwwVZ08iYvcal3cqysbztjYCQy4K/zLCFq4M
UBW1rCDUQIiFwA0uSpfAG3QmEdcwL6IN4gaCXHfe8ai5cVoue4p0WE46e5/ieMdk9e9T8Y1+S29k
4+FPBe0UUseg1NYjf6Hg/8iJvntmN360Nq9UJE8WHBuZsU66c3wgjGbMWgQxvhO4VfVCPEHXjyXY
/r0yJNYXFrI4abnvzBDT08607MqL/PLnr4QPu5prFsI9bdH3wqfCgdGPbAJBFRrRVWwfw0ac+QWO
Gtq6vKPbbvFX6t278sUBS1lA4Co7Nyc6uCaulH6LyYsfWpxxzING4CKvJ1hf0OCoiolOxW7W7QbF
RLhIgOmoabytE33peezAhqzNLrpzSHyrpUFa8wYgkLpnCNXlAHNK4plPuVukYJ1zuL2lWPMJ114q
6LvykiPWJFhWTwtrkc7HXUhia9GnxfVMG84B109XZQ23LrOhGlkIaGYp2TH6zTLbnpRUIRT1A7c8
zY0XBIgzs58EOclnN+jeCXsD+K/j6fTD7jszstHDwH2oAZRzPQLNCFiWcDJNK1TDGaW20tOjvJOH
Qn6VQwHcGD3+tgIQsfEytrZ2ahhnjRIk0jZe9VeY0wO8v9lhTyks5O9bZ6QFa1ZOGSLvFuhTJZFm
DhImkNfyU3Ir4aZl7YZbhtwhgTjcBSb5Llg6nNswA+WFj0MB+vRWkIlgrI7h21TBGme2bXgy4a53
ilofLhjA4T2Ca04DXmM+lj3hKSqCGsfbhnlZM4EhqNkW8+1NoZAvW+zyiXXcy7ZZ7XV425OO6CO1
/otvXL6p0teAgGuO6388912oQL7SZaUpPDlMHtWvFMNVMwpdR4ferMZsJxuNYX3hiZnqBfDMvrf5
wpuLLSsnW95URBDF0aYJ2mzB7sUyvjY81eqkcEvhdgb+fFaA7HfEojYJ3rHLiLMcfsdOTbI8oL7Q
kC9LlO3VbAQBWIUSCmnelk7LGzxEkFaFvCpUlHjziC68RSnbNhCztG8LzYrb+fBsvWSpoUJq+0sI
nFpsvMJqPB5s6tV2sdfEhKhUJNdVNsz/LLBcRIaXePmC1OUEwK5MHMD5f4hZX0qQwZMbhQqQZZSY
B9+BWCdQnMSTVFF6nCBu/1Tc+dFEZEJe9D+q/W1wxoTMcib5R0vGH1wfpOggu+HncFBagVrExy82
x221Jl3haNL8QMhCEAj15w3xvArWxag8BF6xaSaq3wZU0EfR753L3unBgeOY5wFYv68fmeVMxycR
t64dzDUNJdyZQsb+ZW0afJL6XUPgJ+AhxeXtxv4JsKqosfiVdHu1M0JNQkBBt9isV+HO/GDeMvzl
4KCykN6AWyi1a3kchP9+Gc+fKiZTzfQCSmksHT6us5euogE3jMH32spkQm6WFrxGGPpH/4ys7APc
HVSPrH0iK5cNVtLbBegkbe2qsScUES41o3l74qOluR682CazKIqKy3K1gy1NdAvm0JvebE84AN6M
6lq09Drfk+qIC6RyQbvLldVgfoHVFJWSSzrX1JTA2j6ldB7318/E5xH7VfQVamtB0HjJhzh3IU1O
6RBITsU9sYjOELYK7/GarY+SWvulkVcDcJ+jkYg5BKGdZVJo97Q5SKiWl0XBII30WsL1VyluzBzx
B97+y4oBH6QSz00g845BIfwLOSPUmALjq4TdRVKIkcX9rwFGTBOvXvMvf4Q1tEb92DDubz4c2Hxa
MgiORRK8yLnGm+L7tpYztXQih6/xqAYtMweMIVBqa8dJX3B4u7sIZph0YYEuxGbRQTaLWLbkGmgj
0SffZmdIk3n+Zr9So7P9MqLKN9CzmCsb6dxQqbHY5hqpk0mV/Ju0EdYiaGN/jtpW8SB/fM5ZppGt
rGZ8hOojO2zODTD9Vgw6mI7IBXEVU+jbAGcHh/Fq3pXmD4vpa8YbUyG9g8PogJgjKdTsE/+4zr6b
l6GgKYysfb3InMOlLab9KQ3AOwfJ9WPjTsdo/SbwZIhHn39Yfk7M04MK3uk5ceuarPlmWC8xIGZo
KZP3pgYxxWZash7Hs5gQ/lfvdA6GzYU2mf4DkcJNNOy/+qN4qZSAqeHGf9QEX9yOvQVtbJF+KXLv
rDSS6OvIiL1kE5y2K6KyJmaJopRoc4oRSCXeaVd+cnusIrmiV51idrQW5/1XFqRtZPt6N8ucaVUZ
/jxSeMlud6C9vJu+rL2jNUOpTghJHDtYHDGAYafj4xWH7C6Sr+8EdPqqRh72T2vW0LsIBW+EtKH6
0P/up6RhYe2e75VKHTaVLL0gcYuZnjAQ5P4mHRah7oCjrVBMHZT4EFuBha5jH+AZAzqotXlX2CKQ
+0OCE/ZRlcoa6uYffWbtx1skDxJ4ynrS3QX7JfTy7MfYemuqjCAyg+xPjpl+/M8tys5eLydIGaS+
L5HwrLo4VZxj9f1044ADJpfEX1M0tMTmnWH5La7rux1sPl2xo0a2u0WxkoPE74QLt+65lWt4pVvW
1VZO1R4ot2bbTDTf6laSqHkfVuefi9DxhZ5owsK/BA54Mi/pkMCpBYx3kPHr34X48x9n3Jb89Qk4
MtwkL/Kd5+K+OI5emXh+g255pvV9W6z7KnDM51a74vy9gMU0Ahs1fpiKhZcRYA4Y3CX5aAiTuMsn
S8No8NxkXPhz66csZCZskAHAS6qLJ5XF76EG2VZs1MPEeO3FzcvpOWXQCkqh7VlNmyobh6eRC1Gj
6AtGPn2vXe+FRL53JyixqIjUEyI6PRFQhcU8wGknMIZFz+thuPDB9SvyXbtt8xNfkyzr/UAnrQQE
DPDSiFdgJZWJmNgaWLXAmol75fNDycCxVRuB45aErgeMBHSq3D5F0ycgadSTZkqYd1mJ2vmG4rwv
UdqXkonZG/9vHTipQeoOA248OMr6KszHCorcT6GX9iftBN1W7RFb/8h1/gQVuKjpPyYQxoRWHeCE
nWocJoB2tbWT9tUGHwAb0JtsDnI4yfcilrsUtZg1suC5pU+nTmB4xg0yfD2ZnxMbd1kAUR2yVc2I
5rhYmODJpPOfAAFh4ifOIymNobbSroe/Py9y8+UMwzIws9s/GLCcoEWGkxjHHoGuwWBWqyWYootm
D/j2geNT2lc6uX2TFIPdDimRSoK5rf/8H+PhAXYLfBRkVp8akFVWuHUFEQNpIk+CAYkzWRGa+PGL
2xdPungh31b1EMdkIsTogxLFmIUEX5mZJhYwwx5rw/O0CRM2PRTNosiLYhBwL5AYGh1SuoPjxKEA
WS6jn57TFI0L9uyTyR0e3n5UKTJhhxLtH88fmtVwyVcR0iWMq4jADSEFPEIh58AaBb/JcSrm+xaQ
rybrwxeBgkQMJpgVtDMkWALNpqPn7ka6OhEBii24+SZZYmhN2bTAe1L3u+kR/agSE4bxRM3aQwVA
QQPDVkSJeQN9dFOgWyjbPukRZTLWG72dJHyWZzgv40CsDdSs0kNBNkEJD1y3eomso3GVwkjmGcUW
DRscN2I6FV7WBUl9voL21NJQ35ZyyIMBQkyoDKWMk1zEpEvw92IvoJSPSpucyWAWwRlGAIpHarYK
/zM1Em8IJ7DscC2qbRkW3xCLGRN17U24WEBgPzzICOMn+xHs9FYsNqMoRMqi+LTcKfa8cwktSjcx
pD7xKhaoKVGsDkU81MdkZ/+Nv2bd/11/tOWyeswdkHNsaIxfLR6+XnMJ6SJDeYUa76tmf/DYVzwN
uHlgEsBS2VXcMNKP1QdRDw+tAxDQs1YADaTrffB3W40r5T8W2nzLpqAA9Ctf7lc5DONhsH2PBdNm
+xT6UcvKM1Ix/laV5zJwZ4Ot/neXRXXBuMQOK8ohgf4nrQ/oe1OdULV8LitLhw6yN0y99hPbRNds
eybaq6Gxt2mA2//0XWs37nnTa16isFFJq3AXKga/AmsDi1vEJCCbj7JE0JZDlMpw8ykxoWdP2F2n
Ih3WZJAAh+N3lG2mmGon8Ag/4szT3O/JvQQ6Z4WK8NY2FwSsTdaDVd1OKBLe2jTjsF3i1Cl1iFXK
MBLMdQKiMWE/Da29QQkiSugIm3IX496570+LNY8dKuLwf26Sw0TUN0JPDxDIZt9o4Csh4T/V0hc+
Wi+9nsEKQwYNdldAR8PioKuQZmuGeMx8JOJbLLiQPGI4aFiLgf7dOvQPMdVVijyTbB6oQ1XimYKG
eAyEqwOtj1jMMeAmvjtT/LN4PqvLLThOJ5tRM3YCdwr4LMXXahPoQHHhXKKI4T08GC85JDZgMzCO
cjTiFvi61vc8UG2pwmo2X6QjVJGwiIjg4Vcyd8OfmCfPDLEkYnLnWHn+ufCxKGj1ZxafIgV7OUvd
l5Q3qz1Un8ozNSmo9Lsg6UAMuUY0WquhekLEMAbNSR0ql2tSYOtEAP+C7ABHH/J8aODFAwzHqABy
GXJSUEcGLTe8KuaVuL/nOufI0sAC8HcS34fFUs4S4aqnjTd9ODG2n+g5Ty2bT9Bd/QbT4MYn39Yy
ZlEDkNyn5vKKkqwDOlssi8krHy5msMshpY030Pgh6iVwu1+dShYn9O8NZ/k2ijfWul7XucwSpZ8P
RQi2EqUp7/6OARjm2kMQn6Fn+ueAyAVL6UTG53+ZbS0Q8aotNdwBclSFMNANFlCx6/h9mBnOa0Ez
aU360/h3Xd2ZCp40SxEFywKVZQDqCJ33i/Nt48O3QofvNdc65sfXJZApgEU1m26S3T9qHzLUMqSz
9Bu8NuIoc/ptvytX0mk6NiDAoF2G958QfdCkY4lSxTyTcmu360jV7mBvP0Sl3rjYq1Ez86TfoxyR
BNYoE7aTaLYY7VOJ/6jJ72fC8clG2FcH3Sea9nFb/gVPnBEf66JF4goLRc1q+Z0DlJrY2hhTwaPP
jR50QFNptOHTO81s0s+2k7T9ZAKTZJqUrRnOGJKbcTQ23ntQQrHcBxRtyoRmg0y4Z4jzbSUvcy2g
tYav9kZ6TsJZF5DXtCBxQPk6YSFXYRc2K5T3Lvqlao4OtdOQ+bPY2ia3HWXKskvdG21zha3CHkwg
b1br+DHGEPYhul/ilOK2bOorWeUkqjzg5TEmYBfTucNq1qI4f4B3HFB/ltDmmVU8i042lPTy/5PE
W12N4sb+4Vx1HxCGq4UWgncu173CBRUhi3FySZDt9BL+vA59M3FNMCaa8K4yZWfGhZyBa4giJuLc
VqPpXuZDV0lGvrNHyjJ/MbUpGA3Ynl/wa/ups2CXOxVoKP+n2K8AhA8kNxmuxkZVybD1BnmS43Go
FXuDwxX0+4doMlRzROvAUtYSf+deJh2Sf/ewZS2axVJWv90XlUqrtu2tzmQtdAaUQbvjryEG3/+/
UvvdCwb2I0QMNPoAgGHMBDH93BqMTEgy+sdCW4fDtojMWe/iZbemIMf+pCS7JG2VCHlq4daR1faw
ToKtFzBVQk/cFpvW8j7MSDjSPnZT5DsKgSEDnVulrKS+zxTOUjf05diHMBubW4OFtbzQywh4IMO+
BNZPSznd2mxyjPUzPd/AgDpSCqfa9RRkeEHQPbuLV26mI9IY5o6pAW+e0uDXjcYauVmhfa15MlLi
Gs6X3sCq3mAV9uApwLdksEvgLbxy3Pi/WF5Guti91erPGsW1y3hgfb0c7+9EDDGvUfIU/SL9fQS/
lbEAw9QrrIXV5CXSV25YRD26SvZvNzRPFaQCMpPTd+Nowpd/rZTjePga2eVkMjsm9kQ56eSI2NzW
JHNQBK5C60TiyAliiH9KKeqODPIRm9T416aaKgEnysRY/C6GtsQmwJqQy/UEyAnMW3gV5ofdIuYh
6WecVBwTBvzk/8qV3lspeZT7hVkCXZGRkD3YRfW9a3YCmmTkSi5Ed+g7NQx2jntfMhj7RuhRCYB+
Ub7j9Yd+uEe1iBsiA2TJjFYeINZdmrx9R/mPC45gwzAtI9H1NOhqN8jp8wSjk1iym9L58VJzqg9z
Duq9yY8wKZUXSvOAcsLfjskhrolcrAKVNRQq9jXA3MYts/odU1p83k+q5OrZBJrnTPyHbBK4xeDO
E3N7yZbtG7qlrkN/BcCxdot6zr7wvYRiefuOYdMmfQ5THi9r7GhdTY14+Km7Mk52m9fq148ziUSa
mZ+xeLrU92zSaXyv+NLTHHBreiAWMVjOygZDWttvHms8ak3zs8ijJLBc4G2jkRBI4+JOk3QKpOx+
hW34QkahGRdvNFRnzFFddo3c/K8OLsIQxtWJ+uNNTknIAJ05MMeuWoasO70UmR8WHw5rAbfq9bd7
E0s+p/89Iyuve506inznYPi0+phnxrVcY4EhpSu1lK6JztL8BIw7F6MxR+Hud3AIdeMnBmnAPWPB
/+EfxF4Srv/SkWVAWzAjrqkZ2AH/T5XSo8Sh3TzwHKeW04NIm8V7ZAFBifyDxS1Rp/OUWK6oPdj3
4C7Q2w75sPYI9VNNwBiuQGpptbm/992tfAuXw2sOGwwp2wm+Yj4kw9Nv1gNp4Ncp9jruuk7o6onl
xrc//EbkcFyCwco8qx0PhrpS8dNA4p7L2pMGgRXxtb1PZ2aUakAuLfHlqKiKT2NEeZ8rlydyvvwr
6O6CX1HCG3WDY0mvruymZ+9SdKksxr7ixs09EGlAAYKg4hUM0mxK4j1hETdsfxD6srreD0V8B073
Li3xZBxoWfJz2mmKXf7lRMGxAGwQjcFONGCbm3eOjmctUL5M3t4ggFjdG+7LVJK9JMYb+u/BzX0w
7HuZzqQ+TsM6gQyRzRgKFEEEulKB9jihjlVguuCT7gBlM+cpMz1cv/NqCAsjJCc62JGmuPJQMXi1
AzsmZ3Kh462+7gC2W7HHfEZ64m7EmuhTFtK+iMXVQwodqPaw5/P74LaOZcMFo2luT+bX0SbiZVkY
cDAU19nnZy/UF0D6RrJu3x64LvbI8CTZV1kWrgWKTNyvc938cbuL9NGBwOMCwv0jmtV3wKTWLYIT
3kD8Na/KYJZgyrgyCBJUkPyr8Pc9Z6tYSwztI7qwM/6n1IRG4I1qzs1cYbcMG33NbOHjwxI61VKd
LGoz0knu0uavGLL0n7b7k6+YUMpwL0vx3oiwyKifReJ0QFF9AdPr67R9JYVs56NIguOtLzqrMwYt
tJdkStZk69DnDrORgMwq7nvLnz8mDQYyuHtnoSU75l483IvHJ9828V8wGiNBIc6YZBpDgeN/2/Sw
6RCef0+6qeikXcYUIvk9z0hXbi8uCTUj5lHrrNnnECljV0M+l5IxDZkdrq6YStd7p2wbfsuRh/Na
O0WKjSlvLI2WB3z6uXBDU3KVivcC9mdOrVtVc5Q5jjU72ZDd/dzrrvKf9PZZmCb84MszW6GTkyWL
yPNfL3QqL+vy7hKaMo7G4I0xKapIfDVHO/gyisBlfMzZHkN4/xI5ypsbMnajkQCuetucfZAXAssM
MQQQCyfe2g+kAP3rPGFGlEj2EfZ3V3FSn/bgPz07vi3oT7y6V96crmVAURZhJZ67ic+GMMKd9WEh
TAHj+CqRpGgAx+EiLGEnbsJeWsrr84Gxv+ouik3w8W8EwclHQTs+sJOHq5Fxpd7Ou4Qly1pu+OoS
mow9hlXzvHMrlzB2nbKRxY94QsNJPUYwtedu1m8sdxJdcGfNXgTEOUvAn1ByVN0w+nUoEs8iGRHi
Z1YhdyUoK0wytSMbi9S1uZ58NzckNd7SEvbh6RF/Qzm+1jPjlH7ZmElkxncmCgSMeDfUGk70C6OM
AdliMWxU1kkoIB4wAS87TI3UkMHDaLSQzPwlbfcLdsiJughHURyVqJbiSEAIeBQXwWXw8+7b28WF
Tqe1WFmHWpOL5S+hh1/MajMqiqDCDa5WgvzvEM66BYD0iUAs01C6DTB11ub1k5I7P3PkllNv25vV
9EtqSwXu2Y9ZmgqczcZ13zO8iaSU+ntIDnG4cCAx1MXXwDafXiOCsQ1YZ8QGeG01pHGdCRaqyBZ0
Y1Jem9fTukby7IPgbrDsyJQjeiXdboLaybepShW4wiHiwkZxTriAQ5CesTgHQLmlB0hWh6IbEPMe
nUTZPONd2QR7AQo7FU78laJITbeYzk+O4PZG5xo543inNa6HNUjftMCZtmkwSfryfMXoGkuEExND
dewiwKIhUSE3L/En1y5HQzCldCScSmZB5clVNxEceCiRsf8NkpiU3mwXQQ7qvFfQwH7zImm2DJhk
mrwEGYhxe7x7rxDqUtoJnqyffZHkalYCFUXQ/ayTcSpIYPO3lZnnKppZU1WvaY2CRNauX0g4jnFG
Q+/NElEUVIZunBtptAsr2eeiFemr2b8mujplJC4Xhmq7QcgYPWIYEqDs+Pz/xl2vCqKa51DKKYc6
Q6CeIzOSUgZouvjs1vKT3mifKW6YPFkRcXBbOYdcI062Xj8Ifkc5rGis9wtseRJvITcJC/zwaOcC
pfg+Zv0zwtlhiWnT0Y8M8kkGoR5k0SAL4zlilUKVtcijmTQdEQSeRMKv1/X1uHoXnHDeNrmdT8Ep
AXls/xNJvAmKgR8TILZPF+8TF08dQWjo+QBUhbLO2BMKBp9+edbDOZSkKr8fHGCtz5eIBE/ukNZH
ArV8R/wI90v6A4aFUcSpwKU10DUOO81py+rzOp9pdE6BnhFExlv6FRzIXSvFEyf37O9sNePl/M17
nMIfNBSDJYTfHBgKjVJO2qxUwR57aqICWIixbie5Q1ar8VqSDhYhiM9F1lmBsCa19cTsA5eba1ZA
zozHu8Lk/t8SgZJZ5/eukN8Lc/wO9gjy2DSxMalj6NXbAsSk/p79YQB+bK6Ph3iI/rM5OVw0m6Yi
Cu5J/fVSAOib/t3xJJtVCSElDlqTmk3dCd4EQvN5nPD9HjMnkNXlaDDgr77dYxr0Xh+CdOM2ovFO
OiC0F0+oawgTENuNgtw6HxXTGbyrd/vzF5HmbCCDgOhy2vhsSjebNMGFCKS7TzFiML7jXgADVug/
CajoBxtrMx0MY4wPJdJKOngDvi0KXBCAqEsvWDRrVrSS9o69yU2QLytXqYsrc2gOwr58Fh9u+/t3
5Vjx889qvSuQnyrpkrNLNbS5A5gV7DhsiK8qhjZhFxaRLJV+WMNLGqrM6XAk4CUHjRghGWK8JsMI
N+GbRSugg1MPc3H+f1AUK4HUyHOWUIYjAyWCm2X050CUy7PmASPdSxCGjonDnVnISGgjM0KPQI1Z
dcf4xqSKx8+2c8DXJnbR9H4MGYw7rycVrrHKMXG9NASPe313ivByGgWVcxKOdbG/zfVoZb88QF/b
g2j2mVdGGoJjaW3qfTY5WAWcaykApwCkUh04+smYsITTOcn04049+vUInOkJ2qeo6e2wIbk/TQca
jrnl4MI+fG4HH9ZA8KLIq64NZFkRcPuxby8Q5zzYR4OZIQQkvFEmevwTMwY9wDWrpcsaUDZVe1MX
/RMSQPEvqj3iVoQd/MfzHyBPen0iSgACWjz60cXGKlsej9V3Y6XCo+chFGDuipxuJwGtzfXHpPNm
3spQCfAVEOtXhaGc6uKVVdr+EpHXa2Y3xfDuFwm3LzT/5fe+lhfVkuSFNaGLHR/TTj9HrvYRBaQn
Z2FBKILuZ8SWrR7+LxNkv0ba/a/WaWWTI6jgKft3EwJXxL8PT9nE6fPx3sVzXWgMbW+jtBnIOHlH
PsTaAXUawhwdO7gyfm+bO96v5i1xaYcPPifEQl/+xvX2lgZpZKkL6v8KS4DiyhhiugaBGPBFgb8O
NbH7g1QBRhz7j0zGwnuolgYi6y9JwaiqQli59sZ71rbKFcAfkLm0rGtIxlzEH2lQKqpstqeyT4gv
tUMsVBDQW2wNiwXeaFu7MdQKxljG+to+mGG0jWez67+3ihT1CNsVpmlO7uIg6jr6b97N1OOo4UKt
lgTXff414pGNSwLgub5WuLYcB0Myn03MGfVE9ku56SjZfB5pj2w+K77rmMJN+/MG4FroEu4EqPez
9M7rBhDizJyM46dVxMk5873M80KZegu2iBhEnX9s5fNAnAbZfojpP1zehwoVZe/kTNZ98hsC9T62
XHl7mYY2hDjh1o9GmlshUwkvjxJjM36Ylqs9LU8TcfA88CFJfmIvhOs9LRkusaBOUIL241HoQM4Q
RDIhM2f0aEpA+ZixtuVkiVs0pEJxOplrpID1+u8c3Z8JAowg3TZzaR6wlKeR++WqnkuURlX713eJ
O4sOyV4ftRusUSG4vLdVj4Loy8bMG0mwOhEaW1exWmD3bSioS+0evSEMIxKmyztx4xTNfCJpPrep
T5TbVFcDpVluhEWT0OGO6crbBNs9C4LMT45qXLTNTT7bLMBBEUMm5yTFfUR9h6awlCdIrfsWISwN
xNvDk8PRpKEsilUQo+xYOoT14Y6iIZxWz4SQhLRd/AieroXxTnwcoc5BYUF+LbpHcLqHDmv4pZ88
lvDtbIP8OdeJcdNgiUgkVgc4Eey98CK+rNuqGEA4nwaY8xyefariO6hP0p2UZSJXeAwZsdbiMPf6
dmuhE4ETHSku/PIThwAKGllx5QPdVuIX6p1wacORaqjX7D0IXZ033ELnnftMND8hkVGTcIo5UiY7
Ic70UhW7YZQKbLDV7rH1GOhtYt0cDTJdMFfw6LoJHYjwvewquLjWpOdH6VJMyq9HIrUmQXzci18w
TcybLLtNlK4BHz8iqcnYTRsFkb6TwGHBpuNDn41n8vnHvxjfPes7MdYkzG9k1uMRT6tHkGcIsBA4
yo/h9YxmIeySpnDGLduFVDFuvJw5RjTy1A8cKD1LZ3ber0i1SH59sXHnHGR6nN4IpkLxyHnhELYp
lTFdk3zvH3NTyYPmjxas6nxM3mfGg94tRnlEqPtxTeI0WwPWBMqvEtPYFTNIonF43Gy3+SZSg2ya
lBIrBZF7iWBabIIEzH14bzNl1+duqT7yvv/iLWPbhBzEOb7RCqm81yF8KAVWjD1K+6G6JN7b+WVp
WEH5dt/IFKrmM07Xz9a5n+GZTsZMan/xfos1zjzcxSIQAtl4f+v7/PbDSfB4i20OpygYNmTSOjUv
/csRvyDKAgs/3fjr0Hkes9NxNBdFRLmo2jadmQgkaDnyINvzWFy4tncWOGwwKgvT06Jsy6FZ+C9C
yNYSaLGGO0ERky+4LJCcB23c7wY0JpTnSGQ9QXzlbegqn8nfi/KdRmv0SmSz7PdhpGNu50YcF/aK
CHw/1UCdn8nOO63JYaY+a0W/4YU4gem30R1x6J8EuylHqvOeQ2bnTehAnyyOjyqMtp80SvYN6mDQ
798N2MAILWGqAuhbXGoG+oChdgpU6cF4JiJiecTi01wHxUoM9XmIhcWKEM6MzUMiqBlnCXDAkPQu
sv/9VJAdpwMxwwZPuUrGTv1S9uu0VjgsGO9WazTw/amtqISROb2N7fZ0gvbuFibb6J85aRdmXwVb
9ewvbIxS8ijH0mXL6K4CtXfQs7Sow/AOS2I2yma36ImZBdgYHYEiKPrkPPZK39+hIiSsjSOv1T5f
Nhxpj7xVfD6ZpSi69xhos3sk3jI/gy0/Pii4q4xL3/v7nxNfxMgjMfrL6hPag1SoKAQ+yAkozVef
y/1vMeJhz0GQgjFSziVw0AxTlV9BW0j892OtR+dz1Y8KkdTdXqVZXHV1hNCAXMJeSC1uXhxs0cJ0
F3GztvWen5zqLgidg710dKoftsa3adaJalIMwD+TcEYOvEEKYGxkt/fwQRmmFOU9KrXrTYygPoXQ
ZPPS7U/4ff9u8oxAAm2pg1nYbS/x2gZNIu1h3bySO9Qk8AVpP9oeZKYHHdxKcC2XLTH8Uv4UEgaa
ggPkPhmvPh/ImSZyz7cbh4slmPXR1+0TT2msoCi9uF1c4gQLVNjyuFtatPh2hsfbhbETtV/Y1n9f
+gIAwhQtB3l8uHDYeEljFA69u6KOLFB03g8JoSSJc9aUtD5F+FuZC+NxJEgI8aBObUSVm76DRF1k
ocPQfZnx7QV9owSFrDpTEZK9h+/nLhS8QC84bAfDI6GEYjnWNfNRm4bpzb7+N8DANRdEBPPU4sre
eMNC9U+GBDUKnwPVxeI21rRqllzDxMj26ma2HWhWSetw3gfWIz5UXoshYBOZV0oCSpyRiM/LA9y+
EbPEJQJdbpnU05CmxexymQRxtYK6ddQUtahNLWmku9p7+UkavVDkrIulFPwbV09i4A1TVntEKc0Q
UJH8TJ6p8DhR69pt+9V6IQLhG7Rjr5REusEDgCY0uYA7BzKzZB2VqdUxOwz0SXgbY7tSYZ1TYyPY
XS9xGMxnvArGHl8gldBwRxpksaAav8tBq0KtkDjNzOiUdb3Qe3clq9lHcKBO0MBP0H1LWa+GIHvH
QJExhQHphnVYQCkyDph6jQNX0ArECwyxNjaSrFkF6Ze7x+TwQ4mXdv+KvgOrVV4XniNbrn7NzcQq
95Vp9xAb7hUH6fm7y7vdfjUCI0ywEHKVXvoZYdnFTaFdDzHdFpKbzSeO42rIlG9xm+AOjC2SNROm
XDVPDvz/gsy1YQAtdNtLjLwo6Ey7aEMjeEg8S7DPb4w3EZ76OiVE4FLmfiuN0S6JD6WofYcHpkJC
vYqlQMOusiXhsRhkQ3xeqbVMaUiw75A61jfCM1OrpR61SBNqn5TKqZ3Fk3dpRqy2SxO/Oi9CDyr+
/KOFasYMJXiv62OrjGTMA6+Vn+W+9YV4YgRvt1jOjykFpZek3mAPYblgRr8Nptg8F29H6KBq6Jyj
sSGBDfShPkACm5E1A0Wby/Nz/VKH7n+ZNisrm8pPFNnwHqyaeI3j/Thm5xCwA89EUWD5EU9zR97Q
yNcyFLfdGYygHLirX4BW2ZvfIepdIfdL1oKNpDuxeKsdw7/wONtQyp+9v7mo0ZFLNiv6Hm/ppxs4
WmKPCrsXzy8JJBWJNwSVXWltfUGTEy+5Po4/kmfEx6SVPKi86l8DTEIug6zbMFrPHi9mgE7Jtebb
dFgCgVTcYX2sVOfO25UmM843UJRg7V21HBQIp2fR8zUCwxdrRpIT09pINP7WBchcJuJ0t/IdE8H/
kn/fy3R4r3jD0dh8vatsL2KSyQP+eoY3Vj4R4lnPX5kGIgyh9IDd+m/YDN8wkTeG1GUsNT8BjOVb
tBg17PJuBQHVKethiVsRY/byET6E4FBjGn0FZiOgrC1XZ5RMfUdlxGOhoi5ecH6gH1NHupiWWk7b
x32ERgQZBFusdQk3W1eibmkKWi969WS6TVBciXTdu+y3RHYPldI/GS3Gmr2d50u3NFANgcL9HvmC
XnL+xNkrWuX9QrkiL75sZrvVGV7tHyJlxYcbCV0NrU+Mwi54Iv2QoMNFWsWx97g2jGbZ7kgHnafe
Ht9RK7VStz7LDd2jgI6uzyXAIxtcpJOcUqW96x0NXutHp/sq8Q8Riy2upOpa0Udccz1GB/SRjCsK
a0PvRTFUPz9N4ltv4EwdOjwng+Uo9m/ZcHstvn3w6y3W3JoSk1mk+tNzx5UbrGwONpzW9oa/NmkQ
hRObtzFQc30/a7aHzN3SP/eucvaWEhwkm6HKqlQT8BmHTZJKyBZtYVOj0v+hvPjnNNX7e2BWN11+
mCegCzgN94eP6ShVuZumIyls/nxchqsKLMU0KgRIahVLBy4H9FQOPv1sLdaNkKyB1NP6T6p9y2A+
yZXdtBcxDjJFoXBbX7eLhDVGaotvdBVGRwD2kaZcjlOO/wGp1q5TpK+QvaBrSZNd34lvrxd2nmNM
luNLY7SLh4ll/1jZ6RUbXY/oI3L0IYo/2yAsBWBsGqd7/tX8VwJnS4iPff57/ZohMKUtZ3NxbdiB
YCPZgyP02Q5MdYk7h2gyiNJDAcCa8+kn2jxfeyJgEr3SyO+vEMXAMsqFGNdqgUPZfstzVA9ZrG8f
na0sJDQrCWvM0ixeSAatg7WI2i+2rQoVjETNh7e62VdnyBbXXphJeoHuO+l3QNcDhFLT42ew//+a
wvyXlDODbUStSCorGZXcbkz/KFXOie2BHGGmKgZhcwCDLhYLiRmRRJR+5/Guo7Zg8M0X7jxTnDq6
0UeLe2Gup0PNVfQfv8Qq/iFN/UQ6vsZEpyQ6LgcMdQMTnu/XJk2gk3F7pLYATI9A7unUQwNyi9VD
Nq39K20Kk+LysE+j24N1amt8NGuTZy4WgWlpm9RHPQiwI9ptTNz/ePZhIg+PMra4mbXPVOs/osum
CNK1vCHXp5oVdkapyXRV6eJV4QwLrB8M7O1yypF0L+v6FrwrmsUXs+W7dvpyg/IEQbB/smMkjd3o
Sw8h7mxAr8g+q9wMKW0dZJgXD3yC74O+/DH5foBoO3wNUzzCVGUDOahJzAmJNEULlGVsxLLtuwqq
JiOEQIMqVyWq9mO6IBcWap0VhYxTBXA0GzP0NSPCK8h5GlEuVAI2AXIAJhHCj4ECtU5Rmeqzeci3
XrjIXYxUajzwf7oYqhhXaZR/wuvR54wpETx58wzfcXdX86cjA1KA4u1MQkxXvPmk87CgUXr4uWfI
O1pNJZ0qWBqbwkpB2gT9c1DFq0x7/dgCZktf0bmcCj37JaFKl08S3f9yDZiqN3SeSy8v1Pas9hW0
oMnwqgostP/zG/ggWvXA77ouyzHdpLyOIWjYxR441jIEIlVi2g8KdHQkB/kQYb2E7Ld72w/FGQMl
4Icv6N3UzW0RXbfYkoZoktaYlLxoBCZ1DD5aSteGYSxqKTOrBKwsiWBly2JbRBoXEgI/BXv+PS+h
Z84G+Pk3HA1h3q0FVautxXsfmCmqRUvJqex0C1vpuBRlB3yq9v6faH65Bj6avVUknlby0VpOHu02
ok0K4yRc2JIT5+31po9Oo1eOgwkFIIMdU3O2IXor3AQp7QlV0yWMWB3jpKV1X0jX/OGL1ypks7V0
gnZACQD5iZXlhOFy6G5GD759wendWkvHxxRJA/U0rCLvwxz+B8HIRbBQ7/UXiTGdBdGwhpaP2pkV
HoWHbnaldQO8lGPEjV8vC3rgogcLfvQzpU5BC/NHXUOzHZPt14xOxcPSmMmfqjjex9dwpoGjOonR
lvY+x17GXdu9dTDyVV6psmEMKUArt6L7qNiv3ylCQ6F6UaB3bqg1HPmvvlz2aOthy2Xa4odYEyby
pnXA1NUUtOQTl0kdJ3PpWIW8Sq2QRkruQKQ8Vfq68l3o1pMxq/RxXzKSAEYqBNXLUfwbhOIn15Pr
n1xR99FToO7NPtrj4s+U3/lIOFWflWU7arZUJbRPeXCUkvKTwsG3LPuKa7OXrIdg7Pmzp8bLIVj8
xRctVAHbpiu4NhB9/Vjd8KzBkeLGDHTVwfRoEIhns1DYnyHywRdEplMfPv0UliCT/W39M+mnxQqU
RsjjeFp7cnaxZStjVHepIOuOGbfdfI7zvv2fEoHTRa40FdToBB3aC4WASFWBpD755SYyg1qKu6QJ
YXUu4EHGYZiGfZrA+BGDbzLNq2REQu4j0LXLWr/3tUqP4O5UStodt2BBSU7Dg4lL5qnzhBPmyMZq
Tk12uDUz0n195VHKbfVU9Diow+Z7kaXIYjch6a1uzZSHFxlT1bVCdHhlZyUn50vJzzUEYnGDTjpc
rRQtyBoiGrWmIKn4Yg8ogrlJIGboXhh2DvEnGhb/M+ra3K0E0lZFGWPuRxOxPnBPuaxv2fuM7ZLk
wx7mdUahK0bgtPMvjOaT3foLiHZtgw5cXPwzKBR/YW2WQ4QdxqzsaEUtbNiClEoyhflckUd/x/x5
CMqwgEVpF9ln8QO0evINDGCBylrTSU1wly8/+lQQF9x6AaAC8ktoSdGgDS8r7559Yd2i0oTQIyZd
xROz5bQ/Ex6QWr/7171CO2PD7RfNYnr/6MynTAcV5t9pg3YP7S5b4DxKEa/oakTnwfGT8sdRdj5+
YfeRDyO7VoWdgka69Bd3V4KDaPbTEyV7eTLBi5w+3DrtIaNLKGvpOABAm8Pl9rBJdkHp21MihkWe
UBypTqHFgGmH/Qaj/Su2fxA2b0tnJUj/AsNshw87eiqc09G7mKIolVSvUF567GzYjH0KhUaCidm5
2SR5dS/4roSR5RxR+y5fj5zzkpMdKubB7QhGivcApY7/e4jCmcdpZrek449BTwDVh36Ge0a5KwSg
ATJ+9h3PtiXPXHhYjM7iKQdGDkqqYPZZ05S2nvU2kMSUGtVlH5fs9hcK98ikf51nrK9YNOJWk7S8
dU9BYuFsLamiVWFl/8ngJdXhEDy5HePNE/BWQ3GjB8qhIlF+yZ1qf6dhCRMGeZROzI1guAKFE/0h
TkyPKwlcZnYegYMLmP28z04fPVhSfxHvJktJjB15Ngk8JD0dPbyBGNfjQOzEjXJ8c5ac+akOhOFQ
7vOenVldwO8jKTXIkX6RAY1tr/uy7n0GmKM8rr8jrmd183gckX58wNPL/lWXbmKdTqPl3XAsB/Un
5F9Sg4ISGTOKs/RakLQ2wyB61argBkidGKS3zb9QQILoCqsQf9HYomtizBKHfqyMgbuQBGhu4Lw7
2Cby8xklTHG6Gyq8e6uNN76jn0TRCnPVC7Vtag/lH+uG85eWeeSBH3Gi3GvF0rfwW9axUEZTeI8u
Km4CGe46xSvkddLODzT6jZ5lH4O4Xc75JgKUeJfj6UuLNXkUi8sf48KXuwBURad8fmG1E61vFR2i
zNHN65tIqgZhBM0LEL12s5F9oaadDF6bqeYHqxpuGxZYx8HOCOjaZnJIWA6quOErUnhXDcyGLJDG
lHIfFDrD7FEyTApVeA0JjqGBIXH0L3o1bemzN7VY2uJw8LWpQSyHkCUnTbrym87eVWkRmIXmLS7f
ica81O3QE0Nmgak5lV9ykMiVCLOaUf+XI2kBSzgkt4EYoUXqwjXLXG5e/aveg0fcc/5wpb54pyHU
D1E6/OwXdXwzLX7bxrNz5TZSPW9mqDO7irlq/RAYu3DnuyPNAwwdjUFruz/pona1M262bd2VNfr/
Q9f/MWojqUuJCdxKboR8+EZvgXMo2ikhNI8dCT4q617nBno71QFmlfRtGwM2r2e8mSOezJj5kVXS
1y1bVw2J2UVthQBN9BZAAXHO7FTWVcqAABpWQiBMJ5TKmOB6LCofwJGDzAlT6uKYcySqKoTf0byY
iX6tOPkZ3AOyDiRSUcZkGjTzL0ocpnZsNcCGGf7yRAnQzMDMRhjb2OKYH9RjJrDWSaliHJD2subo
u3/fmQ7zGYA+FjpxKzLsNPVLwv/IQhJO6Q7k8p1fXXg3fsbknVbsKz/1A3Zlpvh6y7lI3Xvp9Gnc
0f+o9nar40lDZ4tPeES3dSQ7Z9HoLFZqulvgmrWTroyJQd8mLatwMPlrhA4X9D8iaFvPrdUzSCMm
h2LJA8rY1jVtk6XFBe3cUZ2H33drSgH0jYXjJNh+rodTf8GMhkAQjxe7sq/TSaQAeVVmANG2O5aH
glnc+/bOy763/SyTH0OpKaBriva2Afr2X1XS/Jl+enfbG3w35tiJbOZJ0N8BiKT9puTZwQWwcw20
Ni6npMZ3KTKmt3hBpx4gTWwyBUUlQbRY9f5X7AlUJpSakqjghRFH7rRveRAPLQzURCqgW71ART1M
fNZrcPgwCNzzBGUcjcT2kMCU+ICiINNjeXFX54SsiRHg95iLubBn+hPxnf0tYt5exu0O/8bWEMVB
EVXatfdO/3LZFj7KHxYeuS7KvqMcvjj5BpM5/Ws8MjD7BI12sRRAuXKNhFFBAkNQ/arPNH2DXohc
CktQAUI2C3rmqjy8opKGrBlKcwmMP0hh81/hnjGNwkG2gZ5wdOXF2cuFn7IK2qcmWcf1GJsVceOV
7yno7PMHGXL2uVreYF/ig8Uimgdc9BQfnBhML164f62eKvLkZdwX21+ohtTLw5wZmNw376jojUNn
z2+U4iAInp5VnqBKRfZgMb/9HWpgGOiLyg0cqoKyKmdlik2YQQN11//exn7EhP0XEcoYkTLSIZ6Q
AMk4dAbje24vQUTgjKGHZLJpxQecjB5xj29JMuRtqSMdiSlFKUdFOy0PeVzYyieZOOmc74l8+hvG
4Ux2tWx+PN2R8gFV3hlwoF26VvU4IPMZdqtkro2RBr3bmU0bUz2ET4w1AOPGDxtZUnfQAUlU/1D6
qRxCd4X0YtzTQqbEARv1DSK0YZU6xwYj6KDLxuPe1yqzaxmMmKOJBL4lSQpIUn8cBPm/U6+QK8Zi
bFxxk58dGXBsGu7lN5ZTwHLgni7Pb2Qh/yRmKnhSsgyyk1VPMML87UaGrUAJ0DbO9hSDnFXiVXKf
6nQC9dAvxkQceFOuO1KV4sv/khbnx/2LCchMwx2o2qC/nTUk3f1n2j5/b4qKjXzhF0Tr+lNObgcb
3txrqBml6Krv8drr0mp4kh+kGxR9EQSjnsXpNeO17Nmd56ok1xsmP8vXrkL/ojq6E52NQHxm9wfI
qECfYJtaSBlR/C+KRx6udaB08N5WGIR7F/R6AfL0zwOkzf607PGG5RB4L/iyardzdGoLdcnRYsup
DNzqFskHeNTIYL9p8N+cXKLqSIs07TNgSqLp5RCTuATfjckdBBJ0m7QG+qm1G48/qTyFbB73Nm8b
Q0fSvvfWKb4M/NmTZ5QVrc2OESSUjdBELXyj1FCBhn+G6TfgWtdMA0HqVeC2FVP9cZFm+Dn5YRo3
7D4kNJP/4rv+Ol/8meUyTr/Kf6KGA4WrUJ2N+JBbgmPuAItk2KALkZKs7BvL14fJI+cLzUAZlUm0
hzTU0r+n5d9VvE9xAgp7LGeOqEu91pK83g32GIt+4ZKDfZnwZc+Hd60S5L4uJjAWYjWtkwVGOI9Q
Tv1zY0287EypooFhduAuIFiPEOFh/VFXFr3woJbf8zoeD+Xi0khZpb7LTHbcGzDCVWLWN2MNEcEW
A/gENCaakZzvMoqQCpqSr6Ylzs5GwCmt2oqqotynGeanQuchnww7lPP/7HR2ya73FohJQTRfRHKW
wn77rZvsqTo8v4ZQ4Hcwli1UzKCtcia4kT8S35pMdN16yfYJMAee69XdXyJhQjlGThtoSd+zFP3H
x56werjqcUthOg1EadDUot3DWaLApxrpTfYqtfzMUQpN/uQxu0gpHCT/CAlX3Fe1avy7yJg/33o/
4wb6DJ0/5mOJ85K+dMSq2Hvgbm1FqWLHiJa8vllB62FKUTYFO7YgTH318+5Rz0ANroPgIVpMu1te
CS+1dnZ5Wgg2JsQLJ2UQK29KNiPPCStX5khgbHws2CYmNRFrSUmmVltvmsQ/8uK7VLjtfgH78kDC
5Z6WO+r799aCpefBrJwzcyikniEDYj9rsH6nSHy/805nApYRcStIkjATSJd4jnajjaqqnRqifMI/
+a86K0EnSDXEeZNJcqV1JMETSNIa3/nnY80mCB4nQf2cnhU8QHXKutvzXWC9Oo5Kd+Svb2qHtObD
i0tBhnHmCKKmdh9JCihugrdxhTkskeOoVw9EvUVtbbgXGPYQ3aN10knLGnS7brqTUtIyBELpIlP6
NBNnLo+7EhcjDha032hH3NNEs9/CJefgPfymXDRKNDdDmk/2crcKi8uDZug9NWbhV2L2oLXzRW+a
XUqJ05X8E54D/BCde62ZPGQQNpPOR/YRk8hxIja3yeknzRbHoxeG+r+RdHZEuIqI/tEoDKVXKDUd
HJj/VWIXvCzLn1BEyC0OZoS8MmWKLY321J9OG41Wkg9tBaZGsDAHkMD+vLAysnCHyFTPW4yjEmBM
+MCrzcXCE6ZH3cA7VjmmY9pj4zyRwCuuHSvj6nl7j6a7Ux1gCvOtNgSU2QVBUxFBVCpA+/xp3olN
y8FdL141rZOVqizhtr2P3DXLhTca1vuQ4/49rQ47sk1S5elkNzqKVeoiNcee9T1tZYJv013knxw3
iCaJv+RM9RKXahf+EWNRjHdfWW4HrsgK1e0FYzjEN5oezXinwsks9zr/UIjfbfS4x1q9gxtimcY7
qV9xFWaV3C/rwjnPvCk6bvOuvBAwmjphQYySh2CoVLq6idoN6AhYHdocuC6lVKExa/iBBNWpOEZG
YpZU7Q2B2et9vSDW5eTSJUEbZKBZeAVGUtV3ChtuaG2vlJN2Z4zAaAgZyX0RprES5JKo+x1DRDho
C+ZL9XQRYzChmp47y+OFvL5iZ2zYmNTmM1vOP2f4BftjTF9jWjpSKViDWnHKWUe8YM5uKPEaimUV
+jGB4S/CUiCE0vBqntlkE/jmVe39do0GLEGiZmCEN0mhvSRMyMVVLuCfdY3JlI7YEL6z2SN0P5c+
HRJ5cGB7kh+vqXaTgb3XUsgncDbJsoDGfSPBoQMukNCfu4ZBBZKvk24qL34fHZjTNbuaxjfNPQQc
+KsnAcznODhnOw8AjPKpRpIZg5To80sa5R+IcTB0oZPdc/PhvV7aS+rFNon15IbVsF0C7YO4kw7k
kS8bt0bFl0q0AHlRMSz1p5kcKowKfEmIMTv0z6b3FGUCQMT3r6/YoaT9J8Oe/Ol8NE64SXz2D0gv
SodAQIkd39Wr7RkQn05lK2yG/e2oeTh8vfBYiJZLgYFcVqWML710UeCq5PfSO1DljTOSF7R5y2NL
ElJSVgpuRULc9YukeePhFe5fomfrHpbCQ33ML1NrES36HoyAkr8b9zveKCtf1H8cLQtlX6p4taHt
c7ZwdqmySvFNVRxVzuyxO5by3j41BEWmZYCKbQPyGbYgm3yhDjrEsXV+2fMzDaBBlSKvvKjbTAqL
Jk8dykwDZv9oRZTUE0OX0NSZwRWB019YHBmVukbBehmj1+n4MAQRUKu7VTtWz7zHLqFbPLC51blG
azUT5cDd/6AIor6tmkqxXAZosLBQ76gIvjlWYivLIEwQq1Y7P3l72G/17Ps4UVfVDdK3TL+35Sjk
UTbmdee7hFH41+hTUAJ4InQahPs5en382vH0pThEQLD7XHdY+efQAB1j2jyVi0c3hfu4rSA+Hy/a
BAcplskD7ej68l8DvJbEnYj1sGxW3EOIy9Lf4bBiTBtdO2AWPhcT/ecaz3lgmNjd4uTa4n2nMdbt
RWA6tqFAny/4lmFyP12jU19+g3BTI/RJMrcx0uMZwcZESZB4xdLIeZLAiT8O7SbnXf70lMgtlu/f
zjj9YOZlbkPnqJxyx/QVUtSofP4lbUl3taOLfemidYCtfPMLdC3REOQZMh41lD6YMEM2wU1WV/Ed
6pup+ytA23nporq4fL3kpkD6OOt1SUptIo69QewqT0m0ZvbED8gw6HU04psyYFjcbSAVcS/jyk6h
3gO2DT0kuuz5rwben/0QV2YYHSNEHgTbMhFHa4JZt2h7Y1Pv5iU27nt6Z2lXvmxb40nX9PZEidlQ
06LvxYEZjFfLLTonMCfFWNMP0rGr9+El6AMWIl17Hgg6Qbn5O8+XGXEV2ktmvmhmxWAU5sWH2tvc
Jo1tPym9WmZcqSGuuwGjqVH1sye370Yt+saVLJTCXkzmW1P2AovKb+Q3k5rQa3nocUq+c7vGELzk
/ddQCiGn1lM2EHzjTliWiltJBih9Y/MAuUSrOFsFZuhcwg6G7W8t1cv7fR2bJyzT34js3zKCgvda
PNt1qfWvZec4kB4tbbv6w+eX8ufuTAe7L5LQIZ9NdVpGE7VXX2XaNItz+q1Zt/loEjwZ83HWSt+m
PlBsNwXFao2xeF26ET8HaRRL952Rivy1ZOrEvptvewb9YagW5nSUc1y3p7I9sfgZy8Fa/9YUOAh9
kCaCLxeDCIYOoj+tv8GEdZ0CoAVlJ6BWWJQ//DbuYifI6Z8CmxokdnzazPQVl4kyz8ezA6Aavir/
C8j9BUH3vpdpqG5f/UnASHvdWQ2xDRi+5qTdZqeDJBtTZRxfXOv0NVLQ2X1tixaqc4PIACM+DsG9
em99LS7os5x72JILcIfICHi3lFwP54zCyL6BxQovwq3DEEoMMPzvjuzGat3pr5w1r8cf3O+EFWNf
UvGc/H+n5U3zYcxlk/Ul7FulZ/5YB02+iRnpkji0nj9heJKyAldEDq5Kr674ixirehb6EemFsK7U
dcuoCppqTtblgb47huTviKLUwfWZtpWaIjLr+13cPbkMADAcvd8XgcIX9quVyOiXRKgcW/4pnowz
1lUPcCvqS9qn1n/yg5klaFUf3ZsM+NerjxFZpNV3U46tNd0XFl3Ug3Q69TFU3no8F79Xie8Cz9Wl
RiuIE7NYnsJcMNfG+wA7QYJEB1FmTh5De7YNv4tN9TBM7RXxjfRHvvRIKES8z8amBNT4Hu+w/gRD
j153GW/frmWslje3cXeOIKMIIuAF0KmJ7GPuiMZKU5KCSze2zxdLSFqs8AhzoO/efLHPZZcNhB+r
QkaClm4GkRUjG342TuCMjQAB04RnvZ6nb1ZyS9Obp/4xtU8Zxb2K6BT9NmjCJMmBBgV37EAyCAoq
IfIwBKxC1iV5gjDESEUmASJpSuLpx+pVlRkq81wNa+0cCxlchbci95NyCnTpzb1e9g/CAXYp3VZK
mhEubWIbe8k2TUMrDmLrWm1kUsmtNPLX/4wx4JGfRi0x5mImA7mK91jORLkjUpcVgRgfNkTgcXRa
Ot4UrlDV1rxR1Pksu2zZOUTquG7BP5O7W9o+5Q3aGKabaN9E5jGec+lioYS982Ke/NpNjyunNQzA
HhOY+u5WPpmjzAWtz4BBGF2oRc5SmTP7Cu8KjB6R/4XdFSUkF9fDahEvfBpkhFLGT6xUiwEu+LZv
ExJd9t8407jnpA5uge5OiTiBJkgWPBHCHzN4n4C/G3CHqx4GRW5jbPTmLPd9TYLx2n+T4Oq6lHuc
NQ6FDWNchrPJqiJetn+aKzV+YWX1pTUap28AZKOaNwphFI4cCipvNm/DWnv4Nry2RQHfO5fNQS7n
3TdmhIpLXATlxFswbPNuOAKM1t6PQd4j0UA42zdCCasJo2CmWI+R8U6GRgd3RRRuqmf1MHEel5Bx
PFZb/TB7O4xNeZcdecILuAnbgt6mfxxJD21Xaz1xuohv4wFT+lTJJmBUAeO5Pc6WfYgPABz5Mmoq
xrz2lWeH2qDKgtvXc0HPXjUS6OzCx/6sIlc3qeMrqcn0qJSl0mxyTscaqQ0BxI8IDH/KJvwY65uE
QD9Ty5MsFi5X13E2nBTw1byGDZT8kiES4fV3/dzrzOQ53xwUq1RKv8ETBir8OLbwf/UYEhWid1sm
sUvT7nJ7LpayZInFbllu6Jj6JttW+otuLZwx+NTpBVZHRtmq+Dza+lYjWEiwzylAzM1RRIIsHaGu
QFaHkMgEvo3zfTGPwTZD+g6VWpzWx4y6kIqoxtJB/VMxgnXQWf6Wf/KT72zSdbf+KfBxB6Lhap+k
bpL+60IIGUfeTlBk1rcTRoTBdXrTFRptkkKzGJL3vJ4tY3bL8AAvaIh8Vqw/n+phIWFnTfWr7JpF
MkBJm5x/UtB53k9EMDDMuFUp4ugJonCLY3kJAmnPbVZIfI9PUKO1en9P7HkNaBluFPtQFeQuFK6x
YTgBq4pXcyW9DaaJnFbY9lZ5TuLlJzKedSnQe0W5zJiJu5WizAsmaqMsrkTsP+K6dNp0cfssAV9q
GpuRt7vtX9vr7MiN3/iep2cHl2lSSnrCU4yZUvECQi1Nx5stb7zq33rEoilxHomFSdIcrrIN2Ndk
wf4RA4EVoTodKkxDYa2TSeRU0LRrdS80KRDIZCNIs+PGLgeB/w9drzOPV2dqA9XlZyrWC79Lgnkm
kKlpoPwRlvHXpawGy9i/2RIbGC5ebsWCAZuLh4pPtEppUJbLplSOhoMqxhqxtL3oLhIMEArxFRW+
/DYhooTpatutN2cAt3O8zvAZCR3lJjYIXxUwnvxGYckvkLwivD2/DxBKrG9FDHOwE77Jw+WWjixd
lI0y9vALrNOolY9PJv1b0Y1VwD8HHRqWI/u8LiKOv98O1dVXqLY4NFcai/0IdCB20ZuN6vgsrS+A
FO0RZL49W73VCoQyp+V09gGR1tuHF76xKXSBXUO2Bh02wNMW6xC/rbRbOox5U3uXMKNXHpPIOcae
Ni/Qtpz7roKpskg0aj2631hFDF7+1+WgfauVclEncBAZKvviJxw8gVL0qypoeoCldLF6AYayG86M
oIfjwaOYZgjqIivUiRhL0gBYnJ5Y9BT+gk0kEjEfD1nKp/GR2DEv9hTfbkuH+tmF/AgFGzX7XTK7
DyM1SVdoQ6jWl+JyPnUSViom8vxHY9LUtwnaj13NK68fVUrMcT9RwLuU1ot55xYZ9GofMiwFDXxv
ir1Gs8UpzDY8eUp/mE/1oyMu4zgHyxSQqdDISVpCOyzxC05oAucis3RWvhmtCckiRVppihqni6dt
tLQ2wk1fRHb0nfcO2JIN6WugKqG/mTkD6C+R+AG6pyVOQZ555zJJnNJTtLHmcEnChsRluCRldJCt
kQLantJ46KuZ00RWhMW4UbqB5Dq6+6Sbw6kcn/Aofv/iaDf8i+qvG0xxhOYPhaGihHf8g5bnBdyb
8pYE4eiVHVY+boBAPzyqWZ2jlimAAL5GYPCbPYNyeDLs1OufOUbCOpZGJvSfG68DfVijbGTaAgb+
XdPbqmYps0qXfTPImETq6D7DKJ1E0v+/Vbf46c5qHIfL/z3UVAfKrJY5lfsfpfNQME11VPm1o88X
ZYntmrhCbyofwsOcLCalv2x+ffjuNINTyUwXH2wVWTNMMtcRHQ/E3jDH2FHADDLIUMdpu1Mdu/R8
5neg3W2o8/HpedTR1b1E94RoDmqfALedyejwNyHFyDLmyhtVAby0jmIZdgybIxI1t0qpvblQjDry
5eS2rFKVAsUE0i3Ym2ngb5FWe+EmsAeyezyrHd/lwLBD0O3ALvplyY6yZuoh/fdDZin0m2Tr+aSJ
nIlufk//HhEqcNT6Y29dUtH0LNrykdH3KB8ddpS5DwXaP+s69iqLZffZM4ns2BDdb1u4NEjEzGYF
sEYAr/iiOkXjqBzNn18/PznJ2AfdedZTNQt18nEw431Aw1TUn0lEXFsTyt3IEVtPxrwmcChO+/Ra
CmohUCqhYEbqdYrKLjGA354xdsFYHQWmAIqt90f3W06zOEwp1GzqGsI84Z+nlVG86E1YNLmYvNcV
iRZ0IrRhoHOGJa036Mp8CZ0bVPxt3jWtyGnLQsVTczvneRnRUXjTJDDWPkNu9cgmWErjFpuMK9hh
u9+9/g1D+kbEH7IywVDX0vEYIObCNT7r71mZqaibICfyi1F7Txi1Jg5vceFtA8Nvd7vqlZ9MN8Sd
TAgS7S9vKawGaTEYPSdJZB8N06luc+hyt71P5xwP7WPjPr0Ed6sV9KJAAHMgjStlxRZd2tufnoQA
UbWbGRC1WAfg4sPLrjyVekbfbI63z0mc6KixC7c7Y9lfI+MHv4azSm5NbTEMk/PmOwxHzpEER0XL
SQ1KOVGilcxaItpoPwoPyf9BSQN6fwAAYodz3Ums33WHzkUqaCZYc81d1MHfPEHJ4KcIVRFk+ex3
d+w27PD0sZDLhzzFPNDolYCxWewXeKWcsauG3Z2Gar1Q8L1fHfi2JaK2eIwoYJ34cvw3LGhhhWRU
ihKNRBFA5ZVdY2H0JmojRFL0AGhHrJDuL9/jb1k6XF+LRjkO0VRDzJP5+g6jVjO2xp/4V4US6L8J
hCFUT0ORiCYbzRZPxLhg4wmut90z3YR90gFf9G5c4guKQA7T1IQVQU6qeVOwjrwMX8HhUrsvnMam
AcYXF0159zyxzs6F7EtnqJ+JJwRZPTROzExZNkAhfbet1w8TF3dKnJmM6XU/iLzPepAxSWqFW6Kv
3OuOvAQN9GnB+mt+AUrXJ3EfGX9Pv/7McHc3VNyclo7YTpemCyZo1gKdATKtUXdiq9mVNa4RmqO9
xdIr1d3dfTSo4LDx0yqtRgnhqpGvHTyB8rOU9aIig0rr+EboRVmM7m+M37XY4tkuME+/ycy72Fzx
MoY+bcgt1RSjEcaGW1fTln5cKjIKx/mFyd/rLuFs2w0qXRX+nTuzVXnUkncQQcrDWLn/KptUAIjq
CoNJtOsYQJnKYNwejBPyu1xxFIrACpKZyt+JIX1mAW6/F46YoOCYrZAC9JuB65jRIbo4wSj2XK1K
aCoRwzusblI1Hm1V4rC/VdfGDgcpSexLVrD7qSOf1c3PwRRKPYWy+kw9XzRDoecgqf1ZaMsZbFLA
qAnfy61MOV7jwHg1nBGqG97YkTw2SJhYJuuqFHVCI+W/Ojltms1ZaaxfLPWk/f5SCwr1gKhPaE+8
KNq1oY2qyQTrYeqTAaaqxa9q/ZTmM1f8F9Eh7JUIQdz2esaIp1vaIG5b4/LYdgZ65wUoYweOiC5R
GCtf2g6Gux+4KjvXk9Ad59KZbVdCum8iEwZ8RKd1fbV8sHno5ZZtuQnYW3N1gyPP/t1J3GgaZM1C
ouRe3tRMEW7/m0n1lxfYEiz8lfc7AfBdPhBov1LI7IFgvWOEAQQE8zGj12haI2HmuyFOlCxgjDyg
PvmlnT7i8iY5OKsR+oRGUbkDVJwY+vk5rlQluMCHjJTj3e+8mdoq1TuFKyHeZGG8I9WOxuxBbsGs
xANcPjVDwJVUrRMQlX8REEBoQQ6xsvn5sHlgCt5FQgbVWocHtXgbwIXRodnLBZURN7S3CBse0p2d
Fv+rBzkzI3rh02noZAelVHSaiNFPkDX8L+lyEn2c4N9wj5kL9gy2QPyhGnqQ3zbdESxQhuTC1IvD
QDhxhrv594jmhwVohOFjQx7es4wqAjyl+mEbDDp05S5FIbvDhKQhn5ik1mFybnOam6qnMFaKGKjH
+khySD9M2h0LoHEwTmEfOrnR1nesk427cfoEXjN+GxKNqfUGrf2OH1iNODJuEpNu272lO+LQVOfz
DNNtj2DWf298sudXTFmrU1hUXC7smUNqiPuUq1O+hTyxvkXKqMyxrD7AkAdHw3N38JfRlEz8drN5
gzIsMFvC7bhKQUUKMgE4pEwQQclpkhK5rv7ln/lSoB/7IdZAMwy3+XhE8Y/yVyf4/pmrVFA+EoDv
PRSZalCRnIbhCBBELbYevGdFUV7gIPeTl/2lAmAoulsG2Mrs0/kGqqUPSK/gvG666KeZK5VarXrG
rje4VpcbjXWxEUNmAp3lua2xvTZVpUbJQdPCcVPdT8arCduxLSy0FyveEpsMz+F+6Y4T/U5Metu+
muwAbKDalh+NCPYwaJ7MXTSxEkcbU5ZKyn9tWlRQ4P47HL6n4IKDrp6vCCsJWGZbvg1B0avIj92P
0A6uuj5d9sYuHC2kBYmn1aypxLpgtNd3IPhTnb7NUui35qUHyBLsX3tKT0sJcVnIbSEWOV4THAGd
VpV/PL5tuBBqYot6pv4trcBFp2N4WZZ6EKe/OXQlCppbZrTiNNsYBty+kRy7VjCdQoqBPPSGEjh9
M9p1XhshRHOUJTwC+jajm8YIjNKed2i1mY00NThUGIu2CXbjygKsp1NM3KKTWDZuCWwk8co5lc77
fgwNI5kIjwEMpKJzcahK6JgvEXcD5c0qbvM+bLg2+GH+Qc68L3O59b3mElivG/iucONb6CsiPBmq
xW3bK9gRcpVKSzw8f1AJ1IfDxti31pU4mZCgghIWSIaOaQpSEb9Fub2Rl/oZ+QnZCxPrIIonGWoO
mfm4ahADlMLQxMcC/c/nxRMA7Xsk0lTSsfLm6Qk2VDz3vqzq0OM6f0i+hbh1A9R8qoSbO4SxlQRW
R8gGDyYyXwDEWQERxzZghx1PlkMpOAhMlECy7MBGt150K4Dz+19zyhdlZX5nIx9I4a+qSWIfvUEp
VZHh7aZ68tGOdUfi9Tfau3+s+AUoLTqjkHtma9UoIvxyi7Du6nvnSdhnubkn1efYwR1Vj+CfYFWH
qCWnQeFeQO1Ct79LDl6TaIJ3zl23cq3q8eyMStAt9VQmYmpNEt1X7Y/Vlcz9dirgRS/BLxuMkbmp
zohHiI7FVkBdk+50ayrdevxG1zmuIj1NbmP9rS/d1wy+SeZ8DCmeciYQXP4o6SR4Kl1oGV0qDGar
RwxYQQIFBmzTYJ50diPsq3yjsMBEjhvRWx5ZloaIdqSzLPMzDTLiInGQ6cc/v5gX3gq8giXBTMER
SbPmlLMh5wzCwONX5+/YOGzhGIebGQc8mdl8q1udzPPRNRUvGb+JljQh8b2hq1rDLm7roEdbNHR6
muQRMBbChoTBMhY+1Byy4LDwa0rRd4WMsu5cSG9J3FLwS+O3OscG5g7NIGKB9kFUHkADColpTEKp
S3q6zJqpowbjX9XLb28tfWps7OCi3923Lobh8X01oShIk4o1UxNDRyZv8DkdqG53GYVyIxZZ3bc/
xqegShO8gioCHAMCqJxptmlK8lbngq39scaVzlHfAoPl3dtW4BmLBjL7lNkOrDILnPTQnUXzc4hH
pXAgaKTxewjXQpn3dGhwoiXLXAc2lmokHgQqu+4wa39TR5NsAXvmkYF5T8nv264r2B6k5iMRIlFX
hbRzAbdZNFcSNjVWk0zpwJBcg50hLBVAHhzhGMRl7gVoGsKqLuipks/Cnfn+O2DY1vTedekNnauy
2XEF7wEiAAhXEhWI6Soh0ZjXydqintpUOvdL5e7jMC2C0VD0V1vC5wvBkdLurje6rPQ+au8OzVDD
N4qjZ3+ivSoLs3QgdPu3BbZaZSSV54hEgsa8AfbUSGUFlFFg5BAxQmkO4jL1F2GAUg/N2uYh4Oh3
rt6/rW/4sjXHGMACqied8sepn3b/AL/j/igeQBa30OaJA2iYjOX6WlgoIMZLwWsuCFooi/UpkZ+7
+V2XsDJLgzjLfuEz9cPNl3flt8KkTT/lLAKKqjqmklNUuOFs+Q7/LPVKTXYEW9Xoua7dwjwgi+RN
UI4VcDdy0Ig94vh3xc4gi/q699ZLpIsEEpvcFJT0WVDBNHJmpxXFvPISTAobTRdDhuFFa+/791ii
THQawqs/8hmw5AMFT5610Tv5ZGPj7+LSeZu5NPKiO6rwmOusz2dYCXpayKiE6U363fQA+E3YYqng
+8mQC2gOIT/edHiWoq8eMi6ecphp6klbIiimwUz8BCAk39snmPtCGYGnKBPpmzB0yKXM1D85ciOQ
tYi4dmN8ekSb9T37M9fcDNqfibP31QRyLIDWGmhZQ24yDGSreC0RMNAdakhUpieOKKV5Y45Nc2yr
wSsmxCQQkg0mXUfpG1c9yuuj7nmsfi5llMLGuwcBU5NcczeyqS2aUm1Oept29gzox6oW80GJUgI7
5rYdln3y93OUO3nqWR3ZWVaM9a8u7NkRWnZpbvzhCaysrbJ82v0W1Wl9m+E3fARLLmEVUHYrOygR
uVTQTpvsC3zWj2w4SBETP4Je3+kAoF7tA23kb479pwyLUhgKWdrpYYXH4DsMi1f2XAcJOtohfzUn
K3P9OGi82jGuTX3mKLFhI4aQvBhWa+p2u/zHCgyry+IpqziYA9K4TNiBWVDClX9FP4j3X05SWnRJ
AE4cCtxR7Ejnd9U2vZPBaEMAQGQslVkfeNcpcyHpS8PLwItLDqeVY0m5SvaRnrVLMwFQ3j3Yh41X
/G2LPzJNobTLPRA3OtdgtxzWfOuGihkN8NSQzxkF15XMc9aAxZMOBeb/x5w1D5sBhCjbMTC4ZDsS
bpxpVqxdc95xZGTpkke3kSTGRpHCKPUepOx3rnSEvZLzaR8OwIHqpAT7Pqqs4eWjQFNks808jXA9
Rmoi8/or+2KHjMmRJ7rJBvLcvcy2elfBo783OJYmIexJKjch/+RwmHW2/ydLoeLFS/yY6YEPhjRb
M92DQSoIuiDh0c9Dyu92/fgjva/nxkJ+U9P4iWbkTX+QRdlkZGsSpLf2Q77yAzrASa1nDL0KnrJH
+J27MtCaL5Sm9FxIt0tdhaRiM2GICmfQgJGs7dNY4ZDngXOvaht+tfp6DggcUWU61bSJG4ll0rD+
/EmhnTmxOsrbhvteCJkxrLwGmECcx9dHTw2aHhmTkj7B6gPOvKX9D9kViAwPxxTDLEZPNSmc3UX6
lOQ/A2JttOmbpR5AnpPSA+6AfZ9HdDziTH6XBP39z1zHWFxgho6eY9TvqpiyjXlaZrdTecL7G0wr
cU90Pz4PndPJarYT3fa/FmyX8OQHp7SBlvmGMksHjzxHuOSBk+2wEPi7cCDezC8LLCHZItQm2R69
riY5YSWtTlqdlh1PqP2YMEG+plSD6/yl+bw3nQNzeiwcWj2GCBNAPj+io5YLimIADpVkNqnSC32V
dQtkVtDUaeF6tvNeumisxrk8AssyqZH6rgnJ2rCCcMu9TA7koWEaNFKDg7g9fSX9Lqfzx7xDhbfo
xzatKo9H36zyKoFqn9kB0MFWkrsBhM+ukmIrq4MuX6sdSTVD52skND7A/pCRZqmSqpAYDRpiwaXz
yoni/XkkLPKQHJT+R19AGAQxipHFo5ziCzP9xPCXxxIIfYiywxqNO39Bb8EfZCDn/Sd0c9wlGYij
aquV7F61XkvFYsRkxN8sKctfc31VJER3BrnpQ7ZSSWRSqhMWm972wV9nOWnCgJuFS7D4QSeSbySK
SOKBZ4QHMN2VMvZlX6/g/uDDvYgfDXrHValkX9azwJUtnzge5cBzW6FpbHUqEh1ikY8axIril+tK
Y9EysP0hHLZEnj0B/QrsxjvR3Lo6V1KodGY+2iagRgnW7kWOujbTKqlMsISTYXhw1P9KJKITeyAK
GHPPovlqzbNtVx1AHqRsQibD1LtOo4d/tDAf9lA9vACIt36bJplChBV8bIUj5xoGoVdRWsDF3tn/
iEvFS9whtPFSBfYcRdfnXRS+ltjBYprDwwWKfwkXejeRwigUs98b3MthlWtUXj+x3YMSr2Q5Lsr4
gfZ94QQKTcafW0V6FnMWVFrKwChk2QDLMBE44+GY2OJv9xQz6VCStKtO8xmA8FyjFC3Qzh90LVC8
jQD+wIZny5ilcUczM4wMcevGtx1x52yPINGAXncnEbhL7VWdNI1XyYWKcCVEtXZhAXChFWkFUYcS
zWHWE7ASwLtoNq2fSfuZB9BwYParyvkeBpxmTeKgImQz8hzh1F75znIFn2IE00K1s0Gmw65WFQCz
DdInmmddYWg3QJISj1zy7P+UQzXqqumvifdnTA5L3OjHUOfXApHGRcAmp04ufSzQi381XODJ30+y
oRi5iC3+evljZiGwedPrtWt65gBELATrx5B11hHomygQg47UFEpvdUkE2vBPHvAj9xB6T92/d2pL
kGSsm22H8AedfOEsH8UXlyGDjuEU9dKtXpVZbHzUen1cozaumoinV8eF34iHWN8Wr+NbYa9SY31r
QpXp4eIFK0FfGFlPC8HncyYgka8qDTWC2HkADmGV53ZzI4RiXCRCtqc+qyt5y02h2dPEdVZxAEG0
BoHc2okjiLZa1vrF+lPbAxq4SKbKq63EEcv67B+8zDPBi5UBRzJwOHkVefV4Sn0CH7tHF6P8oPLb
roF+LUa9Rd4Dzq9U5STRsP3q59rqnM/CjiUBL0mtubUlXuSm2M1Uh8AEYftT++CumomLFkherYrD
hkFofRhkUsdRcY4aB3AmWG5scfPOpvr2W7XSVL5Sg2jyH+jTLPMKbuduyBB/yffgixttmU7Yx0o1
GuPb1zVFF2aSsHw83gJZek4e/HhlpzBhDiWxsu10sCz3kE3UffbU9NgewxpShuY2E1F2SNgAquhU
JJIXFIL4NzD4+YSnZsW6kZ3zZQ1ErdQ65jchk75R/zBrn10gY49Rz7eH0UUHBeCWdrCsuG0xrhJR
Fcrit+z6BODQufsCDPJxjsCtt0Nihcg1XcCEujUhUlLDSu7EdE+Njx3RXX+sX//TkT7FWnumNzZC
wSURTlukI632O5LXNqrnx3VoLu8QEPTj0RH/Jm1LP6YKsfk4Qluxt8YreNsEoS+Gk8OJ48Fh1GqP
iQ6e1a6xrZmAKBL9564jzT7Z5i8PLkcfXkNgatp80UT2W1MLyfm46PDAj7iLv225V2akeEFn8h7F
zQxml+gZftwmj9B92euWYFj+EB7nh4sKcGnfVde/ru8MdcMuE4Qmh+c1pHEL4vBktd9RuqXERChX
jcHuu5KGUJToMR2w7tv3gEs7I7uRgVvG97RbbWUX1yQVpdTgy+/eIm8G6OhLm4DrAT0Mgl38wWXV
F/KtuiZnZkhKWcfogPcRhlLA1lA3t1rJz+tCiMe9g0p2Q60oCXM9axwF0RjOOtCO7PwemODBf/Rm
DVGryATrFtB5SGutPgB8vk25kePXwVG7fMvdzYhL7NOiUaX/BOCBCxVbYfbZZDwrvfyagHRla4pN
dkCRDQl3ylihBk/5xn+xZEhYrC7JkOxt7+nrPE1HBs9a+ocJ5Ummf3uo3WvWbi6LBmuxuynoYJSg
ZtxWNEOfYP2MkjE3hzUKj5wus1DOqVl15hQ6AUnnPey6SleLX+5uTeaN2H10ZuQWi1Z+IR/609af
a71j3ITgLZQVbw6/sfuZY/Pv2EngXXwxS4ytNDm6XLwNbM1hWr6aQVX+Czba1LO7xm13c7G6WoMr
BXHvyRiPpd84TjuP55Npj3nKquNAXbmndQ+rYMWI0Lt5/Dh5StUAlIMcdBA6i8aNmXKbTSUMB3f8
JrkC5UFUpdGOt0+pHPMZIWkGDxLyyJGqeGimEayXZk/kG44+rwPcgCYU5s7Di1Fl+3xtGKAVf2sD
qxoJ7lSN3/6HSZjh1iBhgh+BtZ/8eagDBJOLie7UqwXzS9325iJuezh1axgvWDzKlSp1KovaC1IR
EBPKsJVQScyllpukUtlj35mzTlqTt/ZTl/C5dhjr9KyQ6Cfnk6G43+VE5/MD/REWFx8RgAxpwC9c
4zXVr+rbBAFVDlNnKGdHiv8KwnwC3+D9yPYUVdYTM7UDbcjURNJZNM7ow4DslGAgOjjPRFWNdGo+
Sg1qYrpvJvkWXU1cb3vUO52jgdKg+4rwbNwgtc5ZGk9Puf+GqAxWz7QEyjxzmU4lfR5cn5HdNVO4
SE7Wi0Dsx+S99RhTHeq/JyqavpsXe4izhwi+jiE1fmxP7GjH2HI5Y9JgN6WiZ4y4aUUUOy7ympDM
5uP4rlv6qzHGMUJy524n7YOEWKqdaJQLUbl5yM/HidXamZANUuB/Vvv/WpEVcFC+XZUhJrFXlU0/
Gw9soqpB61vTTtol3kQoriZ/hb7uwFM88LrAFqaxz86sTNcaWWAieSmlhbzLDHSOSsEmEpFPZN4Z
adx9vHieB985RjSY02fei/fDQo7HP93ESwv6ha4jajbap16n2cDlZEHW7UBQI9dL7ggMFt0LvnRF
L+VW8PVmFgaW1anizBQZWY1+t8Xl1WqbotES7sY/8H5v4Xb6Ze5FcanFqtDBdS3IHAhus2e4WEyE
bNdWO+D2LyvJZ63CdjGiy4M3ryyjE5d1g2f2tj80fQ8pxAnVZOv7Q/bm6qY4xdlcMlScc/d1zMTy
n8R9MOr+PjoxPAfu40TiRoEkbJCO0xSrFISeGrXCDrpqP10LTZKHG9NKjOYXhHto0y3aZHwP6COm
qFsx7bZ2Z5ZS56dPfwD2hh/ctqwD8j/jxuOFDsBmfUs3jCMiD3PgtC9C/NltIbIVbJsjqfTOZBpC
+9xuHvocnAFxGmd80PIGfc2fY7Cnqy8wD/o2FOjNCyYnF5izX5LJaYDN5yEGopOxynvii1+mhbVf
jdOWb1/frqmx7aek8+4taHZi/ulJXheHVQ9n5WNjh0Uae6bNRj/6ilZ1LIRvsYeMO83XxnhE0nLf
fSk5S6BFZ9bpgj3kYCK6a7jlywAoqPvFxaOCdqWFgHkG5HGA5d9mGgAd1UsxKA1A0QvR+GcQADOT
E8o6XLdV8Aa4puQzl/0vKjw5OPsZNHIdLSC1IPKr49dL2n9VKKGRRW7400Vmy50mGVCGTTm+5Wju
BoE6BqjdRySiMPPHrF32WOrjnJAfwFsv1Fb8GPm7loyXZ0l+DNiSnxNVpNE0yS00F7OA9xiGrCls
f0Ubbc2TpjJtmPJAVPI0MYK43uKX09Ts+X/y5//hN2SrW+Ow9dSNsKAoZ/eOLS0BGgQzG3o77bqA
vZKVQSgifm9AE70wSfy1mjpFmg5lXQK3UTrdUfrcmNZxPM9HChpK8TZqf+Lqkp6mcsb1qvFj/Knf
Ct7aIQW+Jab7PuY6+l8mQcsjRSfjK0zX4lOL9/IIEuhVd7qQ4214A34kicHWcblWvR1yT7tSxCcI
K0imCsy3gG4eYH3nySdhUy7XrT9cE4sR5YQddUenLSAOw/ZAgDADEXYC1Jx1q46kX2YUDFy2kYeb
YmtQwHpvb77q++Y8WN7p1LMp+GWu+jNXKNARiDzaEusFJEg8xHVmKMpIC796Y43UT2sAoxMl9VYq
khO3QRyqKM0IY9687B13h7FA3plCYLinxFgrSOM4oAjdldlB4bJWvR6VMNSaM7XQOxcMh1uqL1eS
kQ2lnpMVdh0bNxPXBUFbymg1AZR3hfbfrFTaHT//8titU6UxQKzR0SNIU58+A7pcIDmAhw46hEMP
wzeqRBJDFNNJdAUzxXcQ+tOgH5XLOKPeLgkc+k7ndN+WAYQWGCemxSE3OyfvQkck3FsnlkeSCMaL
rN/X71d2zDLzv9Lms92wibP/GagE2wPYWFVhBTCdYAPcyJ6Z47KG7/1pKEs3ne6VwM/ggNkcMiN2
UZTbHRNFG9RvDMxWijthdPKEj8afWKOD+Q2uOSECl/38mr01azYxTWflPw+N0JP9UU9Xx8o4TF6j
gErRgE55GxWlR8PRGim314iQHorcQecLPQN3GHjSeXnE+gaKSDnrE2INj6tpjiSKkbHZuE+IzNxn
Lvc2uv0qqhfbVIBsfUAiihjPhhGTFRnmx1f8gG6Ydio35mQ3d+mkeZQvAusxTcMBWlVDpzob08/j
H09LedlVPpvtipAGT5T63FYJCgcqCm3SLuxhpSwtW1sobw4dA/CEyVswK86ZpICKipr3cZaudVH5
CiAyhXOMD50paWJ4+BBVrebr8NieMfQCp4Ey6hE2rmSUh4LYsMJvuwOOaIaBsu+6B19ZQAb61Z2J
CIJtwVrazPBJN9eQ51uSD7aaK6REjPIu1D+WxCfjjFkANf2ImsuuXys6ngVu2X8k2onTYENVdX8F
Nw+vkT9GhtXlXIWrBnAYpU6KH5t3JthIe548p3PTfpUBySlnwUiVaytvp9RNTqVIbL/BCF1e5nlM
Cj3y9FBUFNRBSsyYQJm/Qyc4qlXkYLmDRCV7lKx7VbFE6x33Z8xlI4+EwyP3iB0B5f77WVAgF8qE
8p4a23Eb4pQlVUGC34RQP3KNguOiLzy9Ser+yg/BcMq0uA3/ZejkVHyJwNDA/vIFpTayyKtJGupf
QD5IaRMc7E81gmrnLfie2iyBw7y0n+Jeb3mVGpDG8f2/Mu5EomMMmKcLoznU15Z70ziJcXlvD7jh
8siDlcEL0hn8YHnreGSDmf+sgdhgEXIPWK33C8YSuHvHVMudWmD2l4rYk2NTMuikD8HLbR6sQlq8
8++UBIjCXbFaPCFz8XZDoOp52zcO5t4t3C5g6nzG+5GBjY5XEkUMv+2nvnmnO+qXbza2ROBlzLbe
XaL0Rp0qTNzenx+PgTPQRL0RJeI/ZCCYZ/3KKF7X8SfM66wmI0QhxrzLEnST6MH7dHQnJP7RjhqZ
D4zjYU9WD7KpopkDLvM6HyyVLbtXSQlsF/cQJD+fD8jpEY/P9Vv8txpzN/cMpZXePlJR0oJ4q3WU
MLnuWTAw/LR9kU209OCR8OMtxwJ0vwgmHdHLHCaHRHP5ixtlm7cf6FyVFiCp9A/o7PAsnXKIkSLo
rasU7vut8rJh6OGpIzJDhOiIZc1JFcHg3RsxotrdbFRD/bLZD0Z8XSgxdKy9+Xwy/2VsN0NVARfG
6BDfgHU987v+nYNzwI7J2PQ9tUTd0TcDvqmJPiA79PgU2X86lG8ecI925Y615r88V6I3l8GjP7nA
jpgub2VzFELo+Wdzq7T+ioVFPqNwGYSIOD5r9CzAUe1ZaaXM0/7nvgzzTcMwRURzM3D3q382qAD8
W/IFn8gxyNbo5jSV6p6HyK1VrVNmphTiEj1MkmYAqHG/AaLrrnFWvCtdRtEafDBqHz6h6FjNFUDb
5mtDDrTgrCyHof28NSCp/2UYWehvn1vLA4hDkO4PONyFWf96vjgvcUEc2Q5LUzxIbGjvKrULSvXz
Vi3vfMm5dj4RHs+4I8aiK9ZfHbh1ePcFTAZ3Y7zNR1QR41Ztlyi/PzZxZXjdBzBgbR+uxvZmnVHz
AsB3JQpPEpTz6X6KqSLuc7Ery+x+3aI6N22EI9gdLIKpEWpo5tcfIni7oMlmYsLHqUG2qmykYqPX
hHmMz0xYJVgPDW4cF23QTFGzIUe2Km2WldgOftVwAx+TxW6EFCzevTwZwmoFKdjj9r6QVEN4Ml19
RsQ96UTSXly00//TWC6NyCc2J/BDO9aRfR8pCpaQXIlB6YTe69dUck2pjcxFLW5gpHdrZtaKlOYN
A6mW3rcCBDnmpFo3kc3GsuWz3sdFZDRdGRADyw6ppC7PPDOVAIfvOk1l9K+AoWtbNQy9SBsU8lfL
or96d0/Xus6d/6HroPcAfMy8fVpj4d9IM+wCGt8VrjfPQkpjsYtyz87uRUzgIeqyZok+93mJ3hMi
7DeR8JtGP6rsUBTw6GO2XQn8jOXKaGPPiZel3lysU5ZcX142sBIxA7AHrXPtooqvyks+NJ70nslA
isc+20IuH5ZDkmDu6MoGgeuccPpVo1/jm3fJbyMhC4OEXQO6SkntUJB+N2XEuEe41ZanzPLVBPXS
xSuMUmJrpJCCCj1LqK9kQyteXZir/Rnox9Mx38MLxyE1IMaI+zLFCuyruzdbRv0t96RWqbuPprPA
LWQy8e3tLM5tJ1iOKhrIzyi8kPlus9z37QQntQG3HiwHDFx4KqxkexMULqQR4IDuaexccKD4c17e
xnrQKL5PvlyYha1foEf4KsS489K0YG6TOGpMU/ZBrh4pxaM1ave1HY+M6+yG+eqne/4zER4eQWnA
LzfC4DhkXYldxQfiKnDhGzgMNSoQxZRN2fdXNzKVhNW6qG8RWhlu8qLbn2lOqkBhKKpAxyNURPQm
uKIB/OPWQXtr6MhKHPeVQxDDlkgG+LKBCl2ZIMx38d9aA+3rCOqHAicqV62u0wIX43HgkXaz85TY
flUVe4EQQAcGDIeLVK9FMWHe8EaXLFwMSuNTS9xR0ZY7Uq2qetKTwWURMOtGvrQ3g0QSFfACxlSz
CRD8wvyHO/Do7WoX9Wg04pWPY8Y9ZehEkDMdTnHGWWeeWutfsYmAKOXoRGzjhzNyMvjWfB3YrvE4
yHhju7SrIgS3ZwLYK3ywYhuyszKmxpc95HkcieXMtBRWa3g7hzIvq/abk8MmNgau4Nof/iFg2muC
abpEZKuTodFis05dwTs5/pWTr/40ddD2/Bv9lvITRSK7L91X1AZOwJesVTHOxxSGZEwjGbvfuMXk
pD1JHhnk/YoeH4F2sZx51WpsDtafhAuylKirBaKquTeKu+FhDURB2l9CtKqWMuoF6n4lie1uMqIU
TmMiNmYycBaYBaSO2gL2i+N1/n1HnRwmc+eNgb653RiCbvTp4JJqz/S5ZzkJkQvbzaGyqByqQ+/3
ydQv6PDaq55PTYjvWAgRIsm3em4E3Opt2JIj1Jtrq5x1Xm5GhX19JmlLfZ4NZarllz0AgpAT8rsG
V61xzIGXOHe4GyyR+MeAsTsDgPCx7bUJlupXw6lZVZ/u4BZRfEQEVXaqvTU1lIjz5iNg7ami+jtQ
5BKYwa/Xv/Nl4UruZV/EcNQr+TAIjwigUec87IhW6UpQq9Cgxnk1gWtS/cX6V73oGJG9/wEX6TSC
1wvbcGfXJG/I9zSP9kUnro86F+6fRfUx7dXI3NmOSwiDnUNFJqJXUJoXLAyoNm1qlhMyhzO1aj67
E2Y/52TxCBOKvwnwIHV0zwqllcOFgDpLmJBBZ0UoFl5fxWbDUQcnuIE+V+VhHds43QQvvNFAA4WH
rTKgfwj/Qp+arZT06tXtn5zHN3/jkT4wmX57haXlkpQF97k0YHlHAbh5S3FJ7MKsl6N2ziYXGNeu
E/xZKErdk4f0H5gNiEPXYEBnBkuvIoxKR++AjukC0uitlEqmyLkDxZftyrE7q5ddZ8pOfwRkXMB/
fPiUQzkyp9zOMTH0+PniPlXKeUA7OlTeO9HbroviubAePUgxv5ktZUtQsM9moPIk7o2rBua3bXBD
Cp+fn0XbD7c8U/FHXQCo/DBecv6Qmi2cgHuwfkvSkM7NyzJ4FxPpqbS6Z/IkeHJ5EP9rJR/4t4WM
bAIisCNwYn43tISwPRid835WTOW3vGANsd1JxnMNGx9rmub3Hg4vdbDgsE8INodav3Ltc15pGKw/
FHtYbDv5rUQbqInq58vDDLC0wIBwuwrqGe4vpBLKfMvSPpdT6H6o1V/nMfB6FloV1g5ii3Pquh9t
oiP2y0OS1vO9titnBpo5xY2yeYGg7enr0XDGPQqG8tHDLmyJhS05xOGVoumI/zlwwsZ+KLyG4Gz5
n5++IRLviSAYArcIaHWQWh2QLjwIqzcKz0Teqg4D/80qhIoCB4yYUhWH+RC9mWYHG+Nk5+Kvl+EA
LYNp7pwhOlBwTE5OOmQImqBoHBb/1k6mGc4TfEnDtNng/rr0w6c/B/s2BuT2POPeAdAf/JoTxzUh
nlURizRgArS06AmeUUB6+ZdGp5p6w8rrpinviPUVm3B9ZygtH6kGqNTg8y7olMXYwgi5t12uIkxS
S5UsKYDhsHVuafYr3YZk0tv2DCw077YqRWJklIfiMtMw6saGIZyws6DUu4aLOIJ33RNL//4O9R1G
hV4JBGeaG+i8MYjaVx5Lt0SV6vDudyjAdBjCRxEuBT/ULErrEvMcprwycas16FE07/TYWa8Iros7
n9PCLvB2xMQdjmFJhygP98Hlx+C20Qx4UZD/MDRtgtZ/Uz29YojSXEm7kRbX1t2ZVHIDH2eK91Sr
a9Dyi0tO1Tef09MnzS9ESzlTGpkRBYou4CQxBLe7Dv3lqLdvcmiwaJmaAsC4wZYd9hlLcMgz7O5T
t9HVZQMAPp38y1jMaCXKhPICd8Iug6Vh+l5ZyTBhASSR1g5TfWiluhhhGBrOeorYHCwI2bc5g4CU
QOi+MNGeqmKzqxz4OzChQgkN/h6vKWroKRjx+toyMUXfA5oKPVyjRDoK+B0e90eJb7lAcacWvm/B
etASQ6b+5WSOv3zpsetmnHS3UjT0jQEdLcDvXNZ1ephyo3NRbzHryNgjr7qOqq9SbEnVSFXH3UPU
P36fjrSh9t+mvc4MgRYxqsM1DB3VA1VlTuUCjVqM1NyFLWxZSlagC/ap8I/t0trfdvHKWkpXvL63
5kJa0V//twYAwwmLufTGZtScf7xlrlQEKJ4h7ITzwtdRw2Ye53aqz3O3bHwupAW2O6UdsJPJDUvL
/5HwZrrXsUFMJ9ddmVJyhRxbNzCXTZuIxMtizejDcVw8Pr2k970hyH8A1xp2I97o170GqI3QGOoT
YtQhKbM+fk+bjWrZWxRDoR+NfLzXWSQxMyGoDP7nbXWr4svGU7T+SxEOXcLZty3TBGSTrscuyYbu
7DLFrepuYGNHtaZYhe1uwqAT3TUNyq3qO9zJYZ9ff2AqbQWll5k/KalMfJXWAGBNLr8LuK7zm6Q5
7FJ7ikmK47dlVONKVtN2qprrUrqzpLCPpjFjozWF7cZu97UxNqWWSea0xAsoSWyEAmVpT1HdnjV+
Acf6SWRg7OoDcbEpc2x3811kXfdVTKKuWy3Xepa+ZeyX5qdajPZI0gfGndBBfAotGNr/WhspbSoS
7+YDVRpvHANoskDFmyalFSmAaarsuy4aDws8YB41elnkYlL5T+lOFm0/XCdioG78E0M9R9MPRb+6
loAq9faWcTvyaAFRIvEMg9V8eR6ej5Y+1IQYbeItBn70fznXR3XyKbDyeIc8HnPjYv60xiaAhiNJ
/jF6zWsGf4b99JTeNQmWDCikhiobGWse5Ff4LSTbXvk40K3IKQ0Is1ff+VLfkbfyi00Ra+7LHH4y
tMDAQ2JtJrZ7sONNgFQPEBSCJ9mobUCwcWRvUdqaC9DVORJx9PZ4dq/so7b9/cAl5v2153u+LoJK
51MDFVSRPKsWV9Xg4476lgC7tnVNAHt2OZG/mpX3Cb0m+PkQqXl2yLAqz+Btbqq/gAK9AnaMRvJI
xXWsbT22ipiBBW4bVSCO6ryq032x91RJ7D5vNiG9nic9V/K/1oek97HMld+9ZkDWJYV+L7pTmlWa
MhED+0xhSIUet62jPs6GsN12KE7s+PHIDDqd7Yhi8LULu73vevgjgR34MnffLAHzVeZLpVeuKHD+
Hc5CTYBDBnfW9jibLwaVthMgu55ZXqOyGDq8WRBq6ZYxzCTOg4yvuIxpurlUO0AMDe+T86nYb7LW
CEevm47575sZP8nKX9wWGy6T6qzAiA1/GvvBE0grVFc52GvoGQUv47MbVOL/ysW7gl/tUonTWs3q
bxzwSKb/oaIVSNHRkQqUNTSTpU4Kg3MIjzQRBD5suc69xSeDx2f2nfAX98p0IodaxsjuG0XQvLhS
wT2MCIQe82jXM/z8xeA3oeRpPyI9sNRcm85zaETtGyWPgNfQOg+HCrhVVWxuO/dnRsT1EByw/l/r
GtSsW3+hIr2x2BVnRQxxA3vt25VL2Esynl9jPdozO0x6gIzkWtTBreyxREFhI6rJt8le4Otxd5ac
XW8umk6G+VT5K1z8bZqdfhC3ih37A4LnNQ5sZrPVzgNRt+0x4213eBQ9O1BTpy+cRD6k7Khz5Fdl
wkhMwJbCavJ6/Cv4UwCeTr/7QJUYreEiBlbxlcVm90viX/Rlj7985YJFPPASBa78IPwudk9LWHq3
S6V8+29suEkuHXgkTw52bXnI9o8QpHq5xDY5zRD+slMBfNgS0ShvieCTq5B9KdWczsHUV907G44S
Wx+oyu2vF0ep+maONM0SeJ7KG18VcnX76jXAqG1RKT8KnGL/wZjixB8jAht3DBV5i65dHSNpmOcK
s8xrP3jOCyL3Ng+GW0sllL/6dv9+JHObx5lNnncOuJkwuEBuk1DC4xwq4rWPg1AemFOUJ4Iw0XmJ
wliHRXpomAg6+yjZaL1m3E5Hy5Z2HFNRFTc6L2L1hzcCpyfIWK3OyIFeuy7wUa+p2z7I8I9WO6bj
2mh2r3YTKok6BpPOy6oUcdyEQfUYVmtMPQgosIUiAZ4jfqZj1HaJLLbNhewSRfjZdKhCpKBmSvNZ
nCXkrTOxh3qv2gl/KoTUMJEmF9PCqd4BCigJxKXhMOgmm1FpksD2njEhlaIgMe6I02nYxUTyi+J0
PKEgUfPGcadm6vxXmKogYUgnY5c3nv5DxUP90e0QZ8tAAyUrW3R0dRsdxQP6d0wwZO5HPNHtgLE8
5P66dSZ1Su0A+UIQLgvGxTg3K2t5aeyVxQnziPFwEyWKFVHyu1J1OHIgMM5N4PTMwfJOK4Zulzsl
zMCN9qjt/I1xs37aAEZ7gr8jsmRzqDARRFLBIqVrQSOSb0yUE2t3RB4y9eSnyK1SdbGuPbQdrud8
nRqVdg942eu1iZOnBgthyQV0cWrniZ0YD/RUkIEgaPeXeDQc5exk78PWPu/mj+JaIR5jm7b/KENj
NDv/cL+dhvYLl6Evuzm5SWwA09Szv+EN352Jzff/NmCeDXTqXO7qQREmF6WN5IJPhJC1SYXvuw69
MbZu1Hiuae8jmWali0XaVeYrc4Jy7wAso6byyNZC4tWuxDa4/tYa+Pykwzotl/4gCIpa8KHme06a
dXrlW65WudEIr015C3pluU4AOATCjZK6IZrJGxJcdY8eIx5SGxrUmfuG+JkWYlsJ7oF+oxfrimaW
lpXCGc3X0FJuE0K0kjGZK39WwKJkADBYrV3TuETF5Gl4c3ydDiP3MQU4ESKinIn+evUOvQcMeePO
geR9oC43y43qV0oGmfY1STdNo3+SxNaQOES21rMTRVPocgUvTRDtcVGjLK47ZRW6zG+/Bs+i+wuM
JMRyIk/MIJzln7TEEuNMgM/toN1JUGRSTCHO9RMNPzeJHcQfKiSkk2tDVOkWC+jRCRwfnCe9zjW7
cc3cdybBuuhXdoxZrLhxqkxhNBNKAYINKF0muQYXgdpoQuDZ68LBpTppVZ+ZjKBPToSlEYf2g8hI
3sfLkht7tXbMJQrYLEhbcI6zhgbax0Eata9QP5qrrgc6u/+TbiqscipoVTV+lP12fGWcirSdq0DM
dMk4aH8TzArQ6QMKz04UGF37E2TAs1MW7fIVNj1LcqqJu2RGwedQpy16mpfeF54BKjXXZpz9C9B4
e8ljgxHTHAg7pNt1x+8eXfyh4aeg368bRotyv6sWKKuSkU2ugq229YJGjMoreUVyPeeKciHGPmMo
McsF2R/M21oIDY4EKTY64vWfFuV1aZVN42Drut5dRwq7uPJJrA2kYFZYlUfPaLaMvJMxDgB4OYkJ
+Erq+6BczMXx70ZKYccTYrOQJYYyTqP75Jyj3cvVz9MYeCCWizjpzU6K7fESszHjtfr2tpDdCc3P
uE8Tz5Ij++vanD5SjdjsFDGqQn2eEAacUJ6a9dA2d9E4juE3ay+C9BArpyqWjhzkEvgXnNLbqeVx
wsGkU+3vDD6o5L+EzN836F+ZxOlde8e/+6cC3NBQN3Ge/34erxRtn0Xh40LNvB2MZD9uYsRJ/6Pc
HM0XZ0EclzkPaFmcww7vQwQIaGra2DqM89W7jiIMNdVPEPu3Mky/3DtPaBnuMN1Pj1xf1WugJ54T
w/JDU4UntYXjCsd0C75NyRRoOHLacGSE2hB/vSvBJKjfCd4L03I6Yv1nXTo7w5XkyC6aH7iAzxQA
F1eCxBhQC+MmpZQcciVX5IIZcKpuhaO/sosScdFW857pi2HcmjJz85VNkrB618axallpeoMKd5M9
r49MzcAYAAtpDRFmeCkoxa2tnpKIE7ekTzqpzm5YNejKL7aEIPO9YKtGLyjLi5J8fXB3rz8d3Ybr
iHH7Px0cbza+kqgb9tfC8K+HEbROUSN4GpddR1jSZFy7nzdQtTZje1pOGlRgTernIRHw+FGHASC3
KB1lpLrhzRy58zVY/KBoCeuYB3e4GOe8qXd0MZWDi1Dx14LBI7gRDZCHdFv9rjNf3hlRbaiA53oJ
gzbKUnXr/OYfTlOGKXA2jvgtGV6Kenf0qF1SjUtOQhb1g7uAc9bBBggQdw1oPnH6hRRyyMgt6SxX
7CHadWbem01JTuLQHbqr4PGWps4u2T8/J7rowDzaHW19cqnOWGsfprHF0jDbAB8EDpZqUXlXA87n
oVyso2sovC9pbNDEAYRuudbI8JC0+FRdA9pmVzf31jUcrMPm83o8pz2D24CJB6dYYbCVoY31bQpO
sbQw7fgu68MTvIUV0XRyOaVShKW44/IoRjVOqYzGFUF7uPbwihP4dXJtMF6ZMsUhUp7EnT9cca6e
1vcq2fD+KLl/OK4l2bzD0IZgRKfFRW7RnBmY41veSUbK0Pi5uiKoBuh9XtNdw5ySxJNeBlqFhwH1
GCq5Omp+cvHo5xy8RZqT2qrxbleISKW8QKs8R/Maayw0iY94jWFan4FJ7uhgdylx/Tc8kLfznOIo
0lWG4NnNoGv7tM70i26eBbxAkEFn3ZHVaF2eW6/2uFmklN6IMUoNOjyYuQk/MeQBgbsMmEGGrao+
WTeHHj/jJNEqbdCWkvSoGFi1/9xORchI5Hiczx8m2K4mA8tSnNY/h15HYM3Ey2zQTFZD/pJHYohK
xOKgQ0W8OGDWvCDLOfm1NlJ495zCQkptBEXfFZj58gKImHCIzHkzFaZtA8pWZ6zCDs7hKx8MHM0a
XJtdomOq2a9SADPDnmwT24MiscJhP31wASSsnvolYcs526ZAC6U/uzi4K4lApT5tq8FhArh8y6hP
LDvFqR7FyQvC39C0KMjpDA1frv539mGQTAYGzLKfkFbBgeED+8mnfluMXVsgz4QxNj9ODrY3qSg5
Nt6vXFuh1BlIhjcS45zMv6/015TJHqTFSWvfBl+4YIdzdmwIj7QruEFTPfmlP8tShmnPtetC4SDM
N/ZrymNMxk8lkUjj9JGTIfpGToxOryyaZiKN15U4gwOZC0r8THKu0pHXz60jBstIvXHsam1y9/k7
Wg6cWdgDeceoeYWbBwG6QcfU3vVJDkZ5/+W2JDWCAwLUyrTpjkiP+XK0TMQccCixNnwB6CEYNi11
CClBdmMo4TrDUlrn0CsUHonanF+2PtOBV8JlW2A6Lpi7B0TtAo0TyVVlDRDBONQGDHWBndpmS6nX
eXsxSaFtOMKZX22e2ZUhOtoRevaUZDeTmsu0iGVoT1hMVb9yJaxO2IW2LvRAn6jmc+ArIVsHrzCz
pV9rMMt/Tu90/yNwpU5DQZyQzqku3kwCC0T83vlZPoKTkeRss4OHaBwWf9EyPuhds2Lj0WlW94pD
ouIXtW5wg6fJTxyQanNWbIg8zdYr2vgUz17251uwdOI26gqfS4NfR8nVqEVrXtQIwUTjiEAxKD6I
SwYG9s/7Lny2LVVN/Fk8JzlUbM1bJJIyEku2BroIWhjm3b+RH6AS1wTOL3dpuGDnmLcrkLShP34k
q4PKOcRVB2ulYYkxIGmYElVVW/THaEdREzVE8CkWhnEzyVvGixx2DAK0BnXIYch3Lq/byoFF9ROs
/2xUUsPVxo8b/BVXkgK43TYk6tNlJAUP0zPQi0ejcVgFZE64QkKgzRn4n3FJvaygwN7RGK4FZQK3
ex+b+ba8YzZQXYAVO+UXN49wi0FseYi3ceeneO2s8N1qr3e8+oT8OWWP4gdYDpmytwCg0T/pXO1U
yPZH3glfPQ+za6ud1Fe+C3kb0sZPuVWHAyjoxS4QHq1Iptn2j0JHAG9R+oOaOsPGh01TSzFyrcWn
cTKrc29aYRZ10PGtfqcG7XWHPrzdkE/p8Yg50VSJzVdChc8MHA0kNM9eoNh894rZkPLORtG18XFe
SrxBZcLW4f2NwTuXkXx4nPoLofT8WeLUmB+RJoKUn9wuJoIu3ilWq0qu0IBO9uV9Hedi2OK68Vn8
DsqV5bIpZFrPnARAOVSS5BUmiITj175mbxzwUtROvSFk2oWhRb85tdMrJ8jlS2RWSYTgBvd7C9Vk
hWdviz5PP/nQ6D9l7McnBuDQHYjuAsx2vf+JiYipcGsz3BvAqqnSyYES9svsK9i5SHFgnfd4zi1/
x0QYObdo52aMrbhwYfbUEoei9ZimUEJsqGJyZMpv9ejcUt+ptBSJHWJdR3fjrj5vHkNZXPz7Ol8t
w+Zl2zPUWaJ8XR4MflAs8Ajcmip7+jRu57bYEevwOQw/vFZwtcu8DtjofifTc5VG/dQGPN/elz2b
vGGDG+bK1X8/f7QRAJxdW847Oik9ZTvB+YEyoAvwFhflPuenAe/RASdk3Q9X2daEz2XxEouipzF3
14pARA6l0wkuyPXdCbwkHkGnovARp+iqobl4NTqeonvRkO/RtJMtuZtmSvfD9JG4Bh4Cxg0617uW
qQUcGFj6NTLuTBbYdGQM4JvaensJXNN/wy3VRMI5U7xSaBBFnFQLF3JOut5quXZYujIxgEA4qElk
54hpIY61kAMLrZ93vRNMXSywcdFcs0k5ppYIWlW0QNtKuo1lbZOjdRgn5jFJDpX2r1sUOCKZDvMD
gqqiu18hYFvOKsxCMBMf7dRDw8J1++vyMHDmYeDIoONU6PProKVpQ2L2mr1BljfVRbMSrf5+vPyF
q1Ns3fS2idcqx01cP6cbJ9FqBaQ/0PZiBYXJyweUbX8oB5sJMqg+qdqETeKGQUrNrNgd64FYWiuU
jKi7lYbiIO0id2zgCmyrC8nbgvDQA+r94TRgB7MqwCiaHY1j0Vedfua+EJOi6XVSyQQrkrBvXcwa
VXFajoG+rDIiVWXRkQIlPCLGaJf+oYZOF+BVvb1qFLtSp+/rmhcfFyU58DWyaUj873waoGHZJgIJ
qXeeC2vgfQlNLAeUN1v5+tGfpRbOdvJ+sLbGEcCppU4hJhh0iWuTWZTPzwyShSAdn8fXzwjOaPCc
DUKEIkj6JhKsYiuB1VuHY1oKISPVQitpBA7MiSOS+rfT2FO9FB003nQdnzizkK9BwBja6bxbMDUI
l7Fx6U6oEGBS10iSBJV1a8NrDkawW9iMdO5P6J5pLuQzgivMdu+VzXEG9T25iEIVBYjKnym+Rh8h
sotruCt1J2t9+z9d3XNOIBCfeKPOTepoKwE08HSRD3baDch+WJZ+x7B+4aRxItC5Tx6qPAo1Bcn+
9vOLxOaJUlWbckzDGICQLah4WunX5cOmZWY7mQsmheWT0WGtpGsJyc81L398XJygX41HgD1IXBdr
EBBDAsHzgCNdqQIUWYKkaHic5AEi0IK07a+UYyfJsiCFPdyhRycgg1jUgIhWA0xzbvHci8SdpeA6
mN09pmhgTM2hwdCX4L2XldPYdukWyhrTeJgbBos3pAOdo7z4FKpF3iB7fweQ4zR84rcx9CzO9VbY
i2xQpMopIZDZPgld+DzpcRoFpK8KbXXFJWBpxjhIG2uuAJ4KAI/6Icoo9nwmtx3l30kQUDlXSLcm
WAUB+x7dM0iW7UH7t4sZvZpP8C+V2tajuNbdeovMT/iNfBVjre2RKX1h8q6qRVlWTujHFU/h1HuV
tzsc/hYYafiohQmyOOcRkpfvy8ZMQ/LO/VIzCtvNF3WnTvCltGvJ981v/5F6+L7YlQLGaV2S20Ub
aiO/l5iY07x3YUQl8ozH1V2hLBZCy+mQlPq9IvBtA+THnaamWst7vleAuqt4TG2mOhCjH1KDil8w
8R6Dv11ncUsC5u98mUhH9///nF28LSHKBAYeNHpVqSGYI+wmqYwEk7WBhMVtGRvYZtFnsshRtJnV
90Vz1nLBdxnl95ggmpWm4+8PNjq9bADGqOiw44Mptr5LRWHWD1J0WkJsmgnoY1+Vwzks2tv4qX0f
3FJ4ebJaX7N3g87UYrGchnnFfUKbVUunhKg6CzlE0oXtc467xImklhkc3Tbb6xjqbhv7t1u5Tag4
cr3qfqf0rtFVFCn9t3OGI5QpxfS387KTseFGK9562Gnf58wuU/TnhUbcI+V3NuwXsrYwdO3yqmmx
4uSMWK7PPAnllKIpKjNjyb4f/w3icC9Chb1+MlhFm9X1m0QpILSXt6boYc5JAtL8i2Usc6+yBnDe
yzcRuZECsYp2dHmiRrzH43rxV4hBnipL2A9zl2dAPH3/jliEScpUzp/rJeAsZQYXhNycJ8Tf1eBx
N2/9b3PFB1tei2TqOdUCe3MEIloD35xY6GC+nO7efGFODllvVzN+qyKb0SB+uL/IJfjfkQeTNpqK
FG4xR+G6+eAk/tB5ytX4SKGAZQqevQ2nGcefJLzuMfIJiDB4d+bqDXU7/ENOcuKyOjk9ysCoCNGI
4xqPhXUZAj/JlCrMYYUOpXREOCFLpnM0OCnc5ZbdsCKufAjQZILBqTjB4pybBXrm0+q4q9EgXrfP
qJdli89OQWZTo3Sk6lkKFxqp815YHDmUqjghhDBytaJhM0i0ccA6nmW4Cl4Us5UHY9N0li4+RTfS
FpcSaNdH4AdXqwdhE14UzLWRsgFtHY/M4Op7zHrS1RfATrwF2gNvI2NUeNI6dzgHehBVin5lh3AL
FLmgV+LiOZ83MxM/EvqSgxYmYuISn/E5qdZ94EASRqKJarQUSTndIvFZmUYNPOllPpvlgdgB9rAP
fKUga8Gw7EK/T/Oen7SaBIAbuotBw4Clg6HewufjqI3AToKmWtWqTgVRUcHTz8E2CLAZAId7ThPp
hALdNKER18dPkBbx6QV6/cBeOSv6hfVOGPuY57rtn+yaAI73vbmgc2PDVygeF20jP+Nr/GzrB8Uk
vyuxx7PzcVn0T2RgowRvZdaSR6ZRjt9ouuJHVvMVClkNEKwluDAozsAcNr4gl7+COAW725JjMdxp
NGf6yRBo1Yg5utXhxRDqInrnHSOMHLf+0UeK7+URVGKlStGfUTdGuj0UAnJp5i3B1kT9tcSXc2fe
0I5DGBhratQW8Rv3Nqsl+sQtrEEoix5+ginsvs1XEPAdYHYpyYKdjWqgXNPP9tT82DGSLiXRjl6F
TJoKBm7BjB03vOKJTBu5Ie4jgkBFFOiklcS6FjG0ll+qkXAqJTgLN3MAZqunXySXd6Lrw7j7ORyV
+xG27Y8N+ncnFzXT/bio9xuFJLCED7TpUjijxRTR6yo3960PP76YxoXCcNui9MmaJBgczk/1pC4Z
DQTjmDpw0UDw/yVyBJtUtE2cOiTAofzukrihBk3PlB5klxRAupavzruoKjvqb627OsAqYh03n/xu
AeC07fUHe1Gn/FdRoZ4lHWJw12IRymkWSZg9Oct0KHhucpcvCv9MvVc7Mjn0H5Z8z3+9DOIp/azG
UzCQZoQPAClxSeSPbagSudJxA3a8pj+RHwka29lVg/w7Ay87yDgz0/0jFGLLQMsGAZJUg1ICoAZA
aOp5eLdrLF32q5dYfO6sqBKzrFxZeCtXLbSxMmm7y15eUmIoOetXD3UyFUqevMuyusZa5Aw+xiV5
cnsSaquIoqUc62Eee5ySNzZeV0g4tuEmebjWZLp7V5K0yvDWRYbIcn6lz3ux9RoHl64V02PzSpDp
ObX0GRbMuRU8Gf8qvClPbJ/5Y6uT5Wlxw8DXLMic+ix6IrYK46j/PSCqK4Wr1jTfLgYb+o6m5KCB
EDPcM8PTw+ZcmA+LR7tsZaYi3r9oQY039zfascWZmMKGJI1+zmHS4MJcrZOeYbrxdx+O1a+v38su
aMszVPToJx8KlSfTelYYRGq6/f/nqBt/QxgAM/d7o42xeUq7tRT2OVM3kTKW4YomnCLlMm+MAeoH
sjoFtRqb6SmvjlVS1mqM2J0XX4a6M2G6ZTbKMyUCJOwdzyjpS5c9KDKYVTIk2CGlnlLnOmVGkNAZ
WD+/2C7V+HwAGwfMZVW+oVDP0++IHfY++YvzyfaVktrcMfoUTevMWGLvz90RaATBTYB4Jp5oHhVR
/8Wn+spW/mfeHfRu6/CTFJtdGP4VOe021gSx3UH1sX4A8i1AogS+fQTxoWm5r4J1ZrOU6JGDiNPE
Y0yB3qOv2ORm7HoePGlzmFmZ5ZeUpOAYuS864Zt5Uxsto1ZxRqI7ADzhqDldb+HkFv916gLYFdAh
aN+QY09VtHWops22d6MrkIX0Ado8YOkrRNtHB9f9Q8cf6qx5uHN5H3dHofB9O9mfzREJdry96mKY
A+hRzt2Fyo6QK5T841f8ATndLY58qkU3XuaXL3fMJI+93ECrj7mRDrMC/gUxmCHqMQ/b/wAoAVIQ
GMdh/28uLCMTTR/A6pBlLO8PXY4Yu60z7vkTlROUz0LF3WgoJTYBbbspCaOsgk0OCSipV1wvAuFE
OG29UYeg+t4ZoR6yinITIJUSMHUhc6AwQlTkfHYwIHfYFgkxElofW9MjbROg4xKCP05/V1PhoY3I
u7POP7nQhjOr9i21yWpZn0w9sX5sI91tLAasbaJpzGVKD0N1Xd8llQYJ3jhfuOzdf8m9EcVjuWoD
u3deHcGfaHFeW1iHbfA/jeY9Wc2cV2qZ8eSF3UuLkT3mUAiavzYT6PSuETIzEn4F1GclXMifmwT6
z7afaImuT6avK8FS5LrPCUIvHqoCcPZf5H9uw/kFd8A7adkjjx5VoUx8cQLxPrm9peo7GCKcqNPs
d39MQ72cezuZzjg2Ayh8mmT+zD10IM0DILOKW16L/CHh+j+GJykAD2mJKs89SALLbDeb2aWOwDTh
nBn9yEwGIpGC0XDN8dpep1Nkha27Ya/vyQQb96lN7tpqus08kq0CQLu7F28TAOvRCzETktZ0SDhu
SI4Z/5erErH5C6m03t7FesjV8pJTayfI9QINLAizX3sl0nE4gqeG2y+euVcpW5R2lSpO1sCkZeXf
jWMIVkek1yufahEX+60DEkVaazamHHti3RMXbur8SsNpBGo6NI74dKkg6VbJN7NsajL2o1hSibgi
6Vr2M+7VKyo2yVlecNDJg6jFEYtR7Xi2wufaGjmtqTcHH5EN16J/46Wpz2R5d6g1VfigR3O80v9v
E7nzB927134p4e8Roa4F0mIkwopH9Sefl72xjW9Aao6gpvNYb+lebNBKMkIpG+Sy8g5Hq4JAZ0y/
aUgm+2BIZSanqSW5P9KwpWSGFHFDzCT4Buofy+1YkKXuYB3H8wgfrvREx2alHujT5ptxsZAu9Jlp
tb/Ek3+uipRzJifMubg6XuurzWQgvinKU3chGL1mlCiRZozlUrHLEXL8UX/skI/bjv6/DV2Xj2x8
fUEim2oRMgaOxM2CHPg9bTjdThAGd4rZjRRYRjnQw2dBXsyTHqAKM/SHaGQFCs/s2T1hkioVXtkC
XYKPO5JIy+FzocwUFTNr2MNi5bi8JXk7yfk6J8GwO1IvO0gYjgJI6oEc45ollWjG8tWjj5OdllYo
P639G7EChV27fT7gnChZgxcKxYhhzDpEYzx8C7cYyKeRsqYzKCG6JCUKDSGfCP0hPdF3YY8X6w0l
O0D19iX5vVR3tHlgzOQ3hQCZ8BygPNhS74IDzNfapWDt5PaPW4ZKkHHDifnBElnsPUsP9e3xQvi0
iC+TYIqOQnQCfBmsNBmqdFqGycIxPMhnNvr3oR6pYYxK1pdVnGCpZLtKW/cLZwlKHozwpAUHeO14
oYRRoRfnju2Z33J6QpS8aTIbSYsG6T8//qSq07x8nV8fqoCmIApq/GtNcEdCMb8XClyXisMVJNCL
DiBdr94VI26Zt5pFg83N4f/FV8SiuJTbbPWwtACz9uLPt9fN2LmJfsYBsPhtpx7iBxdkPbfXAeQF
8t4w9xYz2FRrkSd2F91f/SUmElMruSvXxXSIcROcswqR9biAfVzVefxwpxeuwRAsPctxOxwKk6DU
mQLNnAvswYGRPBdXqCFpQstiQPO95iMm5ERPnbXhCpCK/PAVFqbxta/D7DcxFyZmuLoHzIE+mQcn
GON6NHzizYYLhl1gCZoH7xnH4qVRIcTBMgTieEhIoIMWBWbRqXdbjUJDQGF6UDx/1nUxN+K63COV
J6WGxY/TlLiPEN/E6gs/l8FrAZOBm1ggTzyy/fs+W3OlesYBSzhX2zn0V2jAnn75m2uaM8uQQppz
x2G2Elq4/EdFyQUeIZadktzOfXui9jyFj8aSgL736OxK5uwVE9KKlzsoHLc8SvuFMX04iNX30btZ
EqoFEzmc+OKwpJ/yF27Hbtha5QQq/z05jo0XX+Id09sHW8MGb+n+ixMDWPnkts6WC0X38TFvRLmW
3FELpF4HROvvP8zoNO6W5NeIMACeijob8HvWdvfs830Q7KmdmxN5sLIk9r/eVyZjfGvtqfbou+uM
89BW2LIhPHqnFPPVg2+Qisy0d0miVwyI8tUqRshMQ/cgpM6YZ5HlNx4LaSaMiZHpip/M1mgTJpJY
//fopfB6uIQoNvji7V1MlrfX7kCU0UzoLusro+iW6nP0YiOnSgDeBC3P/5CIoxtEi1hITRZiNK7X
xnHREZePZaC5+prz7Td3sx5qCsINp3da8Bghc2Jd/6SccvlZvD6C91K8gNSw+nrTLa8IGT4R182n
rqfH7sBb15p1eR4385HDs2i6w+pTtnEGzFQAJKC/0Ug6/zjitEJsQDg5A+0NC1mRNvfvaLuljDMz
EJZNK8GS3t1t6jeGn2xIUmYD5WpZ2gTZcj7hpH1cyiLv9t32xxxanFbt3Pkrst5vkyL1rj1mMczH
LiBRivoe0jbH0TM0lSk7+ZFLQCseiLRlnBFSjWoQoxzrqWi/B5MCPaCcRI2qJ0R3dM3wXaEWUiSm
kBQG4p5Y9+vYw2qPPvCkT0WQzu+MhNHdAywjrbLSwYUEh34voKVTXsk+kxHbfQFEyYvEvcGJTntD
xOIc1Y+cbjoS27+xszIjmwywdTI4dtqSBqeVnA+1Pu118yldFR1D6mveybeR1Uaf0KtUU9gaQ7ev
QrqcUSyHnqbnp37TxGN+Rzdz6mpl9BXgtwwOhdclKzWjsiyGuDt5mztzrHlirdJtk9hZY4ssWgNy
wSlPfiLkBy6SJgLf2miZ4wO2wyJ+1+X2OADRfZM6FAPNgrn/El7UjUsJwJYz0RF2r2+8+iWpUnEH
f/BlZwmbstBzpObOhQF0t1xgo4jhWt4MSDW2TQZeIGDpVmXF98Cjqhye2TI1hH55fhVfucZGmFNE
n7mC9QBX1fcPMoGcrpoijGGpbisuj0hjF5NH8vnO7f+VbHbM1VDIjPk38feDRO7Dlm2ENcXVllsA
W434VgUZ14sAFByZYUROzgzFf6MbBLPgTioShmFizzaZ5kXUGKL5iPCKkeQ2419hlI6xsk3K9PCc
hF4je8VC24DULalo/mrDIq7Z6itqut841W7oo4PrV3CpEeqAbCY1gLpEc1lN+bomlD1pfbXYeD1m
J1x6D6iCwzHNLWYvPHl1JFEH9GH5PzPU/z0Bw/2bzHFIkxEE7mWCfEyNtpgcN29BVn95eGwb8pQR
J1JspeNBUziWFbpRFxvFMjYcZ2kHurmmj09axlcLcnvXeqZiIxmfrpiq5K12j6Mu4UJ8Rtor+ROV
MT7Xv5m12o2561qQBM5pMnSR9S+ENnP/uFfk+qUTqgSn7Y1QIBngzIaaUyC18AB/tFp34j5RiJdi
igFqt5lARsk8ctXB73KdYw5l5lzjFPK7G5Fp2CHJ/asnZhhOnSVZS23bkhu74IM0CMWmLgVxTqq1
Dg1zxC1HBOD0yBuHIs/+GVNCsVNGGzjD0kJTnQWWJfCv4GRWyPto/jwOSSEJY7BMZYoWshWOnJee
duAC15TApA4g5kvIrkbPGvXV5WinyQ4iWH/V90GdGd0Y4r9AL6gNzD8gLtf7Qxc7mxVc1WF65qOc
LIZn5VtPZSVt1xI0wit1xCGVon6uOpdYGQv2u+rw6hWgIl8wJezTPLTDniUjC/kCagQYvsgSzHjh
U8BuFUsWdLPLt0fZTqnQ5pFCAqAcxD1wvRlXiSBRrp4HbRc3VNy/+XkRA654Lo6J1sfwdRVXTkeb
ZdXPHcgjooqRVjwrCsNLc2n16N2vX5r2u2gNpqZN1vgKfWmQvsfLOqHHfUzrdGskGCNHif5GEoOr
f1sKV15LB+CcAc9MibJ0N7YIKcN2AdhdT+ceD/SPCEXULLRCooDowT67Mhb4ZwKZGgpI16WFprDv
YcH9vl2RXDz/QRuuSsSNaiCH81bYExFk2RcLxAOjxIX2woBqcuJtypGsTBYuGZBSyyUEW6k6zcqD
+ogcEc7GKA6Ebo/ubWgG/N+xQ9m8xAA3uQFUuQmFhN13A82vzyrU6PXQK4H23am1dC72PSMBF/XN
sNlLLGTk3Yor27f+K3hQMRXKasGvR2x+t6PrsXegbVZGS/min5pwsL6BzG03bHEDcYbifjHIH8y9
36nHCUZ0otqcrym5epG5eyhS32OwI+aMGrETwEKi/+tbFSECb4g0q51SvMW/t/GxccCx/PpUAImi
rXhjgdoe1hOOlanWp+b3XWcxlcSdWb2SgI+iK9gk+cBYL0VY8K7HZaJkP6JYlEm94rVaKZ9Y0UMh
54SMzcWIZ4zLnRO9Z+hMeNNNKloo9TqxVuaiIk5nWnONP7Vf+FHHFdTj4EHiO83mjcf6/m0rRlQp
nKc4moZBKi5RIJKc38o9GOCFY/7ZXNSIYGgicpShYMGWMQJvqRjKnz9QWHQiryENWJP2fYUmtvli
T2L9OpEPYXD+0HmODecam+zydnOHufDycqKP6d7mW3VLXmhWeL1I03FxSQO2Z707LuY44tz4zLQo
fscRn04O+rCWpf8Su1jr5F1Mt7Rv4j2s0V3sBqBVlK94BJ84EiJdffXZNBdXReRW1ZlKfKTD8/SR
VntFDUtRD/6dKC8m/MDi/uvh5FvXjxBzBYMBXtPA6IkTlvsY3WOKmrTIyCIeiIgQTfLFlC893QN6
c3Yq2fMIHoJhJBRs26lkWs0IfaPD7tqL++PX+D26Uy16j3f2azRVHwmSB4xpYwNHqdx7v3XJUB2N
SbMbZM0Jyy46glIDe1nxsiTecw/4uaK5jWEGKnbG6Sa9mrt+P7+aTcqT6x0P6kmPK+z+Pj9idbwg
q3rbgLK8xkmN3a6BZuoqunKBWd5UPuh5++BoS6QaKm2yyvpoFMpfL4bR2B1ApvySPKgD6L0XMpXu
jg1qdoXatyreVpi3jRaRge6+TOKq9J/1L72VICLqNZkPipiPfvGdLtCjXtIV4++d3wCn/eQW9ENK
LKquRAu+7GZ4QQGMW6JcLoUrQwa9DNxPWqqNx6fhgO7sRSu7Tq9JUvUaAEMcroX1gh0bjwwTGfNc
hY9gsFGTQAVzt4Jim9/T2c/iSNPzhu48GNL6MQYnHq6z5st/nwvPAr3GtWXDsrkFobBS49hW/6Xa
wpe2RljckcJ+8TRix4tNTFW/XkEE/111EGC1m25qshFRjpHsG33xW0JfJHa0Vhm2P6IT/uV07jAT
aXcUwtlmuxNI/sAoTQlX7xYkuA270gLqemylf8q5TiMgVtre2uMzSnqLS97Hka1NsASJe6WnHNfn
5lyzcS722asw16pS1RSPx6h0/+0bnJkbkgaK14NWRrxFVCrwihDBuU8ddDusdU2n5pIU1ItgvbiL
r9c0bByC57q50P8vsc9KxEjhUuTm387lwCaVYXG08qKsmgMkp2oAy6MS6iIF7PveXHQFfxWpdyQx
7+B5k4tpFw00zPx1py/ebP1X1IJnlQaTNdDBYZSdpK+V9gH68tDELlPSWFQq15tl7V332ydvYepp
KLCFpe8mjN5KvBCS6T9pP8tTjO757o6cQJd2Z/FrEOrrg5V3gCQI948yCpyGgarancaQk9R/4b10
cH1XME7Jhu90F2gV/2bqYz2J/0kCkv+uLsN22OhTg6DttyPnJrnKwTjkK4hxYfxJILB4KFW7gy0Y
hKhvUUIRsbs1TO5x76nM0A197Pu5LqNL8IycPYkM/pqmVz7DsVVrR6r5XAOSBWEhrKunv+jpSGSv
5ahF46cn65HJKS3sMPyNmqjiAOqYwPcjisN2hvD+OCEfA87r/4KEirnoOaF7BOu4Zh6eKxhjToCh
Qw5JDeVFw8lXcEmUx61bewVwXThC5qGEZyannornT00XOKZPkX6VubQY8PAl3CEB7U7mi5hoxxK7
oqZMqGmMK9cgs+dR2Y/Gfrs5IaCoi++EDdcApQ/GkWCtNa0Epyq/hfqOGgKJRVbyOv4LoB+OtSc9
H5Ix1x5HSS7CkvGEzUjzkXBzYfxeGctaYp6O37KUPz5m9s+nBBlpcSZ5nqDRcfi8T9K90QZWx2Pu
k47NI7d+0/NGY4g26se2e7WPyMcMJ+Pkpa3T2iz/w4ctF6WGmq1nvhTGtOeRU0Im3TcKaJahYW/g
x9fzrpzXH33XzbMJgJWJz3cU6tXPYs6mr3E1N6iDdLs5yM5AAHfG+Lw++eaeD6PmtMAH8dTJNgFo
b29ePdC5DlBtVzlJq2XpU0jBI5PyMsF5ms3otnPXmdXFVyiqBl227TECquq+6AIO3O+S1Wc8MXht
WxrJdg4FbnvMKJ1hTMfzWbP7WNZwuIPSNOCOjWSOhYq+K434J6UG1SVYRRpP7Ei+ls1f4yFnzNAI
R034wv+G0ZaJDr+GXuWeQGayzVfYhKsRPE9vssyX8ZN9eyKIzthXPsrN9zm3odsh3HrQ8o4Ozph4
y6wXsUSHe0K+36HBV8gEUgTmS+X0PJHm0KqoIA+A99kxsEfsGfgS3sXWExitW3L5JSHH0Vf0d6Z/
lABif1c7Q9mBFENSwmMC51vW7gb3uhYPg79MFJnFKM3K3a9C3zT8q+T/aQjJFZAPsuWnYlfBrHSC
0bWmKcAOFeXH2xkm4CyVR0Zt4/nIDC7L6bYyq03IVjz3lnS6PtfU3hX7tgbRKLrJzeDbpqOJZZ4a
kc3KA+eI4XlfHpuiPKUl+sHd1+DShisnkXgNfU6bJ+krtPJSE6JwutVYsnHUjwKm9hru+X04hyoP
peeByzXJ/yxt0LgCD5D43CucfHlmvtGc5ufj+vTJIV1EmlTZgIcAXwbybMc/rxJE0CE3cqZm+eZA
RiBXKNh+LY9Io88EDglk/xpLA/+K3BE9AloQiYoPd6M91lkEe9wCa2Q0Q87+qGMTS1rv1XzUWgnp
ZQ44sZTkNHyaq94v+QrIOKRUWvmhuKmMMB1+J5RGEjbprJJSPV1vt9pLdRft2AsLZzXNwjqXO+NX
jK7Edund/ep7sgD0oGyL0kv3lHbk48D6lM2/lJfD1NKV/a+tU5r5ekDNI9GjZigko8ygvWX3oNLz
FQ1ifrU7YWeoomXzmOQ8BECboZpT2Kdw9ugCLqvqH0Fy28sA1pxaWZAspR2uRpYlT23XUwWRqPbz
L+jcRuI5wM/tquRfe6nNVDPjuNlOVXjUIz2Cm0mMPjKEIp1QmrGegGtd2TbcBq+lHIHQtJIM7Fzw
lXXNa+TmMk2PiuD0ndSktkX4QRjc1/WnG1E38Xm/CNxEnM6FpZS+4DqQRCuOc4mmEbc7pdFmZ8SV
APzaoW7gAM0/WbWbykd00rcKNnBz8QgEkaI7FXoYLaiAyBvpYz5MRCekIfVjJSBzQjUtoNnv4LeJ
/Z/4Gpw33iq142XU8hsyXIl4dBPDKJ1qsVYq2teAVUPDSPyYk6qDsTRY65bvMC33xwXC3iah0R3K
cb5r1vDdcSQZhcFu49rPQPFEumRUBSb15lhN+b/RDDQuNOc9j3CyXp0Am9ronQaIsHLGuZVCUDPc
QSq1myEh8jbJN0FJ0ML+6WqZskHUAwN7sR77LeOLgxrpJwhKL/Ru4+g/1fZt2Wvich3qeiLl+Eg1
jZeLFp3d1aRoYbXDJswzyDo8cMqMc/7+OwTnp+uzGgjc6zn+ZtERihVeYJ1h/7FmYF/lY1Go2Ox+
J0PdQgEESORwuQjYVMjGb0/lvYlnSe96i3PNnesNfLFVEA4oYPpKa/J56AF5hngyANJebrFeOzRt
jwYFTj0aHCHc/cOc8crbBe8V/Leur0XSWpleMeOlGqSodGbWX37b32FhtV0qOIssbkqmq7vD+y4k
PtwdumORMg1mKdIqO8CXbNNmHzLKb7ZvsRhzFSSbfUpolOj7DMLW0j9R4uC1X/hCa4oQMabZyhPg
SYJ++sE5SqvYMDLzprBx/Ensh+XUs/RjMbs5RgNg2HLZbpZcGP0CvFPtBGtjsRdiay3sQFV9P4H4
TekbFiJgi5didaoMdlUAjGZGsfHpVcKmtBBWAiSIE1vvgGOQ9YC7DGV9LwgBO6hEbl0315Ryfsm1
C9wuAvQ8kC7t6/iMypSHPYrvIXGN6IdZfle9e3LzMcHvYQ1OvOC+tFuFL0OTjykhjCMZoH2KyGxR
rCKrl0TrbLcmKVUQ8OKiwPDomdxRUUbmTOFpdyhm+x7OLX5rPkfvP/Zl4oFTzAMf3ZBI0MKSNfkX
J6KGZVCeBc3A6oYoSOdvRDEiR7DiuM8vlzU3OdZ+XCultBCqSDh8n5pPibH07RrX7/bA4VqluPu8
cStilV9nUH6B8t58/Ql4R2B272q6acXrWKR7OwIYtl5W/4GlJA8S8OnwE6C0vWQbWhLof3HeyvJa
uIubse67ktv//0U9sDFPKD+9RStnJwtSP0HpwQNGP/HbtTkrMpHd7xpedB1x8k9BGD52DSvpzx3r
L9EF578vYwo3WXhSi6n6SxuAF8NL2jXseC4/EMOfHyHT5EX0gzCZNZn4uCxzeod5g3qL5nneZCqs
s4HeKNXMAwLPCNPcQa+9m44qQ8fUgb+k+/uotjXzmyyVaLsliQEgtgmgNAQi7JYfKLsgyAr3RG4C
EUqHiuC4sx4NP0Fsuj9shxgnfnrUQNI9pUqXLcMEBaTrV4OKQAvvceuqLHypEhCgYA1cpB0ARdMl
PzcvSFLADEngXZ1rnIEufXxiDelkHKW7RlhdN3r8eVbOO3G25EMPDXMiZCoZ0KJgMYtWRDBRtyuv
QC84B/wnm57bIfkQfi1qga/LWDnj47MA8PV4d+Sx3V5lP8OvUGIkUONL/j3A9cbH2zBreYRVkLR2
cuxxTuZw61j08k9DdrTEeADOMbda0ki61wuIeUZw3LkOL/TrgA7zX7AjeIxzdHrfRMHa1DHWrSAv
PVqFjYokb2BB9rUcGdcmbx7YmNtuj71vDoUtJSKcqqb1mFkcffvgmMFvdhb2U4PHNX8VXzufacF9
quh/3Y/cfyFsU0+GwHCnPUK1c1EOsgUv1OtnVwJksiqF5ZHXBRnNb9N9vuJUULI3+6ZDEIznZUNA
RSi5suWxpPbJvx8xP3RxxYYJPu40NGy0EHhTuh0Z2mRt03O/6E/qdCE9QWUgJW6tmWmpRnZX0c1H
Qc3unCAYxleJR41bThL2YLfCUWt7rYo6gZm2JdpdDevi0DnBtjyRY51wmnJ+i5FgPcmPjd7Q+H7l
z7HWyxihKCW+QrdlHz185zHj07gS9UuH/kGUGLqKtCcab0Vu9rOGfm1S7pNqXMmdmxHfMaNxZZkX
hLavd4gs2zWSlyni5oHqWp+o5b3BgXjl4cg7zO2e7TfxZxW+V1vgxaDoqUPtTQQ0KlIgDFsFVsp7
OPNdiwMzdlv4gWQqWjW0XG2OjzYZhZYQrQh2jFYbOHNlyXgj+0mlIgiGMPzkcWIuqjX6OO21/7OB
qL2jxiOdMrFuQGbAT4UAoDZ6QnL1IFA2Zf/zhnt9coAGJiG4d72RNs2DA66ujahslT/64MsV4aYn
K1oQn9iCyMYKkXXRuLsxGafH0Jkq5vGtY8Z+XDR9UER1SWaBAiumgHmf3jEQ4CcQyiek9APmUtiQ
/6eYrfiCQL8LLW8jKAeKkZ2lmN++jVr3fwntVrywqbNUefjU9z1H0+26YUUU6Gu4KEqO1MZUkaXb
ElS/eSBcbCjTSJvRxIeuM/k1S4vQk/cKLezwoI1xB4aITWlcv54MwAz+NKhF5+v7YuLX4j9jr0rT
sOwPPTbOg3xwk2ax7wUoqNJdxkOla0W4FwJ2hM+kEMFPpA/KjZaQHPBU1m10endLbGoMtXiLaEhc
bjg17ySd5hwshU/Dx/sPvSJjGBLafi5IQ+yMZmM5GrPO82uKYOSp5YO8ARFrxIVwxsTtstyn29z7
4AGYDiEHyBrzqhbEXGw7uUENgAW5k2bWzKWEpcJqbBkhwxsbZazOwlMbsFHUcIWyFgCssrP+6vGD
Gd/YEcSRL0cw/5AjsxxiQiIRzHysIRagvX+Kpn/mL7KHODpoDr6P49xsvZ9sOEVYLd3B8cR1Whvo
nyh5YGBUPmqsBx8//1zRJEn8F1uvsQEhrJenA/db2GIGcVHu0XMXl/6r3ONSSsxkOmkiRR1dkagz
Sm6IZrr1W+vT+JFZAT9j39+BYtQls/YbMY2y1D50vcaN/m6Y60+HCny4kGsuL7VK1WYHr3MKBGbU
iZQWe8mucEqAojlc067fnEIJClUsWY72yVuD9q7lFcTjpd8P6jH0lJezLXYfFgY1CAanuGGICguN
K1lA17KHN9inp6yZw8p+cvPZ6Zxcvv2yUFyAV3Jxopnos92C/PEWYtBdMaA9NCwY7mxrG6yXcnjE
IQiiuH+HCGQ7dMAuZqshZ8zfkq7w5bHXQSX1Kudd6xZMDQrjgwDfdktisPQENXCVoK1HQMBz3XU8
kFlM4ugRyVtOQKqWIH3U9e47A5YqfkZf++tNd3h89d7vj0l7X6bA7/Ao1KMf0rLzWmzuYTnYiXs0
5g5O7CrUxqpP8IirAqYYdfh4AzhOnw2TDRvao6vQ9sGfFwvi3miUPdkyXArRjqoEetrs3dJLKav5
GvIwpLTfVy4Tc/J/Ypq0mGQESScIvFlc1NiDWn7hfRZmOn1or/BOK4dB3Gem6UTf4lYslOgOMfyT
Hag3B8blt4gL3BJO6A8APN2HtoqqmxTs8t1EH4R/ZYORFzX8nT0OOfx/sRt6xjYCVjVtZe6E/VyM
M4z9ZXt7b84mvpHynuFNiMqRGI/3RqbmniK0Hp+XwiROLF6iMU6LSr19yuCKl+iOFzRq0aCV9PAy
hOPI7OHmJ4/Qxt7bTZnlL4/pUEP8QRLK2Kho8fD8TnmDcxkht5Fg0FfrFdfyhd1V2IjhpmCYsGdM
ry0/dwRdxsV8A+Dj2u2xuq1yR+3VXuqeQ2mdAKYPjVP8hJKAhVHNLDc5wxnwp7qPOvhXOCXDAE0Q
G/jSFeRugO80HtNLdJ+tw7pAb5rpIrri5JxejmZXjcoqTgNl5+HxUuwVGYW3G/IXKfdPHttT8VOz
s9WfjWQiFYOq7zce00si8wjkPxCZfz9q1DTvlFFl50tOWMgVrTAG3vN3pTAYsoyLCHMFg+KM1zNU
aAsSwPJFHufMMI0irS+qTKVyfhuKlrxI6EA2w4vouRkIgwBLFjCryGxW5u53C+84caaLMnONxEc+
6odNLILTVQEMCTwD2sd/mQBcefICRJxZM6jBjVgJm4ITY6UhNKF3WeDHLmbyi+eer9FQnVUyvT//
41xwg7TTdXzzad6YOzDoXv4zcl8OC7bWBCr6ROEVFdTQFtIio9COn+KhwefyfIIoOGwjfhLMS7r6
72S8T6H4KK9g8aBAYmaJq8cWWivQoUrNGluwnlpZepgFx/lIAOxYua3HHrt9O7VZh7oy7ZB3ytLP
3+On1oXFd7YH2dHM1osU81kHQnAz3VKF4R5jfYqfZt1QaLYUAdDu9YRm5190sXbikHv4UKz/kRTM
5d2DjTaJ/IsJtNyMeKjgfFfOxLmc7ZLXOVaxXXgiZ7WFG2n50kpPtdc13r922pY0Vx+t/tUdYXGo
6gF3L+ORZHMrs95PeUpIVf2STBtj51PK+cK1QWy5ef+XIEE8DLWXKCKoNIBacmKRfGVwwMfIIrxE
Un1emGW9gjmn2rfnPi1LX4yBiPk/qi8YC4WDnnW9iFEgzE9PxeBeU2BN3SUOyBV/DKrFCbZLpQa5
Hkn9wSU9EayyuneaEtBWMDhI7YrjDjdOxtCn0SY/GqRCJ1/X2xnYq9OMT1cE/WgOkGV1F6mPCFnF
FgsdH98doqzXTafT9DoxvHTklfc8i1pdqdf0M/wjj7rI8B8ZUqKrANCqrdhOQYQGL2VAlKd2Yl/q
ZvTYteOUlTWSji7U2sghAx9TpR39zoanSCEOl+qvzAu/OiXIRLH0CYsw/K8ZzmacpW6MDvqn/jyA
nhpllpnJLpsMDKPLDKUelacY5bhQIccEnO0NjeajUMvF/3fvKf7/YU6AH21xLLNafFVUHDX+FfRQ
TmTAeoK/Oo3LYGNMB08d3nZn1BSXFZQp2M6CFMoAckwA1BQ+xizyFZ17LEoMDSAhB5ymgJIkEOKc
2xiN4vw74mLB4DN8mbORUF5NFdgQVO7EQ9uLj+Tchy+/Ujzw8L8pF2sRa9SA67HNR+F85rrLd3tf
uRNYVIFngThgUYQhk8LkA5XZjAKvztWS5PiHysSfZjtg1FYjOQuOkr11/McG7ijoz9cSYXWptO7w
UhFVPlXhTkTd9PIwYu4Ml+hJ5H3i2Fkpm+KgrgPVsApkVwRZEaRPKn5Xvc9GLoCiDLZxdGz+7mod
L0BSzOrs0zUr7e1GBTfqJBqHHbwYvVuWGXofyeGrtT0LN+KQHCHhH562JAzy8B8wRReNCAoh1njB
FN7NDmVVl7KVnVltIuoWDezyYNTHeWQm7Y3RzGZ/piAc7K1mCNxXTQk1BHwh+kZfQeP3hTmVWUrc
XCaXEaVxg4f7KXLwnkMEBGfs//QRl6OMSbz9KIFtoPBnCZFAsrQoQroMm/ERH7+7Elti4v0gA5Fd
lZzAhCGJKdHR9FMOSWiKOkie7LP/HPXe6Z9FNhtGhrSweq40kYiLV5wiFFrsiyZTuMxGJ7e2yc9p
xansoCFTC3uULO7R03AxRHxGEmB9D0UkcRszCKted01P/818t8nk6HlTsToXmXh237WR2AZVy9ZB
oRsDIDnoDnyq5x4qNYiEXLVTlF8eXZMShdlO7V+kjAXeaxAYtnpu/r8+U8pChXtDQgvMT66lLkr5
R7fPGOvKEqJ0x4xzF84UAT33NWLZ2F+NH25P1kRzE7g/Ojx63MyCmGEnW8gVhrswT8OD9yCG08nl
gyrr6IgtjbzPrteclf/KVU33SmXk5a20mDiJ9oUYwNMLehKEUDutHAoVPSVAZtJ83g/q/qgpSDHz
X5VSi/E82kTpkGROLZWkRv0wvcNarIoVnQsJcZsBiMnmiis2cpVAaEex+jvcVlSAflGD0vrvAGal
o0bd+DaydC/HA5Ud49mLxUO/Xl2uXLwBR+ETV1Ezdnt2xGuno2hFxuku+eNOVrheT2I1yRwr0pH1
D6KMLJmSWAyZDRlWlUy/h/Tk++OQLUfD+rLeDeJ+XRYNPi/u3u4wO7haqjkWnJJKtldmTD/sKfKP
BFRrKIt2FU1TOlc50KcF8NGpjVw0CDDbIDsFqclWL4ljt5xYxtd2DoGitohUVozf7bH1GfZCDq/S
C8egDEZ5IF5dQfjblH3LKoRrqSe0pIAIZoPiHCtYOEATkEAtfPXD9KQ9JhiyLhMntJYmnprG6vBQ
vIYF9q1CsYX1e8NC3LrtnbLGXm5T8OKWDkAyM7+7Lkq9OHlb9iEFpcJYz+HiX4Tr6iRz6P7mOaYb
vPotZGub8F33BClk2wJNu90mxGizTtctSvSQG6ig0J5ARD60CmwNd4qdFPHCZw49jNjYlMNjfA+M
6sw6Gxl/W0s1YLHX6gzwss+2+bcZRBOgvTfxB0hsJ0iyv83rP7efAWNjchlppuFuktbcIJeTrfgo
0XZJSIE/+IeKwXW3hJXb7E0Fy1S4jnxs3w1R5DCXZ67jK+QZCXIjAJmIZtxMnRegdYeJV1CQxPDZ
3m37Fs2gUg2KPtpe02QdcZv3pnqjyPvW5YotdHTYmbrdXeMnr1j25AoDyGzF/dIqw2Cyhnty/n+B
s2DtSEFPkXdp4q05nFOHOVQZTCR8nplF7eux9fgnGsKJd4g6t62Atrc+HctmHJ0V1EqN+xwGjzYX
Wc22yj1pXEJriKlGHGnAg6MFoVo8iuhKUiwULCUCR1rjntU80NqD5ys+//nUgCaHnNlOpuEt4Pmx
mHyQF9l4828X2/APgoArjL6VYWDIau1i7XRF0odwJ8mErgdBxTj3Cb05O+7x4ezYJBtn7rrYtCdB
hpAYLWhtHb+LgwNpYsto2I+06IVmq7d3F02vghzIYwuiBWtsh6Lk/9OZKUSNZszjURY/N+xxT3rp
OkzFVpq7tyQKpFedE3dqHux5kciFKtFaFG/3Q47xTtKH3M3it6G3yprHsQ9yAx+GYEZfWTBKLp0H
hSGXGIs3kALIyIU+HuU8gZnaZzJn8EKzP6EFfi1MdiiwD5/FOqzKqPyjd4iDqovb4KJEwHpUpezh
m++5oLTtKx1zRCesxpuSVr7DUiXESOS5I1d3LzVImiRZe5EEHwgnXMVwr/YGG7AiNjJDJWaB1gZW
O4wg5nFnOUh90ePoDEMDxZTzmhrXw+bzsykvH9uBKQowovj6bsPtWZCEwG3ROQiByM/4XrkwRjw4
/j3UxKtZnN8AjFHYlxlwHrRWyatjAjh4Gq2BVQ01HpYByntEWM+GEFfitIAmAIebrZBN6GOwcbx9
Kuk+K1Cu2OzjQcjn5oenJRgn3ziji3ysoZ+tlMVHUcP/d3wfq3yCXycdQsodPz7hlpEmpgh/omRA
BSjNUPQNnGtO8Q8SYSsO4US62WnGg9ECpt7TZUTt0O26QPMGWrYTF4uLGhILLMWkeY9CdMoDq2Ac
xdJtKHT5UqcQYziLu/zJU/8DRLffLzGD9oReTAeVaXOSKxBlu8qCbnbjUFOdkXcVtR/SSn1Dd6g2
9GQUP42W4sIvuPX7Kj6lc7Jvza3K7eqtGR+iydQcZV9o/eep+PVBXSaqy3+jLo93Wvvofr/tWuSd
hTDYq5udfo+/kHwyoTXz3kYr+umRAnZ252PB4kZpR8/hgG1AOVWzjvhvlTm0QsIWSyg9QibABDTH
fhSQd/TGs5nsHjb9+tt2QyH/0wxCWJfKfMxdHzcXDMP1k6aUjizvqdZNtAOBvOgzPqC+CBYuszm4
ly7Zdtal4/NjNLCGR3SSYM9qPQnyNmjMemxDdI+imj1uVOXluqTqiEks0bmJgAI4JOoAcy0M3rim
+EJ7SP6uBVYuwqTxrlx4tKHEIKjoecrl2/06Gn81nzpoIMait/9NM6CmMZCtWJoaK8UMKUdeNSFW
MlWPRG32uxtrn5bpx04T1xoNWqwzsCrrk4zsiD58baoVcUPCyjqz2gcFwcnDSItMNPhXlnT3/IZE
fPOaByppkeRRUivkr821Hib4NUxkKM58E9vRTvglbhjwNnBLpGwjFWzanaRLYVxKdFJmv4lYBY9D
F8keKIdFNKIgP17nvY+Ybk7Loyjg1gTTzhP0RyXiYnnlyb/7SHLP/dcnlDWvWESVuoLLfKVazNOi
0UIIQ49+FDxBn0b7gQD7xIFttOTTj3P7KirRDg+mM+dWagVy9N+XCKg5kFNBxmphV9pHOjCXeWMk
Lpw0pRzxl4QLb10YThE+eEshaO6n4zHUhvGmh1Ib9f32gfH11Z6Bf5gf5cA5/xpwf8fMfm1UEmx1
nqmOz6wFAqZj8OVPySG0JE2vG2mFGcrcpJUcEeSfVUEVmMjPbDyGMWPxIEwYfnyLE1Mw1j/PqUMe
5UJPwxrImTVw1CKrnqCuUSy0oiv/A9Z7Sn88u0Li7feTBicF4Qi4QeUN8u7Oogi59DNNoHqRLU1C
6SXH1mtGvKtGeWeH3G/RNScJfKf24R6KCcK8Es0k/dSn+g+GEhTHo/rxbLGvJpGX6Na90EBrHcqR
OH7dCU6StxYfUCj2HP25vTpsaTr0zbAPix2qTxrbGov5ooMvif/F0DQKN9jDKFnDbE9ZK+NfDFDL
kZRsAZMQ9FNSwUG/tGutJRwoaaMMaMfqKlH6QTP9cWT9bqPCs6YxyfsMTcOC1d37F/9VdEEJiwHA
bExTFz1IUZ98AJU7Up/hwqomHr55BkZsBpf7Q/ZW6kugjnlnXTbbEpeSTCTObfwfPHn/PerScQKp
W8xgodm8gMq2A41pQwOwro8uTrBMuuP8P2MSgFx20/iQ1LCtyiqGmZeSPHOXEbR8E9ow38WyLltK
zV38iStyBQfJouyiUsPFEt2jRPMih/Br6P7MgnH3O8s7A7qPXXkhnAcVQSQWpilelfnjrN7RMqpt
ErK6/DSOCzxa7gt1CIHZI8H8Fxce5RKgO88OkWW7JFnoW03hE0OzHVsDxRYWy/MEFqwTx5tjjg+C
rfWIjz1AnudVr5zS6BPZ0oXlnm5Kwm88Vxv0eUZwcnMzBYzaSpkz1y8znsPCqLW1dznP5kYl23nj
IOnMVMcUug1Po+IhTtUlSpHiIjHWI4p+tJJyuo6QUAfsOq7Yd4G+GbnE5rKo26ydylwgK8B5jInZ
sy2WbvmpcMRt3VCkD6+6S/LLkQgtmP2bCdtxWQc++wy/IL336iP2DP29rAKcam5/VoXNjyBexuYj
YMDLIjW17l9axD6R22SRI69CgE7QC3YcU9cPC3h2G8MaJ1p9JUCYYhUzyYymZe5lEetrjLCrlL5R
4p6SCoEgsi9oxjma1biyN6KDvWlSrRFTB30sxgCpZ/KjLoytwfNJfL6siFy0SZSGRKlm3H/N8ikK
ICsGMBJkwxVAPNn4KkjWmv4kXvb6S2dMnQuY+3ip1muPLdDCrddFMpfNjQyMG96lvzNZ6p8XdzDe
KZ8WNMqZ/Oqk08it0M7aoco5D+92/el8xIunUD0g1eUeCc85NFyUfF5Ab48p9xkmLKHsamXbwmgX
ALAgi/cDY1mpy8KRG9uhXK2v4OlFjICMJaIN2KtaWj1D2/frkxh/HAIJB+K/QaGQZG4iQiRQKobi
RyqVPxbK4PgxQ/qgpyYaF8kDCJJrkNsm4vLeaiNq+KKIRSLCEQxvFF2PIyk/3ukhQglnQ03eqAQI
pZUeIlSLna4VqInWqh79IVEkSdLW8P+ZlLmyS1i0T6NnXJ+OsJijUpPEKagmBtu2qHMdbX6KF+D1
Te6FfFcLTk/eiskZdAbvCka9PvjoVF9KRHc0m+bGWV1pelmKiRw1StT/xJjEvUn8GQQdY598xkIY
hH7iWub7Ud9ZqaIYQY3nioUkJd8nrET6sxWuFttnQHYjNjSPk2klC9Ubh9CpuedzGiT4iqYeYk/z
kq8L3c4PsQrpw49RsZh9LeuKGeOsVKLlebI29CfyWGAL/zz/aWJKLljVYZs0SyP+a1uR8pbI/I7u
FIJzgCn6xLKYm6C+Tj83B+p/wmv1Y/RS7dFyevWlUtIMAXsIm4jt87xYuu8mc6/tbCSisLyy0lo0
Pdzb5bK8qAQyQcsqk7rYQO5NANowL+60X/fipTKf+Dq733tHXIMbiOXrZE6JpNZUgQ49rtNci+eM
nLd9sHqFpEZOoL95ddSuxBC4rMczn7WSf5UlAwLdl4U3RKycluILtiQVBL2xwOk+FyXm9fHrCLnD
JYDSHT8YmBjA7EZsrhIQ2f6XEDpT9NIxYUu11iGYAKNWuE749d1rXoOzRz6ZIT29ve8cYL5JT57B
fnEej21CoBENYepnRyJLJ6DeJAiXtJ/T4gpKoKNlDCdQ8PqVItzSHRMCvze9RHO89f3tMnB/sNlz
f3umK2YwnioLTClCprHsnxNEo4hOhLC/OjEH2RqXQma+wE96uWm4njOz6qU+hy1fzUSLqd6wzypa
36d2g7p65g2wJYP4AwZ8RxCcZpp2Wx6H2sMBDXHfaN8aMRc4266FLoYUvDdPKQTFWPUMwbGxVT0E
VN7bbR5tqc9L4+3DgWRCLg3W+e7N9iqQ6tenRg2DVd0qG58Ci2IeDLLlgav62RxUg3OHmN+ETAZB
LM6GbYMutxGLtiww3bHSeK8N6fZTmOD8wyJTq/U4gdVIgxxcreLGovGoQrtVoMxVOcLtDqg4c4Ku
UQUoFiA6J77b8B5qJj7FXsbI5Vk7wxPzeb5APw7GAZ6TbqUbFzY4MOwE5J1Ve2wHy2HlSwLSKWqy
7kc23GOYbmMM2aK74VLX0HjMS8OdWSmo1JE3NxGn3MQdyP1CLywVQmqsc8/RXs3Ji5KbHLIPD3DK
ihOEOHJOSFuk/1QB+gsJ0fN2nJm+L6K0UR8TwvAkop62WgcTIWNhJURQ5midsegmnzT7Sy5pAFQH
ikJ8j7eTe8vx3eBIH+dQ2lk+8Y4QF6c9LZxHBaBGNT0FdUdaYOWGXeZfkv/SnPJPaGi4DU5FEAVt
g9c/UjEZMwAlj1+2sS3p5gsfDnyVlz6uWUzMtUVQkmkqn9/06mNW0DhrfX/LKFpjSEyeWDQyeMPE
dn2gVGkqnkFu5XMynmKY3DWdMdnKDl0yqiKji4rmy48iAEzF3/moFhAXmafwPaiwFWRYGpa/s/bE
rjulcWXn/VWfxOHPl7CDzxl5LhlW6zgo+ie+UvZniY/IwNDTJmutBXGT4pcHaUEDpxE9NcscFWZe
lMpTFLA4fkFdbl2iYf8EsUgdFtQLSACr6C8Q6JfpINpj4XLGuTeJO82gdsMTRxS8mSTk0IbaSkOj
rLfTsbp55awhPAXhad+C3471FYrONOAp3KUiT/TUHvfOKRmc+2LpNuavECwFacamA1uZQuTfZ2wb
VaEEZQqEkU2cX2PAx2uhLQ1xKaJzJW7pvRilYtFQukeybmBXG6tyD3fdsU54drNUIDfB7jSoZFN1
crzrFtDZcqwXK9j29AMuq4gdE6hoigkz1barCaypek7VCELtfaGfuQtGYbZEQJsGuwLzSSWjXr3Y
WckmstAVIB6w1U6q73KlXY+1t9GAkq1U0cuU8p1DMwOxCXDq/Mvx/00OgKXlYz6YAtpnIsQ9cDK3
EYSekOUBFjfbPhPyX+4iud15pF6bQ79vksWyXVHlMeB9jDaGRTUuS2te9q8v6fCdEaZoTHm0ht2h
aHmBHBISfbzDNMq3cMhq5E4WPaEMADsWTcDVUSSm3YYv3P2lxEN7gNXWEFniVaCFSdFUP+fM+B9d
1j7TQf8XkNC/JwreUxKwDDMFXZjt2kZFrI8UhJPOBG3yV5r+WbUICnA95+Tv6gBGupkD6Fpq71tl
AgFwBO7GQkyfMrNn3+JYDomzC7D0vNMf2aqSmGiQtT45RMGdu3v9pQ9mWlJXXlqrjpRHDCetavCy
ZfxjSjNZwxbM2DcSAc/m/UDz/FGkn8WZeQ8sQ+jrSO9du9r38NIKl3uRwFzfjG5yW++jQZlRBUNU
lF4FOrLjEej7YLU/IF4sw+HmMhmvXqGdWxpVM37pT3+C3tMeAMKYhngJo++q2OsLzMLkhyMAqfhu
ze108QCMKQMWFXXuSRGz7CBKrd0D5cyY03Vn/rbHYpwHV36BvsniRc1+tCNBsBnYLtTmnZkFGQ8j
yyGFCOzj4sQW3TxgRQpE8YtVrSk53noGmXKy7hWj3ihdHxCGYD6duoAkmEhfo6MDDJDRcc+NRAro
mo5bnBjpnUltfmT7n8+R0t/vXsqftYYHOkAOtZT8OTIpN2PTsZAirE8/fUavPOBjAtY8nGd66c0E
Mm030VQUqXY2g3NJMl/3afVcvrgrPpltESAP7+fJ2nKRr5SuJQwDXRw7NtVXHCR+vil/dBIEBJQU
UZm2biRTN+PuGdB0NiKJoXk4mxKMeeWrkSaR7ShNPWp6/XtYpmbt7Ywg5sVsdMIeVMLb2w7sBMCf
PaN1kUB3OpN3NMoGgcrih/zYyAHat4YLrxy0MnCJqjkpVe8Ugfw12e5zNq0gHlGdNkYXC1BjgLEA
qLuKS88mL4UEffKVaGZztTmhXQQYNznU0CV6tfryRC7nCesTso+9cXKTXM8+FY2cw/zph2BmsVAc
aXiD40dzDgA8sw30++dobYIFHVHHLaX8KBSmnaAnwmGXWSOWIR6SZWoQuAD87N7oKQcmCo/zyRKj
pCu98t+O+0/5IBX1K/UjKl3Crbz9z5zUhjM9uEKZwOq9AoIwbBigsJYq9ECDuuIKjL0seynXj8ir
eT59LeD4oVpU2x2p282KGnNoOCkts6q8fbfYTGdiShi1rvmj4AxNadG7DcMC1yX5/pHWbUrzOVgT
SAaJlGfKdLbQyOn+83+SOBRM/APYnzAiYLrRp1Z5Gs/RcekByMAk29JALefp8dlVUSOjM4UlzSS7
MLF9G7/5VFTvK07f9mY8mOrB9WlNwpKfUUgmVgdW9V5sCPibFwBaJoO8367e6CDWsuvVKQvDf9s/
Llbgow+/ulbOogpY6Ich9/wxw9j42uXuxZIZHLEsOqzg3P7w4lYAtss2tZh2g9Qc8OJugAruIL3C
8TuZydjC+GImQQQ53cXxxw7v6UW2Z4Jhb7WsGcxxtvxHravrrND3gmLPciSatP9r6ckEeGv0bHL8
ehofKnxF+vkz4bD9c1eioERnsygAhnasa5OcI0CGPj/+CS2ZepV4biXLUX9sJgljG6gCN2aCkEQl
hGnlH8PZw6DvC5dkAXyRFkM8v069NutFvbgw/otg08FHlEpuE66LXgsDns/mIjabi/AGB7QSBa2X
YyFsOyCQr8w1k7Oslw8+mhN4gjFFbV5/kKJ6FpbyuTCJkx9ncED0X4UmkNDepiwlUFji+rG/tZOj
QzpZ00vCpz7tm8KWlcTj+AwGBgq0U6PqHJCOGjTtLCwibYwE9/UWh4cts2gsuv2DVaAQURAc7slI
cLNiO5Pi42a5mnIhljCdT1Vy8XHcEKCsYMqZCYimM5dj62AxBi5FW0VImCA4/DqFOqWX1ahUiLjl
30GSC4AWUrQB47Lk84QxPrQZxRuuMck+bPTQPMuVhA4yFwNuS7H574I/smLhi0V7TOdiVFC8EOyQ
QPUvFBkiZu96rjjZBszO3L/b6Ww2Kem/i46HVz8h2P5HzqFF0F37yNJpslD+LAJk/YgByPQaKd/S
YpFoQT0Z2fDLKN1MawXBJto4CW9Zvr1EAl9uRRMnHH1wYOQbXNdCuU7CgmvbLukOo6Qsp7jrgj1g
M01/ZC1zKxfTeCxiQlq5qpJe9UxlcB6xTq3yD0Z0kGTRX/L4y3nD7Yg55Nsuw8EFpXiXxZu+ij6S
MdJ6zT6ylZSLP7ydQ/K2JFcbl9fF2PWkiqihilld6f+9Vi44qzz3D2RXtSY8tCYY26tlVFwQ8nwX
uCG9bVYClC28z+/rHmKjSjWeI3e10Xf9AHYvV2urC9iT9/jKkygr/cFoReiieve+hD6obB10rs8E
osmJ2ybvj0OFVrzrc8PAEpuqcR5D3sfLGQ/6PLux79qHoufqX0RcF2zZiWS7np7A6Tn0LHO/L/ed
tNF8LKS8KkoffoY4qI94+0tdfxHt+Q6ReGi6KYm7/P9YKM8aSw/iGttHSVAJEijlgDKUoJaXFFTh
EEaRvOC91L6s77J8D51w4L/3nyzSluqczrvKkJB+u1z71gekxyIbTIxWDM+ihmjQFMk7lB9jp+6h
Mjdw4K1RnPdS8XFsPKOjDEfMXvQAEJ07NAd3tER+pf9X6hIB95DjrTxjJjXvev1z2ZlfszOEqPGN
TP7bgI98rxw/DbSCRWZ7dqriqCA0AKGaU8beTUZgVY1URFlrSkJ4s21B/k3TX1wmbTR2OjkhD6kV
XrAT/CfJLuX1ZTHA8FyCPLyr59YfzsDxCAxX9fVWzIXP3l57GD/tb6A7kIUQHio5cdINhWrpJ/ke
8xbhh+RFmcU41ZEgm5JYD0c8Id4OL8LJsoaX6L2MhoTIb3sV/XoZVLU2stxNNuxjhcLa39KHr13i
v+6/2W/ertvkffOLHz2Wo3pnPJ3eg5stjd/mihBq28tMtUsUKmAqjn+Hn3jE077WYkZb6+jUgmf7
SoCMyRCRs6XlqHaGg+F7C/bxZp/4/g8vvy7FF4tC0bRXtU0t1/ol/KOBngIUYjtzkXBJpPqOfjTJ
NsmgVqPLHn7o3p/XDQC57Po6szmItjqt3m2bL01iLKZojJnW3LrvgtH1kmSjwr6jvsPLNtYVAYVa
qg2QNwP4i2g7cu18Q6tzTO0KqyGu5D1ffsFBMgHtYUywR0s7KVWbd4hWSDX87KltExFU6lI6+wOe
lvPudc08vjLtZnY9h4tnZMNF15UP5z32NMBDLyXuyvAHOYSRfaxQZOXBQm0Fnzk3/jXjLaIKgyfk
EEAZ8UhZ9mpa0cGHFPfqEknGAqpCnSf1AAkqPAmP0GrSWONeqTR9tQVK5CjEkaNZag+vCBJIPmT1
ooVLVrs+yq4PK7g3yZUmwQc/7x/rS1gCr4JyHuNlpwrznyy8OsCMFgK0CFtBgQ7DEr8ZdIpvRskj
ZEXxRNMSdGOQlop+jgz7Wf4O3U/6wC70BM5B6Ktdtj5YBGS9AkbkXiNS9LJXtV37Ko96SXuLdPqw
xMV6RIzYuNjIUxex4nWBUlXQ8pRY6FjvhJrEAj093bLy+hJ11UuF2QRuVgzKWVRR8/PxE03IOvkl
pD8EArZpTtnnCXVd/VyS2xDyhVTmK5b6GINk6jcHfXhEmvOuGEcc9cKNnP7m2OLUnmUQ+ZNIt0GS
jbMxAojjz2tZR8I7TTBAClUP8f/PU145U7SKAsaWHVlxGGNzuo1kYsluYc4wY31nbjzQf/X1OJor
MQv50CpuXZCdIJ+r90t2iwdjAdE8GKMAnLXSfuwctDyYppua5vEC7e25Wm5TxCkEjaABdDgiXFnN
LvZbj5A9zbgPekNPTbiepdHvp86IkRBjbmEDutWcm8SwdCdTUFJFvg+dY1048b8+n3Q69dh244i5
Tlthg8a3w5H89xSa1Fu7QWvzoMppqa/hP+WD6zhlTyb58fAgWN2E3V5XbWy9SEuIdFX75ruQA0tj
wd2pKPrPqtjlXo5nblzYxqGnVPi3tzUpQ8ue1eouvEKJ3VKBadscjNXcv0F24tfFNMX9H39IuHyi
HW4E9P2gtif3HEz0BHtrpBcEfwt9y1E0ApM8IHWca0RfN6mT0DSt+JA1soSqDn2AVI5OM180OQJS
JU3Tdw2R5aO+dBU4jzdnzHGLYEFTUh/t+4b4YfbcabJSQrK6ZB9PVpLr0+zVf+menJpSfERdECGn
BYAbH0lpWYwZfKO3Q5X6NDzFyN5yM1zviv4qDIBPuWk68jphB1RSLQkgkA9lFzKvyCxIgJdSZ3QD
H3PIarkggmXMNiNtRlYIg/Ea+X9WiaSAe5aN1XGS56Fy4rNkmmlqiWjBFKfk0i3NKxPuApEATvW4
gX3+8rB0hoFLSdI1q9UbJgkt7V6pqde6Q6ugQSlDy8kpGCiXm0lbbZRQ5zHRPLuT6SG7X4FIkStF
8GEdXkKAHNxjKBX2e78r0Vx3INDh5DZwplhcpgM56sc0Ja7K/i5+Q4el3B9Y/BwlZ4VL2/Zvam3+
T0sORV31apWh6lNG6MLIhGzfkII2zOf3By47LZwmsb/ALxeLbrF3/LOfI2MDRs6gGWRThZJClkzk
hTIc4EahpzcmZwv2YJra13NBwayjI9DvDQ5IhPG70pmyDIHGiLyiJOMF0INP0K/liQ03CttJ9JHF
Z3FNfGYpve2DnfpEbe2mKLktDwFBA+tT+gJoapQvTBwMZf3/6PRcAvSylGsbsYndPb/pwPnvoC8o
NdcnI49Flx3bEq5D+dLhJwdkMWqoOs1gf2Q0O4CSgxusCh3Y8OpGfvGR+VkkQ7pET6EjUq1V48d7
ZAMArJJqHQdBeLl+sIJWeKE9ZGAj1IKKnpRPKId1foxh3/1GTuEbx7lBI91y1dUxTdbpP/ON8O5v
EsG/cyAOIlVudlYcZaJLqaoA5ScDVa0IEVJW7aM7EB8eBB+EMqwSzynR5/Hm4H0QJnEH0yMGsPiO
Z90HznF7XQsnfdVKSg7gi6EIJ2Z32Ld2Sg6mZ3laepxREC+x8yfO7FciNZmTTD9qG9Z5Y1mzJas8
g/U26Ud0KOOn7PNDQXnSVMv2wleleGoqBpMMKA3VkM8AgNm2NO89ZsmulQyvKjTOwJyPjju7FDFw
YPeywaI5FYanuBQTQ8EUz3oukItwFCGcvEShI/RI5lvNrhJouqU3pNmOha+P7NH2MpSn/QDOw6Zd
2tPQxLtg4SghDlMZByX1G3erEWwYG3xCRYll+so5brYBgRjOsXNDD+veUYjsG0jNdVRfuh8AP3oO
8Q+o5kpw28rPk5F7k0E0Dlr4M9Vr4ZBtTrVlv710SqOGIHtZPZ4+sr4ahYyp2vx8yg7DnD8+O0AB
krIkktFYrpkdBZUmfxhqoxu2JsFiTfdjCLTrdDY6KHHFczmBefBLKG+xs2oemzvwPfRXT4AhDFYL
3zQHHObiR+pBYiOm8Vg9wsrNAeCUaH3qTrIorJNDIq2ZI9qdzs1rZQNrJLzSTE6XPJLFNMQ0Ywst
SuZ9dupZd2d+IAxGIoqb0QwogpP/04vl9/pMP0rODlwnbIS9/rBYoVCKRqzSURGiYpCYfBILw8NW
ZkeyYeca5NLepoe8GdRE8uEJsdwwGNc/tLe7nFIGU7kHkGO9jq1fzQPgQ9FeCeIa4vFJs8qEhcno
WUQrEPhWCgDcbrnX1aRLXhmTC9R+doyAH6ns2i8kqZ+TzNDALhb/5FYfj+LywrC/TrgyT1MC5OCy
r/OaU++nJ9qhNsZlDK+W+8QdtCzTYCyWJGlZbZrW8NrF8Z2L313vvkiZR1d/o8TP2uCHFJGxEnCH
PkyL8QDizNZKbclYeAHqg1QoV69vSARDYRskEFuzB75z+7Fog407J3SH0dZ0JedW6t7FIad80TZF
8UV75f+t4KEOQTEB/kmE0DIebp8ddXj6BlXIaCnGA06RoqDLzUNKEPTvuex5zGbiMPL9LObXA2Ut
2BvNgeIf8oshJuZKiR/6vk2tK/yHzdIXfC4urQPf6qJDnIL2QEwkQ7dcP7NYjDdmEHrfXArKPXqM
xJ7dyy6n9/U73V1ZE4DhCGoBX4XJeDjHk8AJqZmsaR/S3yWjKYm5IGOCZAdCy6N3vGCge8kKyItI
9Zzh6GfLD6k6fxPw1vq5EDNVSlV6IAYc1vRWZ54ldUFD+GwK55bvyH5yoLw8n4C9c4lZuxmh/KwK
s3p2qd/RswrrZjEkzbiX8D8dvHczo+SEu7AANfVFvoDQBfkN0Br4Wx0Y8/yjKYvvh26iFmucrNpF
gtuC9ofqHECptgr2+HKkpQPvfW7Bymdw/EN7cJ11SYr5i/A/u2dCiBhYJcnI2n7BAsaX3VQ4kLG4
7BmpTfemkZhs7KDKR4KREL4Kh54GLIUcYYZuf3yf31swOSGwadAgbFa8FU0fsUU5lYDSModg9VYD
nTmUqEltotGjD5UZ6ALipk8MlVaxWF7/d1P4bC4XpT1d3oFpVv9BxfvYWHjDBsJxxgDe1PgwEVed
/bgnVhX4Tj0+JIdorurCTqoLJhj38/SC39RmmRLfQykn9ozlJljyeRC1zrlYjMxhzCcSFQbMrtxH
zmOOQ3dp4K/nAEr7OLWxKIc8IyY1dCLvYxkSpbEhZb/eRkVngObv4gQjcu8HV9sMfkh5SnBZg8tb
pRvobx7KHvd2qYYqpriPIrEDs7krse03YeFh7MFftsrHB0b0mXKRqaf+KfHn9HGnUsXxq5uPWV8H
gl2LNOvjL/3pxlUzgjCtptR2u06+q6ybgFNu4rvlEcps3iuMCOrfxpbxj5q/9jh9Kkgo7GbCjehB
F2AK+meCMb+6AUIrWmwfrsmeuVPiW2UGpPofpDkTya6itDNtNMdrkik4IFjCEIPdIu60MWv15iRL
ISUCgOYzCB+6n/AsPfk4Acr0b//ZIdJzPllfAg7Fxu/FmLOyujLiIoaKmRGjmtXzo4wAsE4lVYSt
aX+0E9uFMregRosah+N3A7dLt7jC92Fn2Uvzr90zPDWYnmL6L7bp34kXzmtd5HunGiZIZb73BHAq
c3pdxGr8l90akHldVWLhQ5uQF0veit8fB0YuJGayQ/V1J8EoL1Oa7BxkcViflIp2WKfGqmPYwHRg
M5P3u99uFoJ8uKa71yJitTi1mhqV7GHgUEaA93+bk1EbAlCXhechixm2ZQQ4Z4rpq/FjaDA9iqab
d8khfboz+XznHQdUFycbRQreeijgqr9QScRyNgLzzvdW3MikGi/tmq5ySwbKDJYLk0Gw+Jwr3loL
17z79pDj3SA/r38JMrT8/hKNEShKOKhVXAOmnxGMsjtgxt1sC7alcKfbpV+zlgqyyOAZn93qePup
mwIhso+0N1WJGnZWYftYzYL5hvNykf0RGkdo1q8Lato8bYTwVe01DPR1iTqZrK93TISOxA5TDvVq
4MutD0djsLhiMsYw1SBSyHgmbb7CkSOGbiH8ZV8DA7Q8DR6MrQcgzZ4SHrIlU2braDRUH/NtqFqv
0zXCHzbFndkalyUOA9WNdaofkDIYfcdMJhhPd5k+J/8kYR7Cp41r93B6fj8XGrn4e8D/mRdbum9Y
HShF2BxpRstECk/Wbo3+3OU3HqAVvh1SpmS7m37mIUBT3QdsXF86cluQL66omyq7VB3K5Ey2uh+/
bOu8UJKcf+cCsLXv2DYs1db7uqkfEKQihIlYvmSyTVLNg/W5t2Wm5a03HdVyltlIVXW/DQHa1xZL
HFeopS8RAU/5MLacWOCRmyhyU0rCgijq+CzJ0izoh+a5bQsRx8/RgWYT+rP/BrojpU6A+kRiXziu
Qhf3UNvEW916G8pwQo6dSNIBeSOIPiwWi1sxwMIO+swlKRdxneDp6+NhdOcD61ler0YB4CbQeq8S
pJ+OyxkU+FIq/HkH4vV2e7qg4z0AOHqMcSqkXisOI9zWneYHzIuInN2NzdDfLFkcnw5u+nDusCBU
UL+IZP6FsbDwXaVu5wbsvGN0h1Ipl7eo0lgBNXqUpWp/HYqEUBAFOUsQPdVI1N2hZn3mFAoevt2C
76kJ295y3Uo4EjUsmNE3VyzuWBplmdCan1VkavopqfvOfdWfnMJFa9RfdWwIEB6h9+LqWBvbooae
ZqoTckJ3Dwq1FCuQm8PZuDFpvEoKxD7Z4RAnfOlNgihswAGnvgkn4NqLahOmUEjMxfBQRmbH0j2d
SFIbTaQ6g4t7NMIqIyuwEivnVkPh5yZq6AmnboDHhM/BNF9rYnOHcodCdou56RVRkDmulYOfUYZO
sm3RIgohTGqXoH/2EmezWUrJa3vdeWotGYxoTJEXcitV9e1S3PTbPFwJLZOc1bOyDfNZJojsMuiM
tszLsZ8ghy6cygWMpvNA2/SPd8woE+M5lFcVi+FrLp0TKfR90H+iI02xOIuKB5RLOote0/igfjnP
SSuLx9xMHFFktSsTyxYw7HNQ8MpWTNzlvOYcFhntP2Frm/ajLs7Q8P4YMUOTB4dl3jdskt1MT55Q
kIMNE6th4H28xFqkuHwoTwPYFGybAbW01cZyxLeViRCR+cVmFA4DgGtcQwL3WD9YEaZLvVUt7ef+
YIJtHZelLiKZCGOWp50zqczX+/2FROm5Fs7czy77/4wIaUgpiZX6SgW5GKnlqBa19X5H+uT4oafg
TGIFngW5pmXihSQZxblgN/SR5/4+t2JKISTVh7yros/5OXYDAfcGQz2vX/IQ4AU3Ip2XmiERovDf
8CVla+1WSbqwqazxCxpReO0eQYi9Pg3OLFtzY7mnDR6u8qZbfvATXp/ip50O/Wfj/A4ASKfr5AKY
FaeordWb/VEV1NAAD7OAYj3bMdcG10CosTVihG4vOUMHV3Bk7xr6roUipAtK++N1Hoa/2m7BdnMT
0xjxHS2iBIdcxj2ZkENT6/pt19Emru5Sf25Lm6v4it4zo5zNJdEGrGfPXJMw/ZmB/GX1otYkjGUJ
/GsQVXD6s0JlNHQUp0XTSc9IXkuzWP+iNy0TvEh6dmgGinkS2Ie74bAq3wa7zJY4eoRXb38Z0ecL
n7zBWXLTZv0VBVczcR3Hb1E7NNkUS5N85HWhXhRWbDS1tAFfOOBWomBxPPtOjctVEkS2CmJHjsnW
NZxCHifdiW/XHFwktPlImFQD0FwX+c0vsLdmxBk9N8O4Z+pxIcsVxHaYc0oGmb5sc6iyqD4ZdH9n
DbGMUF7lZqmFmf884pObgZhSgD7orVthO/030s0/WolOy3Q6T3MO8Lf9hv5w1vQJON4j07HtUbDe
EFwyKQWInjqLzO/9LvSWdmnVHuGiVITWvzQ34XIQ3O8FHd3w8KyruUUI1BHvZooXPF/K8P/3bq+O
zlArYAstUcv9pHkvilEmETzqSLI7hEDmhospILvbQE9x1rzqWs7vAnv7VAf3vLEj7CYEEniQd3AA
o7Y3zy3ItrWCy36AdtkfFZwCrSjzl9WibcVu7yy6zAUph/zJRpxQios1sMaAc8wv6YK5SS4BFl2x
KCE2AVXBr5Exzqi1ud2PRBkgA7tBKhH4xXTEUoQg+tk2sI+ORx/OdtdFSqoHUHbTF3o6Azr1q4sX
Xq6aqWYNnbAwU5bwH+fy86a9dPRzmvvg2C50Ok8z0wNKkeMHKMn2/K17Ahkx923m7eUhkDDThgCX
FRqBwT9fzT25ae7plImSFvlO6Edi6uqfFs/lk3FR/i2LKwZtQs1paVEWbd7LKeEWvHyg7uxUyXu1
oZRfqROQbMO+coGxf6Yax29AGtHqRF2GLHbo3pU6HIZr+f6wILN7UxT2ld8P+qY0WAzIMktfx2oC
ZWrbUDvKqSCtU47BeHBKXXlTY15AHiNYPuq+RGoXHPTD+2sKBqONufkCqyVcSeZpRPjkNkpBHd82
ha+Mo4Iy++OY0Q+TnX9+p6yiE1+N2d0iKCa13jnwfTL2hOxRuU38bp3oEKDL9Od8HH2iH9/Dy4pU
D5RUiTtZhwXs6DbFg3AJkBzFSU4zb+nJ/zpxPtoCStsQebIhD5JknBozkuQYj6z6k/C4kRJaUzMK
O23Ti3/tu1JJp/w6nZaImtuEhLOH65Ssmgj8MTVWZiwb+giOYRq/JEUoG+lDys83fw+AiMPSvki7
kLzkCkgStw6YFcabIom7fgyFoGSMK6mikguU4LL9886XXEDhXmIh3iggiptp6KGUxTKxFohm3orJ
Y7/JUgjIxQ1CGF97t1ptb1icRQ9OnrPuoEkQlZrYWVavh5Vporjq1L8gKZAEWJi9zOT/J6/v4Tdn
LDcfCo1MFk78L1kLCZbiwCsNrlb1jg9wqZb35WLMYLVy5X0hp5E3/DUGeIiCPXzpm2YbQbelTBLL
fhASubvw4LT718niKTLrynT6UQ0IUfVTv8JdcUQyF2zkp84x4vct4U2/FYCD5NPjFE4i7g1xmhar
Olf0YTGRhoGJJFrnFerI7exmGQhXlMqYJODf8j8agElkd4a8l2yQ+2kd0BIw4ZDfTCC/huILk/Ud
j6yyyREJW/NeteB8RnORcJli6JSxoJM6YHkr1gt6ig/M8AJH0V0iKemfJyAI77QTJKVUus/LZVBi
4llV+ptBqNrz4GuXUEEusD2M+XtQkOVtUfo147Tr7Loy+fCXugICb1hZ5kjlrqSFsZAaLwBRUKUV
qus77a3gRNqN+479ilgLeu3b5m4asYVsPEqAp+TAW5QFVNofbZJQ+I9O6smRAcOn/aYGedPBM5xC
PHeM5MS6/78KyAwtfoxzAHpYGFCf4TeNlC/VBCPLVOsBeIv9/gU85rTYVahtB9aVi+XPF+tyzJBD
F16vXiGyjui84pOU43elrn0vhsIEko6Y43/g3Le3Si1FnbmzQn4mUkfrA9wU5kmaJ/zmlgKR3ajs
yR5yF8fCkmDzb2S/I1PMtOCkVXo2phjKuCBXORIBgmQT4Kv2piHjgmJAuwDwSXvmpUQDdORU16rq
6jn8OmLI3OPMCYjEK3Csu4GobmF8kyf/YdHEMmjQ/NUDfyL7jBBZReExjHCz7YR5Xr4IBl8JMZdq
hA/4x/RAv3CBE2isokXOHVZrfmA3KWZmU+4OcWT94BEl+g4nxXkxkgaBuFKWG1h/G/gZros87miV
tqdREEWIgR22k7g079E/KxlfIPy4XUj9lEvN24QGGvrm5nb4fVVd4x3uEq9v5XlZaXNBfehuo/rq
uR/hh+FgOetinYK0QfOaF0gN/XQ8k1QBQ6CEDgo2qGsUNePxB3UxxKkpOi+n+ZU841HgydA0dXTt
TM8sOyEUjJz9yc6GhX8vMiJKjJSLpLrx8Dy7W32f6BVrB+W+i9R+t4PW7mWfrwFLfNLw+HRDUXFy
DmbBBHCqZK1ns1W2DyTXzqkZ0pzefXvqTy9AbPx8eeyUqW2Jai8qONiF1f94J+B5i9O84E3PmCax
A7ADcoREV7MT7fBaPVoAFsZPXrrRXCaQY5XiQa0nxveJgl55kj7b+dgwmdOtsDbUSMdnpq1GrC4t
XOe9021sKbzc0a/tYYZJBsKTU+KFqMzkDRGxkR/rU2MvwFX/GpNPSWlZrjlbif/vq4TpdU+DciBN
JPsutovqT3nUgfp4/nuMruobz/44FQM3zUSm1STA+P4zQpiG6CVl+mr9I81CeTvAVtymKrZ6V2+c
iqEB6V5y9cFPvRFi1qMFFBjprRaMfbYzRKh4rPNdwxtCUKZVNKK6qG9FmR570lE/2Qnz6Bp+eVNZ
WeI6CkVVT1ejeVRlyAfOkWTG71seZTn36WEflSpWghJ1vvaktce6paNNUzy5rNLkPJa0Mv/Atbqw
c+VOv+/ZZDMxiDtHOkl/C7WnsMQXDhDRFcTHbCUpPDaG2/ieOYupl1rGWfCQtDbcCd+VSVh9XSTQ
Ttju9bVCcziqDSMRukyFo5Lv7aIite8AyWeodHZ+1gUwF45r9TJpgkqDvP5pC9cKLFL6+yQzJFkA
2BGyeoeeECNJKhSPOgBSN/XEUtEHjV+50F/ekpypJbwpYm9DyGcXfxoFf37/8Pi2avZrCL1vwlar
Qp0pyQGFKlKeWxb04Tq8+/OOSwOXy3g9AYUYqWmC0snK004biHcFez9/6O+EHaPGevbs8sOThoM0
aVwUqjgkk12Dgd3jWLUlttuoWrFVlMLUVPD9Gu7MZYgPMUKvoYDbb3Qcu62wUtboAPSni51nXD9i
9cU2oCG7Qc9MhXejh1tC0b7k/xyesKMDBzC5rR0aX9gGiS45my0JQh7DvGO4M2bmK5s5T0LrKp4J
Qy2koCe1ZO+UlnS0yWsR5MmBxE6QbwxxNX4jfEC9U5nONnTXxizLudd39zDsa3S4C2cGVrNBrfSw
/nc/Iwsh8ofpS3R8Cppw50uGMhlAYIZTOjevNi6CQtTuGk74PxRnr9XCUu/2wtEjnKP2HOGTQlEU
DLY7N67lZ/+L4zXgEiyWIR79ArqHB/YArAt/1PQllPiqzHOhG5ZGGm5b+yK60M8weiXgGzsQgTvF
q4OzEMsfpGhiqu4dRZNghZfqjAwDxmUjslt72oJsI3Xgt2Y3jkTDm0hqh8InmyS9AyXERA3NrzBt
8HIXwFszkYcdYdgCvk0n1yhlhKk9K4uQnRvp+MUPBNpWiyTgihVSHNdeIFxNZHiggh0B4FKyMdym
TZ64f0YPXOBAxgbWh0gefDSBMEVgr1ex8qNeLnhXl3CAINM3I6jVnq3C69EqwgnBYOTqOFq82QSe
RlJMeXNtp4nZ67yqXHiGrBg7aEPBKO3UKk2H8TSPSImdff7q3YBTe6iy4fEpD/wvk3cXgJuculeO
UJaYQv3CPe0Sj0Bnw/7u/tWo+qjxsjjejXNtweF00T1LUSuV07qBVs4JOm2b1xkmCswnMVRjTtj5
sB3Yuj1raMOUqPfjzuP0FedTVjyrFwvbYgR7o8pk07i/akHdKzQ60FWev4zNCGIy5Bvgd0YmDgV+
O8XfMwCx1eAqV43+STm6Aqf2xGm+PVzpQ768QzvpghapiKQWLI0tPMT52AHm1WLuV83pwTbfuDM/
R7eY0B1P8Djur3G7OO8i2Hi5pe0Bi1Kkepw9+kT/AAHMrtCNOufqy0avrT3XZ5F9q5i+j0cQvoyN
WFUZF4bOxqvE4z+j1YXYSeVOWmNxjuN5SmbzrOcR8w27NMgITFsJcWzPI2HuD3yVV6rObap72x7+
oAWAK1JB7G2fmvyB+67nEmvCWfME2wRFmlOUIfX/cTxYg+tFZrmRt3XwGIm5zOiWc3bolj0PwCx7
n6p5/uOvzoAQrNsGpiCdWS3UPupu9FjEiXrk1ITdP+MFxiNjA0aFgvwCyYrzzS9Ra6vTi4ibhhN0
NlClPY8QMSjdWjS6D8YQX/ldVx6elF4WvX0ne2DYC+6PPoN+HXYo8YfrDXpvf0hgsOIdZB0svfke
STYi9tQ43MYEq2FSBEqSXdK1xHlbWegcOTljjiqaG/2H6LAIDCPhZNfvEzhuV9YJ8k/QsEvc8dOX
qX/r24zMDDMjzqoOJahdyQVxMEUqbbdAm17N5bSiedhiWSxdrSkZSGWg73iQMDs3jIh2JdxLtGYD
tLF1Ls4MhTM7JzFdqWTsbuJPE7LDdaRbNgPMzGaGBYx/8vEqaiZj3vI/xhQc0jl3LL8gJCqWACd4
45qA+Jy3RlpnqCyKGPRxtmv5ZwB9cCo/uEaRlG+N6PQJm4y4myNe0VLVT6VFxUg7eUa+lolMYacO
7gKWxvTUvLGT/6D1UL1Uy30ZEd638XrObjPkLnmd4hpsLfkDxvInFFVUO6SAxuiZT3otE74wYJF5
g/lqcm+FimeQLggdQMgJvQmsh1BvhYmFi28gcoHjXWE0lrz8QpfU+pjX0qzJ1L0Bd5sZ8gtYPQOF
hxghWU+UnTiPJ4OoIdiEzBofetrULhS29WYE0o4fQSrembzYSxhKnC7rvmSbtnh7X2DNRGGljT2O
VD27FIhK4hO+Y67xWkU/2PVtPyE5jWoNIjcGSHbl5JdtJENbxOgZ/aJsaLAOJ+eS6Lgo9u83RLqU
KvBBEKxebBqBSvXjvCZVoQ338atbWrl5hmBGSMZvsqIA5jHfdMTxQVcZdw88f7bFkBYK43sCmJ8B
jDkF8ODEKxDQLMV5pRWtBWJtEcfO+U3Y6cxMM0XnNhu4Q9Q/AK/LLu/qbUvFPL5oypP9rIIeO0nS
PamZ2R0d55tQTByXGrJG/lGyllNTNAgRO/W2qefMoHOREfbII48ATBHuGqUbTjQVQ1DtcsZNWGg7
1OX+9jOn4sCFskcKE9lV7i4WW677vGTX6berQzyOG2w527Y+4y369VTAz5rw+aBDhxeYH1NnUCGw
p1WSeyh/9Hhn+5Lu8Jz2I0Y01pdeT2070226Hyygg3GdcSOZGG3BtCzLPnFx+gfWCO16z8oAXQd6
FnrbFF5Eb7Wp8+3CQ4VhwF8AexynB2LnCLcUkIMdZtUgmEXAbe9RjIREf04CWFnfodNQqLAcJGgH
gID165oRn/eaPxhv//YYGkYyq9aJyGnN/GgZvMfdkdk/VGzWzGK8TQPomT+V9kvfOSKEoI+slV6a
9sE9HVwVBHXxWFKvg+hvIeHDNtNk4d0VaxdoqcY5oGsCNGqX2HIZUJFxe+O2XK81OyIPoLZny6F+
XR26ESHs/ESgl0uzViiwzzXxZ0kSn3jDrYQ4NQ5kOx2qkD1btJ2NW8oQ11TFhfEQgVdqtDBq0QHO
77tGvJqoeGJbLWDkJ+JMZWpeR/gZqRtfOHwLXQxp5QWCS0i6jJU+It4o6ln8GxbFK0JIv6s8TMW9
YMm5bUWTZLslK8a58nqgRczSpdLF8bI2Uaq7bbvpP4FxJcboINXdppkvi6/zf/C9QVxy2urbiz7s
xR6+KF2FGhYMPYEsSokz1LH7aFQotTzOnS4r0Aw5QCPtgX1LBKkyAWgIYjiyQXEYqeg7ErXyP/Rh
ukqJX0ia55dabZVqE6T38Zx5q5wEuM+MEH8VcmNOGmkrSYr5mgtMCMISmndwi32ikejzud0wvxaN
VbiGL4eovx9YNRz5K3VnwhSrg8wnvPhO+FfeE+A4dBcTfw4+lm1gqTTlhZMvljrEnwTDFT1hYD9o
6uTWHBN3Z5K/lPDxFIO6P2FPp4y73mlxotMgGak8ulArp1f71gcUinHcRZXS8yMlpNssJPj/mtks
Z72AP5lgwQZbYMrsp50h2lDAzNLYPToZU64ATWbRIGXwVc+t9SxzvZMfa++Fkvw4OREKEqbZbwOA
AgJqOvaNVbT2YyuW3hIWmc1ed7VlpYLXWTWGSckq3RnkCeB9tury0eIZjCGRsxczelX+l0LiVMv0
I7h4qnbTYVLbqrRnQgUfqDfkk4tit1N99kmlM9LK2/VZuRJ0aedWcZLzgQHMDgjKTZBIpGedE3gn
pPJtMhapddX17gqhAJmzEFu42Tdimv6GxRUcXza36NKdVFEZuRAKiMEiiGn5mxs6jv71bboOgMej
OJSbpeQi1j0YTpzkIGAvCWG/Rb2D57MfOMRNsqKhSOpitnpDPUF0IRR1Ch9C3PDGrCCGKA2FzWSM
NZ2BYZrBjsGOHZj3dq2kA1F2I9w1kUFrsYR+X//NY8LtbVpCetT39mS/EFFH6oL3FkWZZAnw7hSF
MlKqgeV2FREeovJJQ2cYILCjak/d4ZEFYw/riJ1lXRV/3Mei0HcXjpJ53bL2+3HARZh6O3BZvJNq
reWeaJ9ZzJPTGBO80QBjKiS/7Uh0jW4I3PmEiaQiINbq+ujKjMF+PvsNDU6WIOqXb0fgoy1Hnrc/
KI9I3SaLcBlaUbz8QoYH2WTuXjYctCz0rQ7KPhlw2RT4sxF/dzidxCfDwsjUr3x6zOmq6ttSm02b
sZKOtXPurJy/tUIYeWkj7TOzLWMA7wUi9ycNpZ13ZrihEq37h7z8SDqvlfAH3V9PiTTAWc9artMk
hxG7Idy5YDULy5MQKJDCTa2OWnWMGPmzBWKHfhW+J2ZXowRKMPZKDG9YNvt+YRGfY8rnuA5EQsCf
QhLHhEothI09wpbswi+HTL/2ZvbsbweRjgrB4njrErj0z9cMGwrEXTDI7KXnnHXQCL4SgG9EVnpH
mX3EQbsJgEpFHmYkdVm3ModIIx3/KKVpR2gidrsDDI5ejHN+nK/QUT3ITsOKFBiu0elXprlmsi6/
zfftGXTzHXg2zTQ3DHu5az0YxT0Yk38ea9zBoi+lUU7TqK+R5Rlimpj38M3mRM9nNFTRnYaOVK3v
rYM9zt7koCtmF9k0Ia8xIG+J41PIkYXBRGXkzNwKVZkuZ4Py/pchCjOU+H31TYTGM4vJkDK5JSI7
z6VVHty5PdTHgeqCSqwmOi+HNfAkzN4g+dqW/NNyTQ0+GxW7l/hzf0gKQBWR9eF5rbI0KIlYq2S7
2ZRunSH+PgMRDayaJLA1Qf76h04ZQnIk78ufiR0s4ft6pM2ows5Cjfuwffhdxwh9Z1hqZmkSka1z
WlJFrnHj7F22FVcdQY1GXDl/6F6YokY4IxJi1EaDiCTxBH9hkeQbqSNeRtPqUllgV0Y1Vcv7jlas
N74pML/IaZ7CqoKhzEp6AaDDvX5FlW+a+aG6lMfJePkzpf2h49OxV4bM5DztyV5WQk0q24iSDNwv
JGjCxOwnyCqZuBRikwE0t+WA0lXsNvCOw7dkNb+NNSt26J4PHQZWKnhdsWWa355iCMKA9t4KulgO
gIGkJAQCw9zXiomY3FcZYlMCJsKMN8CICYAql4Edb6MzxAsv1tmPWDuHsO2+aF3NNEfMfftb9IK5
4oynsVeKX7mBayT3PiIwet6pSQY9TLFWQZ1ROPpqiXKmrHQ3ucWiq0v7i8jZjZdI1JbkO0qvSUqx
6CzyLeziWLO8Oe6DaI/+p16rEQBsCvsYxyQaKG9k4f+k708jh+d5/pVs1IANd5qdLBZ9T67bTLYE
toT53Y4uhxUhqLgd0eDmGV0/gpOBDXthHh84sRZzoYLHMp96ts0jbM1A5dNVvW3yKlwFAMdJXkRn
ESBcNmVzw6z9IHnDZ3zy8XrBHWcAS7igWwu6EAn28Wh35KW1vN94/PQVzXdA9qgncVXQLbHv8SzP
HQJrSgskC4sP655z4jr9nHqPSRqhRaGAzPBcrrORk2R0ByVM5bi8Pedekm8H90DxVEwagPPT1TFw
NQoXKmMQYJ8ifyfTNU4ueLecTiz/BVytRb/bKmdkqZ6gMc9F5FtTj2jc+IhjrcMPSpabfUeeznf4
c11xWZAdWMumQbqycwK57lLZB3zbqoek0RKzu/xR51HG254WYfeoTHPmV8LfWP+99ZdMRCKKOec3
KJNJW9HT3Bf5y37RHO757CYcdkEe6BEY12rAgIDMz3699TKmUjr9fQHvuGbSAGWGyWkt13C0ZNLf
pKBqKApFc/VQZdSfuicEuvsnk+97qGJlin4AM/DC5Zy4pJd8iOJIlZb6Xy813GChFDOwoQ8rl75N
vRpgzuDFNC2omCI5E6FG0uBW2p2OeqRrUSk7QcjOwYYOYSkPMicXNZKuf3zzXM0ABlY9wJVF9fac
mAUqzy2DzPgLLf653I1luXofoAQw36kMdmWlbHLXoOxNyMk+SLgNbcT7ixX2NpH3wJZM45x/IbE2
T0XIdIMBByb8cLrnWvXpxVAEjw7KPtUr7bVUtICuzP5jlMlXD+foivsCuqW3dwlmARYdazCpcilE
H3UG2m7BzotzZPFj8UYw7Mf0HbISO6l8qnivL3QRLj2A2TpdOxIdftK7I2xS3dL9pgJvs1mwD6BR
oyKAXxmcKWoqvxe5wj3+zFtKSRgwtn28H54LTmwqJq56JPuSpVMkGTgjA6tqRtkhlir8I0zX4cIF
I11AtqllmGnPNTW0CM1l8wDjSyDDBcSFcx06EKL/kDYUF7bVMcrvAt34DPZrAcK0+jGQMDrkO7Gc
mxcUpf6jFUMmAhnGeU3T9DBVQZHjOmID0uEfRWJ5H5w41lkwksXvs+3S6zVp9v7pVGz5SKWAezxe
X719YCPE7beAcLc4eH+FiST8jS5my1YdDA3hR43CLovk/WpQXc8T62FnqqhleCOB7mXXNu9PrPA2
4r1KuXMJgMpoj9UXJaxvotoc1soVNJCENi8XFN0vZW+oHakRg2dNDr0vbQR5QtDHpOyvgKAJl8iD
gx2xfYnD/SFTM4pvEL7dF9ACBQehK/D8u3reBu+IzGyi8Mlg96ORK/766Xn6/zTIyIVztD3wlaBB
iU7syirLD+wSELWCFsPoNdPLQytfwe+X9A8WGo1+asGMvXaT97dCmse6VZqsUGso3Vqnfr6f/ieQ
U7xvxCV/nVq7L9pDqI5R8r2DzFLsLlM8GMERMYSuZCHbvv9pWl4LSvM+xRPQEbL9BtFrcJGQjLUa
gxDhs+oudinV8IXU69KMnWlPLBsTlUQ3IOUYoKYX9o8QXQRi0rw4E+mish9LAZ9tEYMfrzZJP6d0
7Lf5ZBLV3mf28h7xkIULdCtGYU6HiF6ma60CJvz40kvzPgu3tC+vHp97Vl1z/yTQ5+RDit30+ghR
tvDWh/h52hWbRLdeoipuaePjv07XEZnsAFYSBM5Fqgn54Ce3bbVH79EGLHAELrq+J+u4i/rPxOGI
hOB/jRseto3aEIxYo1gi8G6CEBOYZdssnQ6YdaDkqUhJzsn/26M7LM4wIqAcEI6CCjaJ3LgcbwTG
2ncIp77PmlhsnUmP37R8NeL5TOCVG/xa9L/F8+zMR1tesgd5nJw883vBZPh7OOaMDVBxqTlyttFy
UqTyEfTOtfz/e4ZPH/I1fnJpySsnfz8quB846imMGDszz9ZJUXeAdrjWj+vd2m85MhlReTw0CrFV
wqsK9gVqVHBNAfknP32jO4pZhpBc0i0NGgkfgQBSstA2dDYz9DeqJbdpxpPnEdONfzI5rrDeMNZu
SQCFRt6wxmQUbCzc/7Gqyec0sA1GOOnRdyk4H7ZArd+4N/LriGytC0WUgXMGoTMxwhCuGeCGDjwD
oPvySClgh6GC2hNpeBR6q0358PlrdkrCaoaHFTfQX5llJ0k4vy6x+G9kzN96kQ89TZmIKe8tIxdR
Nc2hutNIYS1BwhbqJ8VZFxlrk2lj1/Z1IJY5viQ8Y3dd4Xhvi1YkiMkrOBci1RmkHhxG6mlo1OZH
fPXb4eghViiwzAub98RHno+Vn9k7qWe1/tWjgjdk0TgJ33v+gP8CT+Gzyw0FnavG+acce+vCuB0F
iZSqUr8tqYpSx7nBNqL7SWZsWx0u6Yk0AZUglPO6T0wfZ82Et6YEPMLn/sIIXihUq7UowpuTk+OK
M3PDZVqqVN6v/RY4p+MYBPy/MxUQBhTjVVHeUp+7Vzz0sA2NHQWZnGSTdqcpT97f/jWTY6RNyIo3
CjTIlreEJnQVwsr+1OMy/Y8A8D6iGYF10MDxtzBfeAVtiQdLU90sAxTWGGE4VTr40Yx81VJbjkL7
XHUFSn6vR8fPJmZOjVn2f8hPQ/oV5eQtFxY8976XERKhFYEno5cbkZ40uF9KcFAuwIdGtYocADu3
u/0V7qPHz6VgF5VLQ3YMv1JLNPsl+l1s+3NCUWi5VBOzrvfy6QCdIOe0A+DuYVjkgywqujQOlxLW
LvNCcu6G3vt4iPh0EEXluZkYPavrWSsv2Wn1q80gpyTyBincAElUy2hdJ1WUsZxuC41d5I7phLjc
O7lhtoxBfrH1bP6MVkfCVfNSa6w6BN92L2ZKsW+WorOxa+kV00vNMAF8T8o56Zf+8HtN0ePq3Zaf
UWqsFYZQiQUtWQi5XZP8B6UefNQzv1DtWfNuqVbs5xH5hX9WVpfpXafoi83Q/ctMqyh6tRSMCfoF
BpVt2Yp13S6dhmaDxaElxV60odlpX75fRkz5Dqp8Xt16gYzywgAQL5PguyOU4dLqdcuzaeph8bak
MXfrTat4ZB0LbHBA2ewUsYhWA8Aw0SV5c1oTtEPPcLjAmx1UXkStDeuujXEGTHtcDiZ3nIwr66bD
4Hi6Wj5sR0Q22Ew+OkcXYDQEhZqHIL1vSgYkvScJycG0jBQOJlECKZ38z6SHDhXTpVVWVEYr6l/N
99LaxVaZOiQS+UPI7iOlZG7FRLafB+TFsd7HYJWWIftU2WDsR0B8fqvJDJWFHHRVCY0P3bydQIrN
tWYfl64S6BuoZBSmGNo6coLNOZsMhEYHipnyahMAxnpgtLHdOmFVHPr3iVClMBhJw7yaniydmrq/
Fso4oQpGNZB5eqtlwTjvqaiv8qpMb9uxjrxEbO2iMq3018nm9R0OMYb41A/w0THgk+aUJsNYtcR0
iVEXLQ8MzNWVZwZ1cZiBU+T6SRytwpJPXGyailOUxhXpNeerxAo3/EDNam/m9INIB8tMsGOjIPxB
s0IjIl9Mm9T5/8KlgHR4vhe8m3WyOwZYTK2GjuXOfnzF3P0Y9d6r5ubQUvxAI2m92q6jVXOCDGQp
YdyHkkas4sMNKz3K1EEx/Lmag0BqD97t20NY6PWfWIoHVszoO+wXe+LzO1+FeNeDzfoOE/rHj6MC
Xeleqf2GiMWE4fJPE63odogOUcKX1VJhEa+2cgpjwY2T3BYI0WrYbd0bPh4InqJGXFhQrEHaNraM
dZtkEDcKhRERpTL0Mp97Cn0GvsEBR3IKMgGXD0hZvLRtuRAH4Z5l5dVUrXhnzzxsefp8hFyrom5x
ylVZPcqj/0fMfGvz2PjcY4ML3NFqMrCZon1RstPp1BAXzr2a2RdXV0SkB/a+PAKhUpB3C2D4aM39
S4M5wfk+Lnc+TDWQeQkD3Q+9ECLzoFYJ2iwOrQA4A6iTiIRkOd6WVmvdSIGemPrje2fDsgrFV7CF
awrTwsueaGRaWdYpaPkYFhugroFPXJtS6kP7SlAz5IvSBAo4q0JzwSym/y+F5nQ3G3p0wN/PUl67
zT1HnUwcUeI615zADr5Sz773oKsqoj9I345a8b05yyStT/9FLK6jThT7COFRMgfi4a/jWGZ3Wxmw
awulUAPt52fWxPcugcfoB7gWGmcJepXwVDeR00npbaAfvcVkSPHJG316vZt0sGoTAGRDybpGOQT2
BToUKAUMOw5AOq9wZf+XiHCIrw20maQFga/tSJvr8y6zL2vf5Z21oPbSn3OM4LL3Iy8WG37jZ0Kq
7wsuOHfIytiSV3/bQgRyI1eNVjWwmBk51eXl5rroLZGj8IrepJ01mGX+LXk7+doa/2rap6V9+O8e
VCk+DgiLVBgGp1KCn51XwJpcQxj7+jEbQTBtrRskMflFF51OM3upgXPdyQscmc70omBPCPrtz3tN
bh6StzM0fuE1j2xZSfg796pq0HfB+xrNnbFmSvot60QUOIyaGvvm4pdGKflebJJ38mjkbalOEhSe
n1TceLYJztneC2Rdr4/rE1JXmll+0ehD5UAG37mvrNwAiBkmfEtDMqeJIsl9EGa6H7hlgeSXAPB7
SVerqMqibYa9P/EOVChl8W1h8E7dd5gcYrFfjef+qrJs4kUYdPQWvj++NvZl1fKSuDKW6/W+/FrL
cJjQ/exiXRjOjSISrFEEjKGB0t8s/RraggNs8zhn58WRFKHsRez1A6UKY9h2Xj5HM9Y69JWHkdJs
hxmaMWMLuz0q/wxiJAKnbq/GbL+SVshSPfUY6bOEijRPvXNZWAIHp+YOFUGDC7gJFlSoOq+VDkk4
n9xN3hTDBgDkXMdvQZnGVpSaERsOKIo2/7onbKmO7WgcaAPSX2zNsrND4AmRBbz44rrAqYRV0tkb
DYdOjAJEbFV8Qj2Cy8IkOjH3V96UnMk9VEYNiqN/ak4tLibPnX5jxbGc0gtbJZzTKNQfpk9KeaY2
+mDw0y5sC9JW9zdbQhQEmywq51NGrjKoxv2BiEmgWzSbPmmDWpa4RHoS8pSNpJ8QDfh/e4ERTBNi
gRSqR8iOc/Yc96b0r5KSXqpOFcV+j58DQZXQDqWjch+7IKZLZRKi+qz2YMFvtsYBA0/sgMNK55ez
remr1fi7JpVS20TZPXrq3qeYIcvnaN6uYK6TlzxoDYdNK0VZDxGdtxv1JFjuZRhgsJmdDCjEPz31
KKmAM9iRZTPwWqpTHmFOD1BCW5vv5x14WvK+JXJnVDKp2nMa5ot+G/j0y2jeMEJLXMuCZBpQ6NuX
slSgqnX/JavmB82oYMFT2nG5HIgReMpHrPY32rDZNueiU9vnxu2Ai1or77+zAJvtF8FMlDJ73mLL
C3xJO3bMUrAAzUGVVGKwconxLvqyTTjv2uC6YKh2KPzxpBhPGXZ6vaBIY9GzyMQWxINCqbzqDyAz
31pfgtI4TyMbt5DJGtiz5C15oqRAhUkOhHHsbglM+WmNX9uOcMy1bdech8PR8piRUT5PfNXakcwL
zOpXZd+QZd+Tmutua6brl7mfsO5BwZrDCiXiWtJDJlFzVbSp77dw1X+fcm2SZAvjSOXQGI/MH4fq
D+lP/GWAQsy0/t/1Bfpd3GouDeUiKdZGfL6Q8m9OAwRtT68NREfBtGU/ScXnL0ZcMQx84U3pefSP
2hIRqsYvEvmtcGd+DHEBCFWkJ16kcUVp/K4NezL4GUhj2IAfi817kW6ZnDpP0P8Gra7pBQGcIFi8
JdsE7JrSIyEctrzYK4RYBZE2msSVa9QNAPNZiOT0GIE6f87SNw6K7qypsl0lwGfuSX3eD8Jior9K
B4RmxinpQ2EW0ObrgP3uknePk0ASXQ71GJnincwJeRaHWWw3UrOkxblpn1oqHQ03FGe3tAz4mbvy
6ruOk+yGmHaADhfg9D2S1OwVHhOskVNolEEsekVvHIQbiVEKJlzZc8fRz134u+7Cit6YgDE9OCkl
q4bEkDmOUJ4KCa4kEsBL5RkhavXW+VflP7Eq524oLoJrbMVb321JQlz0pQkNTer/O8NMXx2Xso3t
sNwCpUUp/li9gLvCyaQsmeWwP6Wvme8ftGdfLNqMgFNOJJAQTJe2msTy9Dru4m2lQeGgchbQ2eVx
C3wOgpxyBEEmr1TkfYdYdyJtxWpj2mM/7CcB9EiOSXSnyMP0721AgHhK793civ61J/WHmVwCsSLk
OqVhXneEkjv1ucpAvDZjsL6kQdvVze1HakH/benxWdH7vRFJbIFsGLIw1MGZszL+etrZ7K/9gyua
I8uj3KQFFoLFgQJ47lctmMLStdTSlZJFKFrDWvc6uxeUqRkq2kg/D2oci9zSHs0vr46B4IqgEqB1
2cCxRZx2WT1w97slOqnkRMmAOu46Ib0Y5yaXpwYaCkiVELssTU5fsJxU+ZERpFfX4HSAhPd7Jw/r
HinFyCoAFxdb6x2rPi8jEIUNPyotBaIXAngJi4IONE7Z6bnAqdN1wMVNUt+9CvMv2/5KZfycF546
xiGvGNIz26OnPWj8eOxDPgs4Wgrz+HSUM8yMeJRc3Y+khrqVG4mILGOKPmJAKQhF5CevfONP+OdZ
n8hYPmwO8NyZL4vbmvS0IGRrPJP9rXWGYgCQVjwzkRZTiIQf8pbKmLHFQWK2RW8ng/w11uAl7/GR
sVyWwFc6FQ/ngdgCrJTcr3Bu6Bs06TbkHH8h8cuYyjnqDAwabDHc093hJ6Gh/ssQ1Qr7mqt4CjvA
m1n63YFxpKoxid1SIAM8NVasWyz43JZgv1P1IHYD4SyS25vEFVgOEu+hBoQtjIjIZBpDc+BL6hmz
dHcJax+xfbzQ/XmB+VIAf3pOpw+4N19UZawtETX5/6sUEoTCKpYabYMTYbcpQlnuNqzb9BFJbx7E
jTNkBH9LArR6FrjIxGmETz8eeBuBX4dH1ZIhDU7s5ba5nyav7Al3HocHxPc6QiaG02WNky4xkjwN
nt39z2Mox7RU/CSJbH63ebaoQtdHh5oRmRhaeAmoF6QrqSASpeds/drgr6QIZhI4uQHauVXdry/8
+6nEGAWWNo21iBh7Hd9gRbnQqYI/veEWwEpNH/xJ3ZfS4lL4f7wkPdfbBG9n7yad3f33+RoGOJ48
YAVB7aHBgidKUsRAoCatgd3+scvL0Z7oBmets/ix56IdRjYsfD24sD595MuLhLxCyW+rekbCf/L8
c6QRUR3bsDkhm8X9ygaPImWxWAc464m9W2FKKnTaRHMdftNrVHnm7O0xNhEuttI3lG8zmPAU+JGK
pGrLspzksTbJfO7Zw0HnB1Gd0kQqCqqZN9aMM8gvxTBKDlHj08vQHyXIg5QL6vwB5idcIDKg5aBc
9VpK0A9I+JisjtHXvUgioE4rl3yC5gfxZXl+M6rG+ea45Bp/ldo4e933KA5vvZtzhx6f2aQ0eY+F
++IlKKFhCCmIWr8YFeetxNB695nruCzW17/9FggvqZ5TCR9hvPMYiwViSKm62PefFtMaKsdmxmq+
J49guyDQP1tkHBwIyw4rt4fUelUmK3LySU3TGV2UIhcFIJ35eUAqDePNYoFftRQvlLAcFjNfoP6k
s/9N/Kr9HBi24ypPAYF9SRlzXef3s9wjmR5MZb5cRGL3BnNrbcP+h70rwV6cudnMjwyy5X9sjYDP
PDPyVkvv/iuIK+uYBjPlrHVqW/HCZtJWu67W38eHXqSnUSmfR1Qbuoctonn7JKEjyRQ1tBaE9bNN
5C3CUZPdmmnI0bkLu8NYebM5hZv6biI9AmRmSgwHCIQZdMXu3JXbPQXBZ7qqJJ3r4uRHr5s2hbBS
2K9pfeH5ma1UcqRZzTAZF7khNEVYCvpCLJXU/Fv6UySo+r4CaHyuQNnPd7/5NRqYCfTyCjKVAXyT
KeKfIeuGGyNCgwHzSErE0w419+MdVZMhIT+SYQOSkid0ZYy2rXpF/YVQ6ux3zgAzlRB5vGrJIA25
NynVf79RqG2ppWUN5XeMg9x1HYX6jUdy0EUguaMQq43I4P9i341Wuf5Qb6OGYCFUAeCErRmc6dy2
jS7TQL6D4GUB3cf9SbPS4/+x5pdylfo8bad+oJvG4+PrTMsMFNBY5ki8NeFwhN/e3D0Dqc3WFoOt
coT0Ljcb8XkSDJwCrzDX6ozYyb5DrqvNV54/yJ1uw7EgYeg8jNP+zrAYs0kYWoeum+ULmR7Z7m+q
iDgeRDDNXsGhN6WAAGBoD6zu6AIuNiZwmAIy8zTsQXwutAqkrLW3aP4+LnSyS7D1Hwdma+rcHuir
IrvFN8/4nuTaISODvT8F3tS0PNll20VCajasHgwuGwAOduwq9xCjUao910iSmYUEMckDmkY2r3be
icreVy30/zjzQ4GtyGpGXisNyvA35w5fPkT0yhi7kKAvze4FQRN+MDkUYPfXxxAexEb/H6qA8xpp
N1H6br9oS8C/FW2hlh2IIMuKzG4rgMd7TeBPVX4LfXOLjjIzyxeZUYwwtIog65+pR656AAGG/JUA
x/D1ZJuOKkg6Jf/PvAI3HS095xQNwzMXNCRe9kUD9sUi7v8JhMEMmCyuxrmIKdpBs+wdZ3kBbQKr
pCpyXRF46kZdK+kZmiNOmTXUj4tRJZDJ88NgM3nRAbTk4qrIFcwUJee9wD+8J6n4RpQ+WPB8TB7K
HFJ+J4kjBxsojaGFFc+dxX6+c3RyvuIA5M707fHEZebXi4Bu6qO5TFxGzzg42p0a+QBfc8IH6Yz9
uI/EPxC6cL3F3cm6GjvsnxtiUXxE7jUc9mbZxbyp1yjv45ajiK6VQDqp0LnbRIDlHzv+uHjcTv+t
zf4YhMQL4Tkvs6eAQR/R+788aS9ONhyg2oFqrILJ6LztfVcbfwUA4WXzRh2EwQdJ1TvvhA1CH09H
h9wuvWoyFG0Ua1r3e5oMZoMu9cvsV1DsAJdhT+YJ1A9PBlALVINrlkWe9X6VZN5ha1IbXvqK0cXX
OU3v7BL0vXL70XB9ZkwrsxyQCBNUF4xomeq7Neaf/3ig19EmbGYWza8lDkVT0y19hJQnlz4qPwv0
1uqQ3rt+bwEkyYoentEUDe607OBxEUrZvgcqjv2YX1L0R2R7YNQmOdLIJYZUKjtyxRxSuKPS1F40
d8SBXLXwFeuHT+lqcHY/8Jzx/DbRneb/BA8i6B/xG/iTnUD82vab4LR5EKMYp1/YCn5izGwBK/nd
EMMXqtjWSCNE0huW6Wx9hF7AmwIVjsiPZLHLitLdsao7nHZFEzOMguOa5pH6n4imDGzGYbw6y3g9
yIpZXeH+E7Sg80RcRLv6oP+EE1W28TMptZSwIHyH3WdE9JAorsUogPEVq5VmsUzVMZgZl+AdHqqk
sRdzN1dCAx3n18kbXtxegcn1Jv99y03NSFu9aYHUp3+eIiwph7d0VkeYpyZ+ajWrgCqer168eyU0
7MSjPWaslFp1RUPtEdtf5S79zOTPl+0L2GpPOQr3SA6N4xmAKlc0fjrqlSzwk4KgR8pYAnWdiV9d
RATPpcTCuHw/rgDFn1aHKPl5RMAwRF9nK6j8hkROc1Dw1M40/c8ahdFcC+d/+agwxH1opcc8u45F
SE0XHHXmsLZ6wEbfYBuWD2lLbbYNEwrI0YMUsh4ZYFoOa3piV7kpDTFR3QSJGk+SnQ8m6KsvPFkT
nuLzMZXizhP8+ITpcrskFS89+M7JRoGRHX3QHzk1tlQltMqDUk9YQDOLXP2EQiQfXip+71t23+TG
cv9uDXUWTVPByqZh0d0dLNSatosyX4OzVsLpVPZk95c1Mipo5VVQ3eQfhGNTkNVaDEjhTJQ9vqfx
CBmFhtDWC4QeQYpx4WkjOYC8z5nEA0/VAgcGBf9XAx0ZTOEv8ub9tK3u2INH1xej+WFTXMVASflz
vVa8vWPBHgyljWExq3qMw2Sc5qdAMo/gDa4aKLTm4U2/XNKO2MNzVBPM1e3gbW5eb1Ndx4IDg3rm
UFv/fDYgvMryMRTPAwMM956CII4wEqNqMKICZfFYr85B22G69yES0mkC/x0mIu08O8+YhEgyxhzx
RTDGnZoFDYfqRbPsPwOBY0qnxu+arKt9vVeItPZrIBxp4m43g5B6xRyyDZLuaG8CxVRVHT8g7rtj
qk09Ha/K8Z/y3VE+SSOgS0pQ1sruBLTy//Ep+YvvVasPCF03owGqtnRddDOg9WMS8G/KK++qFrpk
XUVBDZCKv2m5WFkoxPLu+2LqyK930WLlcM9dNxkxNMX0nf66zCYi+7EzAx5Xl6N3O7jdaQOgkEqJ
d5OH8Bo1BPF3pQd5nWBFzrpyUJ7aqAOq6PU45LCtVaqoC8zNCXTY75m1CYnSIqd1VBOw12Z9hi4P
G1OTN7Ytcc9urye35Gk7U2wjUjeTldKEHonb+XG+nyHRyhrhqKqdAerjKDi13StZWGA2J0bBBi/q
EV/H8TaLrl0syotC8ZfrpPmuSJ1R9/I5t5oGl0OA8tGMS6NstvCz6/YGZ7iQPPewHitnTRmZJcmC
UwhdCaYBXDOuEK0gwIARoE+Cy7TqyzPj1k/SYGcMqv3eYmAeYsDKtK7v4KEFNMzUnkO6jUosjRxO
jB98kTFteOgdLDuafFKB9qOlwFnFPu5Nqb0GV7y1Awae8Ve8u3iXJbSFPbkvdYwTaO/h+eNngRer
fM5fe2zSTlQxI8x0bdHqMqkebCgBuu6kZQT/7SPzfRDbUWZfuyOq/vfAlDBer4fLYRlWmx2sV+8w
WkOqG8O9lJ9UjNOH/MmA2nYOPC/T7cRQwHcnLJs4MAvywSr7yuQ/TNIrhEjFLmp+4rY3jc5h/kqt
DAPgLZgOmuwe2evt1ryuVr0uEyZfbAoSpN+N1NTqyc3pizs+Un0m+ZfDkc+eBJHOcrb45xBENAGk
isQ48yPPWAVPi71hVbBKUApP4vMgCN25SrCsNhNk0ALTUWhTsnihDzXopoDogX2o0C+igdKBod8i
CTaaAcOXr2wsaldduJJ81Lz53SklneII2jvPmWBhrmnJG42wOIITAvKhrFyY9N9j2lRWm/TswQgl
0d0fqby2YJVjTiNPb3s53ncEo01LrnHzi7VjO+r5s+y+PK49xknQhcCr53X+uu8jDDCq+XXoqcsn
JOJn/hTX+4AjGgikMnstQMQMjQ5hXnXiaTINUHdHRZKDjZje7SmMw4a8IjSF/HaF4bYT6hFvK7EO
69GiZWPX+CXkaCPWwsxTd8V+rno//LbJ6/XVkvCtdfvhUfEm0TxYkJ04CP7RVCBS/qp7j29ndtVe
NJRBH9/FKFVjiQdj6W2TsdTpu641sUxSL8zMj23ij2MO1+2J5orHc3gdE57LDhgRHkJHfxIvAvN4
X+jNf6ma14Klbor35EDeuzbcDMb+uoFdMAeSCcMIuYLtIOs8aC/6eGWhekGTcbrnKGQWxXgShjID
0rzxx20KQpN3eV2Sej0QCDdSgy7gs57cqH4KuoeFzL+mHcA4Uv2IWQzPfTGlY1F9jlZ3NgRgCH/I
GG5hIWeZwyUJ74MwSTBEsuk3S6yv6D5Sl8WkPK0x8ht85oJLtrX3c3w2LRYFTs8SLy3NS9bR29pw
3JPJ/mBxGX8PoJkUvIpKkDv9zP3B4uwhd5GvRu8PMn1aQ1p25eFiyAvxXWMWXP7E24nTjE3qp9rZ
r8afWiDYjnwOjzHC3R90PF6s5OahE/pygDu3MpRp9KMI/5HrxCoWy71j01fsRRbWn1buwai67ECr
zO/1FvGDjgUShsJouJ2Huq7iaDVMqrQDKG+EgZBiryb/Ml1aK/XHO9BQ4mMiDDT4QNqCz2On/9uM
3v9Qi4aIVWdAQlW7QaghWmAZou1LPwZ3duA7EGvh9+CXIUdPr7dJ14zHCah+dyQ7buSkzcxiFfQM
XmKiF6zK0D8UmtkIk9LGaB6FGd2F9yKIkXp2BTiSoBijdDcaHfPw6Tvp6gyEIhwOXZTDoaTNt4Ts
CmHB7U1vIwL6I53oi35j0T838BRHWR28IjqTqeqqEopexE67VurtJar5XSbouxl45JLfKmeG/d7u
7P1Wv6KjR77LvyJePLn/m5ncrvqCTQM2+tdHZf+w1ATZ0VNXbIrOSKK02e5yQuanAswwvfpApjhl
dYscD55uN2RpegkPBCN9/3OypML2aJUh/IQr2MprWke5LHeqIPDbJ7HCmBrQ5H53yZ82Vpkcbgzk
TWyJ+MBb6eNk1NvWtKw4wm9G5fHFAVoPhR1qNH6DiCRP1O8GzVBJ5j8cBvaVsiN6JdH7RAd+hOtm
dXgK4n82tYF7RJYh/M4Ywc9nlrIMZvjgUP+NHCkQhiWXxEVpEcSG+kPMkaAGRfKAAaKHXSGVdQeh
Q6GN7rCUm23kL2DZ/q73L0WNEdVH5RRqi5i3djrCF3DpqtLrwbsDsWkrg3lIrZhLIRXpWP8ghQNE
Xd/c3e4IF7KnpAxAou8V+ksts7F6e3z+PtY2wd/GsvUwK6ZcuCiHXBOZtNudDwbXWG3qB9GtUI9F
ctV5srNWy4KuL41QZtq0cY74n38yK0C2fHoOVqPWNxmBeuytaHF1GFZ2RMcMnU99XIl9TVAi2fgL
Dw4atq5g+3ZvXZ/wip9vDR3rpujjLwY54ZiYbbu8ASTEj44I/1VFv06/8wETpIZXKitOPfCgbsBF
lnjXJJCJ4hYbGcgxi4j0YWb6NmujXPT+Qxp4W3Q0EU2I/kwKHoNQPrrla8kPnruwI2jhQVfbNaao
RTOS2cZp/cls7dVJsSxzSFzuXM1CzpGX14+jaC2uHTZz/xSvi4tHQAYtW1JVkYIJlIkjn62tCeAF
OYY5HGZae5c/9FCJMpKBLC42i645GHwbAKTPhpjww/npmKRTf2ps5U3d1tvJKqbI49beZj26tVcy
xr5y9KdxypEQTImsp15SC6kUfIGqVz0h+iRPBLvddRhQEboI03SVP3iEs5Ylht7pwJV1+ntGqvO5
+dWOcdlAvI1uqDh66wF+Y6OgRiusukr9upnLObb2MaqQYJ8Ja8+nDEadj+W6/5SjW5aPMqafB6hl
Hthj20GDkEtBrYTGN58V8sKR43Yvl6x3t2UWT0bYolbQ9g7rwQ9Rmzif2Lr8HO8xZ1+Q2QMZLjfa
FlrZrEI2QUjIGD/46bJExswKt98gSjLoIv1u0OVMbcSQ/x6/tXJQmdsqOh6NGN1AkGIbWc1UgEG5
i4H23j9sZ5DoXzkQj17obkXPpD4LZxhqmOVlHzncl0e0Py+1TsMyFLwUXSHIOHRR9TM5ftERfv0D
trobygNfYh7wuEDHGY6ohiEKAp886qtwQ/GF3PZysV+hCt2aQWf7Y17d0y6fOO+GwkPrFrBfPGn8
a7K/rAShZ4nXHoft7XaC9EXDBawp77WRVvDpw/lOuMLSf2DuMbd/kvbxJLN+5opWMQ3oCAxtqyUY
AebqtrjonkrOLVJiUPWkXYpMV8+vltMBGAWpd4YBcv2ibn6HBvOi7w59LaEghj4g+cVAzOwpDlDw
ph85Y4gbbGCj4VqbYlMgfY8lb7ofeCYYqEjMCBZhcDfjFU88YD87s0ltB46jlnqutvIfTGIezkj6
RlL9dCpv0dZJSvRHd5lD/ldZ/k2WWq/vvpMhawAY7Lbq6u3SpAsjhzfJqrmP9HhpcPvYfJoF61BC
K9OaV+LSRTTibtOAswy+Ka8fPvAGjK6FR3EC+h9nuaLtUNu3PagI/gmTXaFh7VeliiYkq7jUi2DC
nt5Gh84n/jMqEhiNpXtzSsgd52Pfgis0HWL3TVMCTD6iqoQWj0PbUWPGUNi2qAlnB1gjGZYEMMVs
mm15mv+wHy9xGAhCR3ciKpm0BHXXFjvyT1KtODbgW1Hb/3pxtvOkWIjRtcAmiurcRwrd3ZMQmyTy
ZAkq8OfjxR53Do+f/bqRYnv3mslv6tkj3kVMKFah6UZI44W4asLN5AmB42+D906ZX2wOi7OGTrf/
HzjAdjIstTleW0duiHUewq6fMuAkU4vyYJENM74iajX7yt9KYApyKEnC4nbM8oZ7W2B/Q6F/QUMH
ZYD5wDiSLyBE6/9UgPsII/NsfW61+bTYynCDiNF+6JM0jWU+xk32uXcI22YaviPPvFyZcJAu8tuc
DFqFtNWkCHTpDLbwtr5Kw+f0zt7EjFt9uRdqo2vsMpciyMFCPLi8JdehnJBz9zwsQzgKVbIQSp1v
RmkR7r//QPB/vy5N9RN+FNE621ITVNcQ0L6ijeKtCy3hX6GDTfaJZRd4f2dny8KOkHlDgOh1/tMb
ccqmEFHLOxAL/fFG2CPZvnrG+8OqHbQ4VqlF44TinfDSWef1x6ZWxDCzDztWCLUNTKMH0W1Ib6Iq
TtIAfPiCnnkOGthF8yahScF2/xx9XO3ZsqIc+iq7MSpAKwc0QUqfaIFi3mdcEsG026/0MYbu78T5
Q3TMwXOCcxoVT5mlcuHZYNFCPVAVhlUjjGIOI8R4aZRYE4xkf9sUbYtLmGnYSJmFyd1DrpRZNral
ekHwMzQ5gCD6tfOr1BCQYI3jWoaawEQtuLpQl/Gjfn4dMjunNu0SzWfZfOg0pJoI8K028qb2B9Ju
Q+whQ/Fhfv6O0gu1DVk2k9yCPCetSkOAq/lPIni/tLXvGx0rXyQ5TDgp9Pbmgt/gjfynuECb/e//
dXgoXYHmJGYfhp5vxwaEMyoe/0ha0OsbwCjp2EtnKhOTUXI4IsvpbCtb1lZtsuAmGrYQ8hniKorx
FthgGIy2brWHJrbE30u/OhnISBMawfgf59xf7u5DzGgJU2YC9SjzGASpOVkfrnYDQ18QuzeOYOnP
R+215jhKQDfUhLTeLhqdmnU1+igMNjzb9F1gG2rGwoqK8GLJzmbba1cjFDL+j3RG8jalRNxGHJ/6
wz0NZUX0zqsIJBKdbWYktKGErWdPzk3qGl8lcpevGJIJIuLcK/BkxBNJwOVGNXwdy+o6s+Zx1iS3
/jpF2Bpux3QfrZfL1SGIXYHSAGQRP/ivrNVqHk8LXevaxzqTsSosgnmc95afmNy9gRuWlmn+rbM7
WgsGlTxeYdXbnW+EUbuPpvG5CWnD1UL6c+elhZohD6yHEXzKU5LVhkww0LTVVsiEgOGR3bRTeLFw
/hcDX1Uv5/CBIn1JmOcjvqVcYtTChcxUoSsA8thc2c1YDIl2clM0s/UGP0AsJE7EoX3QrMUv1NgU
PfHCltAqiLrJ5+a2FmbI8KHocNPEQq5EUqDwTpbgqeCDtSDuHALv0cLJO701Cz5B8Eo1iv3n9Ukv
rO37wM/61cukzBg0HS4xjKRp6Oz0PainM1F7VArVeYdTwOIrNCnqD7Z3WSsXAZvSUH6jEWxer0yO
lS8LtP71Kxsvb9+72ATtE1jWGuoCK2bHCZrUUxRvnokHb0WJvCQxyYsW518AjG3/0L5x8vCMfoYK
pRQPMzKp+/TsYhcU2JKhJh+BnZx0OiJoqEVPbxF4hfYl8sXWWXMrFlb4nEfZXxcf/F1pXF4kJxYJ
Nhj1sXtWPkQdtEdrfzfXzVUEKnccrRh0h8r0gtlKmp0ogp8OgOrdhu4vqEhfcQRLIvpUNRaOlUmC
CLVYC5NbS/WWHXAn4pMpdmBizE+Cm56nQ3fUjPjwZhfvhGGPMWwMom3wBX/7FEmo3jjq21nA/nut
fATaQW74FERGHawjee6sPe6aWI+E4KDl8Z+maa6a7nGbF5ToAMd/nk5ta5VWmOeGdW17bG8kBbWc
oYWw0Xw91n/Ilc6bJNykPhFWdbixh3Md4aZCTgwlPnmFojePB9ATDL5JXHAfyBWXDn31HpgvFJqW
gOz9Kp9R7xuyRw0m/H0dU+ucgaMXpDimZN0sR/U9NijnKCo7qK9urxOBQQtD0dYcT9ePTMYKKLy1
Tk+CapBbIaZ4Wgmhara+qqbPO/qjN7fl2ncvKITvGZJ2vSAAo+DoUXChnyExu8zrrYSZjjxCk01v
nCwSDfw1qx9RlfbwXanHX5w9qxzFYsJ+yHs4ZLXCmvk0dntb0+fGdYAsM4wNwN8YQMG2t0b+iAzP
FmLfjAPNHVjp/RViM6SscGX8b+Ac82EZi5hQoNceDW+MLO4tWfQTyiCmtmg4WzLNo/1JOn0IGGcF
dOtBxVdQ5bjS6w7kHPAeqf2Bd9Csw2wHM+7zTANPRJfzxT8x3CdEtrrqY2IhMnZD5JIDmiXukbDQ
EwVmv3mxkiYIVyf632pgiNloSHRktZv03I3+FFDATChEyvHym/mkCELZlv+5jjv4dZUWo3y/c18s
M/18JEAfnXZZi5KYM31xGtRne6vz3ri1t7TK/Qvrxxc9XNIp57PEGwL96EqJ/PWoJ+PZsTnqc5iL
mRMKFkXE35kARx9i4K6DWeS84z41ie6SIgNX3AK8DXdFldjPYdJ6/h402N9vIGXG49GZfmR6l8tK
JcHR5bu7DJfBrz1QbKmLgkea3W1pS5e7OKcgNjMAa+nuURGTlldsWciB9GbnisQBiy6NG17VgXDz
ys0ck/ne4sQPDk5iBciALJQBH+Veamkj4myjuIGCIgjDXM4oV2wYO7b7QLvagCA+7gSFLUnfrwBC
X4Rz2MXOvWzQwIxSl2vJVPU5YsjvmG7ELzi5A4vnGUNd994EiCrnbgs8FX+jx2yhBqavOc/Aln+D
uqt/UHo+6Kla1JjebanFlY7eat9n91l9sdfqrFgU6wtoC7MvhlGmhlw1byqcIaJUPCn7PpeTh9DH
tprksRFSX1NfoZa2tirgfpzM5aV3kJy/7Z9ajn/uP6Mjeo1DyU5wg75dJ7EasP2pi+tf/J5XMzOe
h4PzaC89UWvwFUtXtSTK+9pDaXKsdpZHKw1On32bui2QB1YJD7nnbVCrczJq0kx0/AFeWdgKyDeg
DK8aLxVHC4hpqyFPOFGiZGK+UPwyUtnIh4H/FfUDC01OMANlVFk2lTNFmfQtu1cPEKaN4+QG8+lk
bcH2E06y1aE3KWTUC4x5vbHAbOuq+XG4gdNPSUYCKf8H8Dipvv12MA2XeQpmsRk3qDWBAaOqoqGu
PJrLFop/AD7N0EzXrBYbyMCnDsTBIafiY9OCfEqeyD/2OgIVsK89vBAZXPT4MzRG8ZL2Wi8BkSxG
sjFs2VCJzwY5NKaPppdjacYRwjaJF7IsspbLsTTecaFOWD2z2P36lTBaKxazwbWnqwkRVIFbznNP
MyJeQA3Rep9jiaAUSxt6I1audM5Q5Ecximk7FINJQoasbfPcUXeEZVuXqHQC5prbT8cASw1tcXL6
OhhdOxGeUvQrZBZhYk7UyzcHTZiLBNw08des3lzxzXdIUmmtwIMpP4Dxig/MqfmO/RLolC5UPbZ5
uBwyqXUhH455bfPMzKmX+uQPVBrhHU/zr1F/DSU7vHjgA1Kh51U3FfdxDiMHfo7ncZwN7yWF87w4
yS1opmKUJur5RlBM1rCnBHDGHltgXyWzK+desdB8SOvkPPKeUUjEsv8cQegfciYFXSKJGMReJgwC
c5FkfK/9Csd6wJX76qAvLete0FclG7u0FU+7jQNFwWwXaCmESQikQfEAOd/XAmhqVZO+x+2V7pBy
ju4p8MqDirhp396Gri+LPuRGHBdN7m2IW5DVB5kiYUfhEj8tg1drH7auDfIxnMoDKWiU+q7ksxBX
DXjlPPkiRZ7qs4YNZBynJEV9ycD910vuweRvQnGbtTDYKBKCKATniItR7lqFAJRHDUyTaoO8dQQ+
Bdv1ng/00/q/Ee8gsUyVVF4QlyAApdWDoxiiwHWyjGK54jHc/IVFW4UQTuiHCcdJwYzrBlN4IQUl
2JQSDIud1679UNqUbpRO/56kju5UD0hnJVBpZMVdurniT0W3/0OaoNdIgZt2BuukG767y3I7/aEJ
YBnZirK86Zu8dU0rUDlNR9G9TVHU94hfgx9xmUwh3C53aOggMQzLcjQ6Ich159IoJUKV0XSvhEbW
nrQMRNcvbDtjRxps0KnojgISjkCghTGAP29a+2n1Hxp3pnY9x9IJsNsT8EqnCHXzuGbbmew86Ttv
xv2TiK/92V69g75kK0MHAiH+d920ddfE5vEqvAxhqaf+gv1XuXQmtadpC5HwWreCUWvT4jrVnOgo
Yd5vgMp4AGGdbGdvEtNs2GS2rQn14ScIvCC9+6BpSq+t9HMsghvkQ8MopgS6nVl3i48pTCX1GIhQ
7EZKvJmN0GSvL3qwg8+e/mPs4/KpU3KOQr/7jKGgt1BJe08eT7ew0F9bFY+Z8uP1OFSanCaGiYra
E/wdJ8cdI8q3OWm3XEPm9o+ihA5K4EmfAmfgSbf7uqip67AUE9eUiMFhC6jxP0y2xzAGUw47jrDB
rGr6+ZHyyMhauqIPwcMF5N973bUsefBPuDhpzsQneM0ggVjv/6f4+v1RmLacFTuB1IaYt7xLLiBh
tHcdCK9FGqWfc5OCh+1rF0F9Xuxwf0OLJXkHkSOYmz2MrExSB3oY7W+PafeDLhZPSOTsVb+WoHLb
SQi+r7ac97tKy/musVOaJ1dZp238nfXPRgL9Ejs+dgfxhkTrCz6c+8BdieFaFh65NcbcpLbmOBm7
j0BgxJRcswwaJ0EgZt7aSIWeSEMTD+ti8A3mhFZnvJ+t3yPaE5psa/xNQlFp2AP+vhSWmhE0UQzV
3jab13nOKY1w91AFzmPoBaMNrK0kqZiFKZdgclW3wb0lGVOrVIJltlRMlemaKbDooa2/L8N+wd8W
6VGNCFda8QJBolt0yNIrLqgohTrZh4L2wVVgOwOoO+8G4N/tFNYUJFDjlYE4iHpS4fifE00qHsnx
6eMgq9CpcMZRy0+nJP8ZNdZiQ4F/RsiZcaxej6axxZNtc4CKFHJANDh1dvBaNANb8r5PvHoSGTer
4Wr7WqCl0lIYQTtR057Ag0UvYrWKssM7OYeSxTPzjMbxXNtzYIO5lP2AQZXWYx9k7VZDL5cS24Sh
uiNypFHdZD5WmzIR7SMlkWlFwDmhrMjnZMGrodjxWedmDbXvGbfLZ9SV057mebG15ST2hyfemOGe
DqK8AgVeMkmcf8TIxkMUku7+/woW1b5cdrkRmrkGa443zzzboTobSzoMO653Zd8IIdUWsP4YhnvL
wMeQcsb0QqTTE2sIqcthxP9s+ZJ9RnmXszAvOXtjGDJDQDR4MlxtJM7bzzEAA8xgUwrdGoLwW0uK
tGJc6VY0vV7P4C8rphlhqkrcU+VpyTodRcfPrAe2FyVTe3JWCsn5kmGS4oTj3/g+xY711nizcLQt
zXZmrW/uqvgRG646lfnahC2yKT+XEg1uDeO8qEOqwSMZU2PjbeIER0DbEhmvKAFnCwVPlk+I1rIL
sbLpoyJOhOzwyneclEMPrZxX9t4XYzT4aPxMKzj98AlTDgaWQJo1Kiyn8cvXk2NzRKZknvouD6O9
eDj/sAx9tIeo5QWu+g65hxWisgABdj5Hw1F7BB1rxr8U0T+yjGh36nRR/Yj3YL0oAqPCfi+uq1MB
dOTDA/Zs0MpG1JaKS6lbCZUk5QnorJOoWrMBV++XVVc8QrKf7Ugzg5J0c0cpGmiqYKC8SJYsa0AB
8YmNDTrQvxFgZ+s2n9bDoufy9S1DRmA2ZZMdZzRPXEMlXetSC0dMDzLtnwwV7DTevMxrFKuHxE9g
fgBthBuNoIyKLu8bKW3yVV0wJQGr+mBPd1cLfy5eJCPDZMwzjwVKKNi444BwDylyQtsVR6B8iTGq
e17kbg36GVKamCNdF+P7X6NhNSit4yEG3h+qPOrQk7omqU8F0T/RxrzTiPN3me0P2c98YnWucoHA
aqsFtD3eFfZx7pkObpWXxfP6zqBpdhX8yP/6B1cVdihRyTVlfwGrFTe+kjyPsRGg4uSDDf4MxbNO
2Bsn9jiUhjiD+rx4mEmCptda8oLyx03BDhvZKUdLUL6TgrO73ZERgCBYElb2NyLZr1gkhflD0+dd
zVHIZLsZbAb8Xkyt2/fRBltMxdyLB+shqxf/semOPut51SDSFGflFNAGiAQAL/k00YUY3L49x5Vp
/zlW2RdQr7sIwdZtG6cQiPLQLg9EOD58X2z58e/ULg4UgLucU2DyX3ggUSSzg3n/TV168JkbfVA6
TXa+cFlWpIBzuLFCgXEy3b4LQwwmmQb84ZKkroLwebSlwbPc8itsz2dn0/nuKWQlAYKxfcpQHlBU
vaPvVlQFN5SShjecut4RxLBG1q5l+Cv81UtR7Re8oApYJuTDxJ3FlXw5hrBCyV440yhp4LrBohaH
M62Xpx67r8v1QfbFdA51ExXeMMSg/wLdQGl+4n/WaIuv8tZZrIC0za9ZToy2WiJofzLF6zclncs2
BG3iqFEIOYSzN0W7heSRVkevQIZz7RlNJIsPg6nebWo1XOhBGYXaYbHPZh7oHgG6bq/vJ/2t39jc
WRpGtWe4c4SOKwoP6IgLEzgYb5KvTVZdfqjZKy1M/eLDmlRuZL+BCMe031GqOa9GzxptLuYjB1/C
zq/5+h95lKi7HMr1fPrW7Jj2n6geq4p8e4bQpbXoie4nmPaP6FpkVnDO2cmSmM+Wzok46efUcprd
VekbyxAJNVyQZRlNlSzddEU1lrGY/bHIYgyeaQkIZLGGVVdfE8YZnv1kEGYbn0q71BxykEM+MisM
uiAo+3qEsx/WUVcZ1cVd0NoipVpgICE1HOPco1xa1RbditGQ/72cjxx0gOhvrk3Ro+oX1HNlUxZq
xFOb1fs7h81S0izQaoA72kCU0opmW9vpYw9v84wlrICnvGxT4V53DKHsQDQsg/h+MNgaRDZHLFwh
UQ6v9JFhWwYku1sJHfeHe1+1ZCoEbD1ylLTIrzR7Puj0e1ziD7beawUDJ3aD6/7PnSSNt03d37PR
55a/fytZgMLB6m3aN8ZqytSEh8DTzTgugr2e1LRHXWKfE0HSZUSxsz/wif65iUTeJFnuQB00NAz8
C6mrnx7NLHeqbr0ET5ebXbVH5J3e8dbinGJAzKSdYwBwUOBUrgarv+MRo/mSRgvOlXVo6qkygrB2
ncpDmX7211+HUG5i/OZlRIKPacNoSEf71y1j4TMxmcNI0F22Loe6OR1GFtPq0n3YjjLPJPJeee3p
Ag5ynQEJtIEI1hdaUwd7JGGBMneMjyFGp4kU6U3j/eW/CPvq1TZbuIJaH2VIMgMgeGiPPMzPRXr6
mpfYCBh9PjFCVXyH7kCPdyJW7xF1OYyERSp6KQJFRDgdHHTQq3g6e7pGrGMhPo4+HE3WorKKb0nk
S1JvfVnNsxZEr/6VyEvfcbdEHyg9toLmPhAI3MhxxJmY9HyRxt2ZvZ+6KamKz0GrlQR/+hiwnaWw
zMfTBFpw27C5riuVD2gMHGN8MjevUeg1ew/rDIChVOirDZTCIeVsV1ayGIzTmxs/syZe/1z9btUF
VYuoQ+2ZifjsF8LDCapkZbM3U7DMMWwCXd+dUdymvJMBWZxTULuDjT20E9WLnIO9aflb4hakYFNF
vr4nau96DuKP5mAV1mwEFmVfyWtg1ZQ5zvTcZFMAKIftXDgCzXJembVSIssY/n87U8wZ+TqSwsHe
u871m+PygbJzdg3g4QhKkxU7TF6qdmBoRT18UybuH3tj3YfZKZNJpPnfZpz/6xEWJ6P5KwtXsJ+7
DsdcR5xNNmBf1RlkMuo8nSl2Q7GjKTfMM9VO/ZImOLJbp6Euc0iJAf+4N+vttzdGELzZDresWmFb
Hiw/9snx2YQHm0FjyFjRmwMOlt4B2EwUKEvkIOyi5oBZmWwUj5CFV+63cX3IFm2uz4wmdWaQEz3H
qF7HYT8U8f/syVWPAZmkphkALKj+hN5XbsNbGRB6U5/pLrCWAxQ5/KpO129zTTbp1+FGGBHu+OZv
0o8IRNFmVMSyPjMYSnEcz6R0IScZAxzbYWGF1mV3KmwsznUCa9+TQjwsEJtMGujVnPRxbY5Eyunx
Mcwqw3Aabo69HNj37OpiaWtFkOjejfrKNHltbk7pipqdI6ln93vp+V5F5rYYaxEi41BvAsQZVPE2
1E2/32jSOlL+4H1tf9rdlU/fbUmD7flgzlfpKih+hsznMSF1hV+117rdHZ+jz44HusTYs6omIOIR
nFOeGzWsWHug5cObEoVW1L7t5d8FRXIV7UkMgcIgD/JkRnA0W39m4NFnJCcU14Y7j1iItRpjvgvq
4jdwXDVxfYj4FD/jSShCvU0aVlb+TjW90/w6795ai1qL+mVKpqr2lOKgXLWGBTURdGhBZ3NjUI6s
MJ521KsUhqYJBevP/lD/dDBABRDkmWt7uAUJ10I2xEElmx/mRjdaqcJ44haIsCl0nIfeqypzmAEA
zYGNCpsqa6FKQ1bVn00iJuXXDt8lcSAefVxUoVV5AZYRleiRDPQZigeASQ1tR4f7NoC8y95p4FKB
nMqEcXr2KsPvaTNNM9fbCA2Xee3cyiYynus7YupernY4a3+mAKruBLqAuHuaJMeURdfkR28ZZ+rV
oQuGKZfgYbCJclG5exyetYLPWzOs5hDfOrgbrTSMSmar0ov1vnW0yfH04oSSKXjJlC1JY+U0XBmu
2ArZ595vilywtBQic0klOQzKNNq7XHXnZsaWEy40D2PePSs3S+wIQULsrEMkugCp2wtu5sDY7HAN
WeBiO7Fe7xnMdtUlO6Vlcb1dEQfh4PqHJ4SSGNKaeZVtTXVWez8L835ub9IRqEEJnE85gtH3RDgA
5A2DxpQuWMgw+iR3uBMe3R/P91spwp7WO2ID4LlJwjtBvfXsIKbPzXS7r4n2Mnf/a5+uGdZlQRJQ
qW82tjlU/x90nIq/S6t8Xmjqunq0U8xUprUlXq4leWQt1hYTC9dBSXoUSs5J4y9DMVDwT5oC1c33
bAGXSr4MVyvGmqG75DyZEy161X948xX8beXBW5dTofGBJOzaMbsv7jOt9u8OGX7nx3tXkWwj5fRR
L7TkEPYHfy/xTGcL6EH6sO2hOhX/zbjuYkGLWo0+0ejQnSMF3O1mE3ftXw+dwsUQfQ0GARkGPB01
o7VwGFxjXdW74dBL8Pflu4BIF7YQSXK6FIvVY1ss51nhV1271gR/SAFkhJxiH8YuEzLcZxavkEcp
voHrNhAFpf6wlv/84qxAYrRh5UnoVOZ9Fx6FSgVaRjgoooRpoHl45pIme/kkoxMLWmQaBE7HLyqo
rHEkFECHNAyoFuGF5ZIL0e1F0KIXXQQDv9c2U/WElaOgXBKf8QSf450djVboDqAfHs9i7K4RGUYD
PDwEK24PM+AOEIyE+C5vsdbzsag2dpIt2Lo+TX8nS7+qqMJvR9XVf4/IyFEwRmzMSgVVCf/1p64W
gcoUHPvLM8m2fAVKow/hNuZebrKv9ogaGAC2JUdu9P9wDYKvpN3amXN71AQ3FS5ZaS/eR5eM7WPF
RMolbRQm9FPRxJTkZyfVYmHpSKz9a0CXw0ifbgZcDDdD9o1SxXDoMRzA4KQ7flh5d+7yjbFVzSg/
EwSvt5SavwN2WItPlHpuP8PklSzvHRI6CL0MmD+JV0vt6FYMqSCsvYT70++Y/ib+rLiWucvy5mXe
0RkCeX46AOmpwxOCfFeKrENqycIGRuhoK8eN0jlT2e9bp6RoahrmFvHWMDIBcNPtyZbnqD8BgEyS
y1kjIM5yd0KDoP+2PnDKiGmx7wXmWHyFiylmjJW+KkeFmxgAJUGVHNdDUs+XCR4RtlNzJ3IIrEqN
7QYclL5ApR4qY7001RBTc5Eiq7tFsuldJWGE4x6cJuwnw3y2FZRMbgrXeRX6K9TKE43+PQVKwpEm
MAmNr8FYlEFkk6xU9dk+PsicNFWXlZ2C332/uOez73lQKmMXOZvZh5m6Zy+KJj+DK+2QwDA8JZUh
dBEUWllTs/U+yXFssVdyFY+gsAan9ZrIwxSaSvfTMaYERQTPKuKIn2sFuy1qqi+4mS50BgXEdc2z
Z7H5+qNTLY6dSK17TYmkPcLfKAsCnbRr542gD/pGSMhkkwgPFSBpXuKqMVoK20Kqp7/4vkWzieGL
Gf8br/WiEhnbeh7gNEr4K0N7PyksbyFKB3TNfMq8HltHbmlN7IbR8APc7hs5gtOQmESz4GxSj5Xp
P0qjpCyiFrsly6x+5b83SOqqM79JRqeau9MYyBOYlA3np7Csob8fWc8szKU9DpBkl7sKHAbxwicW
nURtAOL/7suVyU1PX5xe62xqObnfPw/N/IE+rvGNzDBJ/BgfjfGiH4Av+FphKHTBxg+U+Y+ycKRf
H5RxZUsgizAx103novJnZpRbZscHPWJNKZvdMiAPX5eh9X3dy9Z29Zh71lfpkdhre6/2zFRrHtVK
+zWSnQl7WVxg378q1acuWawTHygg+Dg/+UYfK9bvpP2U+1kkR2s/APIjyOrRYeqhCplvkI5pm0lC
6wGrZ19hjtr+8bUkqRAailSArewfUOmUEWTJw3EQeNQHsCgRnTXmW9crYQ9T9oh1V6ukE5/mKp+M
CPJzGHdh6Iw3Btwkb/fpiykbnlBTHW3/iah1Ox/oUIxbXZ6ygiqON+eOcrbQ9Fo5tMUDWRYhjgCA
FV48J3fL3pNT/Ze/bsp+DSmIHx0hSkBsKfaD72Q1LiCIFVjMJoeFdgTlkeioHbKN0dQHMASNDktc
P1Zozx/COj39INe4ntnYAkstmS75PLwsMdJkoz/M9gJSP4y2zJvfSKlt5yVyvbl1ICVY1Y/nM0Ue
Wz3rvzCM0VwRcp1Sh0mXixHVGqm6PqIuXOed1+zDeEjxCYTcqjhnYd5cfx5y48ACOM6TjgyIgwbJ
ktYWf6JH2uJ7k6ajF01qtbYodF9/xRWHk7udpG8VfyBNbOfpypMteTSDCkdd6ddfjjKlBIjC4Iaz
ywfNUPmUKyRpFuEUtlAID1XzLeCuehM2jM5Ai4oEryxYzVVNbw7A0x5jBS3i8E2TpNG1LQWGttfC
KGd6NVtTFkAK5u/nhSgbQDvn0vR15cFYUc8KTugIVF3lvVyxkuRnCRwvUTU/3GBLX4Fh14MzYY2E
XijiAgRbaRifAOX4QUY1CqwSgVnPawSJs/v++yeD9R7TzzZ002r9xhY2MI2Ur/47kaYlDtB6XtKu
g8ssDCYkWahfaUqP3dlJFyGj/C8FzcVJ6J7NfvqqkmWV/fys/mC6Eu7+yVkxHqsfIixJHYj2VXTV
y1u2Lk8uXBBZTbi3cAWMwbK8g8F81RZjI7kf3u2qrgylx/oGOXdBRlyNqSPL0Za4yvAT/8WsHtYb
AOwsWa5eT0lgioUIz9iv3frJK0bVbeF8XH9VvPeKiTRf0SgIl+uy0J3xmk2BVjorl0nqx+q6rw8d
U490uwRUj5mdzncaa3iTC2S7HDcUwKRHEc9j0Q2zyKqfubC/MddQ6UD8E6TkhDWnv3tKPbDyGrTW
HJ+R/J38O0YMljAYnlaa6fyg+qSjzKkWJVBxuoNcnbTzRhI1SZBF0mzoz6paMFZ3tabj6Arut4uA
wOxGkrphEIKk5ajCBUAEgOJeBdGX3efXTuL3rqabI5XiuxzafybqKFb4kyXwzk7QNu32u0LtQ1Nf
FCTYtiFWHkroNJe3iOVDqsdFdDxkcovo5zZHq5q4iZytnZA6T57vkpayMpSVrkMbs2Q/DZ9AxZmc
cz9DMaUM2LW7TBEuA48HAwaztaqpQq1c8JsDnD0NHD6gKFPdboGa1IIHM5NC0GFydfjn7O2Fgxfo
CrUadIIS2mxt2GZ/3b5JXI/VMsFhye6VRCxLhzn4rrH7PKBTeNyXLNORqzq45JC/SPIMJFcaNsFd
2g1v02071ugzjpUCUvkGd519ObsPyvASVl1M30caM+7Dr2lCsbmZclwTphA1HNmCdtlt/qR9EmMc
OdzL0Epxu5cEGk9Io7IS68TsAVgjgX6ZW68d+iag1y/2OpkBPRiv+gOTF2lty7s46GxwoQaUk0Ai
rXqoRVrQlFF+xmJKc0AnFGELPCHxIImeSQMe76NnnUnqDrNNQXvgs9IdpkUCSX5vpB3Y9PG//YyX
JPESFUu/9ON8AahiSfgXF3qZiEXQtz+jnei2c6kmcKCqD5h35X3VtWy3NPTwN7rRysrefjzZHege
HVELwjsEjN46Yqs0EBkeBVd532/0n6AMEBi0+3LX1mi0s4em+MBx2yi0iIztc8rLghieKN4fjNxI
DyytOfTfAh2OT9WB5bvYYRrW8K/zWKLrt5vyvexQhdGTcV4VcAE8i/HdbQB7yAAlivLjpg0GyIMX
MbTezdSyv50jFElE1g68v+uSfZ5n6eDdy1NSLKqNmkHYXDxfzkgbHAOBmcqjcT6lB77PsRFZD1+D
V2i6RHKwwM8Vhv7egHaYOhrlXF4oq4qczOI5n0g35cw+8IPNk691f1ZLA9mag7a6+mziqlnwhAEb
L7yQSKOzc2dfPl6eqMc/NXzPXB9DO0+qcepyU7Ad0AhdO22OGw8w+hDPbhpgJuxA3UbZ9CVfvyHW
Wf59Kic9djXJPtidp98Ml6nxcE1QHf0zqpn671Cqnvl+axqoAWUUZ0OeduGR/zBh9ms25zHaj+nz
AyBm+eeTNy/nckBIt/bvEXC8dU1RSGNx7yLded6P78B+M81bilhyri4u9YLcQAjBySl4tjykrM5U
Dr5r/WiW/WvKdE4tyqbZgXYQToCyN6g+p8cMPW5BuayuO3AhzQcxkMkRXTvxzVxj3ggv4Mg090qu
kchE7FPn8kpMjwrLyyNG9jplBvPhBvSKSfA7JugLqaLBBY54ambChyHq+nQtVEAz9YJmUTotVN17
y3jFVut55+agGPsY4B8Z63SQWOOn7zzdB1CPaDG5KNCKrHz5Zuv5LYLIunTFf+TE405kdmATrFPS
3pg/cEgV1bRWa3cyNiG+qetATQMcA7lCxZaQ2dP6IXo8So+ckQsBql+W8iVJBGb+EPH6GMo77hbd
M/BqUJt5BZN6Rd8lSn8bxhcUvOiMzrctF7d+EOYfsTAMJbhF0cuIH4OzqWQ90PFfFkIOK9eln8Cc
7pv1Kt+S7wmoNm6JCu+/WWOAm+nGj+ThCEbVhRNNiNYnr3jb2aFM1WgMt9CpWsIaa4P23J2J/6Kt
cW6ywpQWEBhnBLWqR03sG6Fu7g12DSA7eG5kGBu83K4LAKSaeDRp+utdFNSuaTfmPgbEfFPRa/Te
6IK7ZEf/GkD5mLATjmwYu9LmSw1f5754TU9kOL4X8w5OF7YklJHJaDYthqyPFGdiEQW4NRd7eNMD
VdteX1BTfBJRd49KRR/sf9D4Gx9R+8uoexk09Ao9rEGkfBQbhsaH8McDgMpfefY6gTB2OjcmIGa0
/G3l9EE6cGcdVkIh3PFZGj4igT9pCavSUKJTaHUL+MCzdbVsPSFaW2f6hVacrfsPoHEFy0J4D+KY
gVaKQIK4OGCflFVHn7p87l9GckC1+K/FYLBZMBLCpua/ivUUOL287mphsLsJ4W32rRVLj1rz9MbM
QM4QB4NcZ6KVde6P2J/Y5iwPWt5F/ySPWEuGM7wPYy1T1m/lT637BxXoNlNwPaLhPqhfFEWh53uu
14AuCqhdgdnzKYPIcrzzEGmaxeZe23hN+v9tth/jlfrxdWSaLY30zynWg2Or12LwwyBUpT0FUSXi
xYKetHrnVQWobul55Y1EWyZax25uHEen2U9bJZsKbfzXV+TfrWeCXPWU8NsrRLPZYb7e4+roe9Sc
G70CdxmGuwlteWgan6V1Jh7y0pc0EkMxz5+MlRMxXG57NTaqMxJMJz4hKzI9DOV6oVvm2su6aMoe
6jzo6Rasadb8c0gqpzkIskY2zcys1fQwRjzWA5dzywmB+cesTTD5d6xy26cr+GGVDbnH2y8Y/K0o
rml0b8zoorqNRAG+kxxHiAxMEhm4wW0aGaE3tvvi/U/moBrgosccAn8Pu8XrfEtWrSJB5GSBal/v
123E+D1Dyo7lAAu5b0pOigsdS4U1E6TGgdmd/3ynJB1s7XwwIPEZ5//e1XuyKhWyTMb71G/jloi0
2uFcKEPl38w7gMD43B8mU8rYVsAnfwRnq4h2km6yvglv4yreLCVbpk8Yl4WHkRRuWgAD5/MwsqnF
PuF+MKPBBJc5Hc4CADRVobzvNhoJUIY8QORC+wViV0fPoVSgsVxzO34hCbw1tqiiLQlw2l6JDpah
MjFNNo1qjOsmpUMXkDUnhOgcBfGmv6KmTXGVavV/edyj7QE15JJ8DsB831dOPcWm6nuEi3t8GOFh
2KgCnc/eC+s5oVgU6To+7cbjwHdRXGyF+wbwFPZk61qIo9w/V+9pnuQz3WQVNklQcV+LKgWSm5el
QA3+wXEDeNjqIpPmHRxJGkINU6Dob7r5GymLVw2JxwSUc8yhTC6Xh8VR3viH/FedvEtH4CCuUGkG
zv7m28Z5IjDzevLRxN/POgCoVscef/QHXYc96107cmE9R4yLmyZISQ6hqTj+oLlVTIURR9ZQyH3Q
DHolIEj2gSJcWum48IgDkniC76ojO8pgajbhsFnqqpC7swyJf9fBjJQ7HRGzYLv4tfb3SUgCImud
dJ5OqcLnW3SknC70Uv9dGsi0JodJLdswMXGCHANgKid7qi3mMQM17hCFLo/Pb33fkJpXWuZ6zkFx
GdRnE1R/7olWmY8R8LrVXS0xE2FKWLitMnGk2Ul6od+ikneHrM0ZC0ENQzULpsqzrXifwitzBvt4
LgmCTuoFASXEJkG4tJlBLzowRkwXP/0d4+BCTwL63AIZq+k/qxfYjeS4quD0szDDKXFXbNuG6iMW
f0cF97uIUSpAso3dMIklRYtu5lcwbhs4D9V+BJqpF0qiPUl3KRpUyHfw7QgguH83bbLCYOuxbpXV
vUEgZsil4OS13CZVtkud4nPN3DT+AX/Pk/lVOoVVOTe/Wd2aB9P/I9HHP5GWtWOTkPgV7+TdyACV
OIpKeBQXyVG76XCxEXxcnVvf6+LhRllkwdOE25XMon407QPpeDolc/SQnnc0mJhgw9OeCbVOaSUB
GrkZzK836Stea0fNVpCd+5fq9mzFDBTmL9ArRGEC1Ox62y/2DRX0rhEvWLWkc5OdbNi72XwwXcA6
RhtLkWi7+tIdN/QbD0T09YAc/IvnfFC6kym7GYv7Y8P5TMiuMp1rnRCf+xCYtnFDQxc2pQXFvhtJ
VcKvJkDcsQejSOesXIZMWYO/7hcvqsC7eK60aU4AVWvAxfVrXa3tWg7LIYp88GAQPG0glU8KTXaU
KV+DkWCQ0ogg085qBaWa0AIQowLzxpiBq39e1PQbnochGu+X6jJcI36y1op/gba0HvoDsCEmmlb8
NoqicP1GfkMjykS4hHIyf+uY6fS7B7ACGwMf77jsugv8gzf4zUbu8ouFlUcvark/bKFBc6ds+Pg4
Y7yk5l6FcZqOI1XE0JI+dZuhe+ir8vsCWrvCjmwXwIfWHa2oyzgMCTsf6Nux3u1X/sheC/Jvn1Or
tRAVm0o54YHtWbQ4zXvXOZJlHoE5e4MzUCPnHwOXwne+hzLUWU8li9Qto6h+cdduL9UFdE4K0ztC
AUxU5rdb8CqIEX7FO/9sxEJ9MLOd97Fz6prp+qmdKVECIBOChAneNbfnp0dN0Gt3j221u0N+anOA
CLt4+3owDXYVGzCDUY5ITAXHW9kV+NvJaAB9jzGnPYnTRrQ8dGcBIbmnlhKyxzKl+q21hyojv85+
58dsWB0lP7zT/TMlGeNEn+91linFlJw6vixs16GXcdytd1v/EWMoKr9c4/eiy+Jn/BI4mo+3Sx6I
1gK9C70GVYXSwyeP8BySd6Cyt/jW9St1yJ52+oWyvBPXueyaKe9Ly+qLp4re0wWcj6tbE6VeThm0
RwJgI4STo8MKR9AJoEpvghHnbUFyA0oUXA7k3XZevh2E59VK7/ddbTml52Lyb9OuAQHFC4nWIi3g
Udg+ueC7eKv2/gluTfo0edlpUEk26TuwFXo8I48lfHS/PPHdD711u8iuZkOhl0pjf+xRMiMwGqYh
sM4cIeVKb2DggK6m9YjWnf677niIkY30SKJxMxAYD8fbmn2XnZs/4jIZKFm/fd5Vk6NA0aLqGWnT
Z6cTGlRkJCwKjFrOJ0HWO3HoPeKN9TiB3xbKx7GejeW9qhDew4QWqtwabYNWHKG3wbX4TwkNxufD
r6Y5u0Ke7BCj5JN+s0tBgfJLo/pvh1UC7bNaDyGXFszUbzch6eXr+DoeoFGUm6hIioBX2orBxASd
vOUDz79DnkrxSK9uE54Y3Ge5KRKcmBB/od8AsUswy/Ex4X4EHVFnltM/yQfewjM6iQurpwsfMgkc
N7R405q+JIX4GrXhO+nzhg8qtWeWsiZFvskw5iyc+Gj0VCkxoPQml0f8hOFraAvIqXWg78+m9xBe
Wvl3KyZmYMcef2/YIB/7bk9achYPHCIWVR9LcAFBo0Osuf6+WLqm+MZlFWQ9Hk1bcslaeZrnnPmR
1dovKvb32O+/9IkZ0OaMJ+XRkHarT/dkMMRtrZRNri9lnj7NiP8ld3yTG5RZECAMScHfxThf4FTe
W9TGLlrykbyhTJYBMrJ07fSnEzvNTjPZdb0cqge9kHfZAALNbtcKv6qXh05S8B5c1bqNlNsxsPTJ
+1nZ+A82foKHskd1AdKRsBvQVOsAKNkgZepCxtVJHg/y7hA3qyiHfkUTPZ6zhamhGPzdQ1JYTh7P
eeTe1bk6v60v2YDW2rKMESQyb4qzyl9VlgzETLXvPB2430IKqOyYLIVIebzn/Nhq2aX5jmDUiPfP
MJKd3cVKTgfxQCRI/GRCMrf4nfekzivnDWWPrlSeYgLSu1PQv0CfOduHjUVQtnIOG1XNzjw8UPpS
ETBTNVym112NO1Jkies9XdjNMvPfKiYBmdulLw8Pww5nwcl9MFkL3pzyu69vzB6QZUrjP5x4D/UR
e+HW4H5itRBXN7PE2HyXo7m+X9Ny0uxj3v27AjfFLJSjlPMdN4de0lHQ1L4sOfS3oT7Mmv8X5yn5
D1vKXgh7eRYVfyQt++rBGPpQcujoA3SnCxDv2Xw5gqsQxHOYrXFW4Vm3jwwlY+xi2vVqyvqyhNuX
Iib6mO2U4RHmVhWlc8eyUorYH2+0aAQytTuK8tacMGQit/L0Zi7HbMjgxNcGUeKd56LLpuuG9hb3
Xd6izlB0v1g2+Ni8V6Mw348iFxaBdMcefDiw+H3JvGD+sLLeOZtnhscaIpvKIySarSh0aHDBNoZz
ShFCUe9Rl7HjpycY2iDlGiV5W44pozAm7xWOvIxkFlyPcSjr//7h4bH7/rsIEohiEAivjkR42SYi
dAbrMF1EgV0Ybn03x8j9QBIMIiHxZEOXRpgTMlJsKk6gOD6wwwFAhkDOJJwyXyVD9aMTUJShLg4q
m8pkP5p72r9usv7PKX96H2x9AJxaVi2ilGyU+O5/p9hXOJUPv2mxMpAjqDKYxCmqxPttRYJ9mjde
6RE1On1YThycLXJBGsG5SxZTGo/jdXVupstuUyzi8KWgxFDNf+l5sY3XNM0d4YR68v0WK8EpRxV+
RLKur/DpK5Ij0yW0s7N7RmTjscLxt/T1ti0d1CHOhkdQOfaLGW9qyABzHamusdjW2yNVvogQoD7y
KvVkD9AbKATZ4WlQBJebyikCrAotzMUibmjA81Z6mToIAX5p2dZpSfaGgAwUoQma7yf2lDPlU2zL
2z5aN2Kd84yzWLXmQP9ag8rlLdL0CxZPV3RSJNcclv9JmwpUYM5tTnvv1CuhkO7n0Gk5EYTDYzdW
Lba+tr0G3jXtFhwEQrH5gUROA8N10l183AmoXEO9KBcizpFsymxSKeKdWiWXOwxgKD2DJbuw/3lU
L7OwFueXrMIU+k28qJiQ+KQN7oM085cAcrmx0NLtGp4AzmSPQnewYqoXHsBFVwP704fD5YgXeJJG
fMD6pRMkQAOrYo0XP87ry8SvOTa04oAbZ6IAOaTSLtBxrSY92kXECnciGlGOhX4BJPt0vwOZp30N
DAFQ7cfFxk0Sgg3PTs0HAUgS0SJsXs2CuY+rZdPeRr7h316hmUdOCZncFqu1EHZuHaY7opXoBvkH
j3vVkiTT8Em7pKsrvf7z+lQrdQyc/8hsBFALE72KXw1Za5u5D+rBhlpfkrYlp3atjg5HU/lj2FQx
05j1TRklvl3z1vbiMs0s24PqzyocO5f2l++dmgSrEgazgrHAugHTx65uPEqegjnjho6VG7pNnQmX
S4jXnfQ8NttVPBmPQg/G3eMLUI0ez9BVpw16MS8Xt9nLGG/ek1cXhoh5GSLDCWZ20MNTHgbF6kFR
P4YU2VM3GAipz0/CeEHBCmw5TLdsEGjHQnBKhu2q84DrbZEKFguc3Qrs1UcbeQboHGciNDTgYGwf
PF4t2Oi1zz1tsUwvLrgWIGvUXGaDD6eorkK4A6yShCU9NYcZSGhh5hW+1LaKtwl1/Y59Sy4lPa3k
/Coy5eGcdyM3IBbMkZjUniZqooX3T5rrztO+/wNXeMymz1uOIcs5usRQvMoMax/h2qtnBHMqPFoQ
KOLmGOeAFCRbwiwHUdKSOSKJcampcviWQ62lIWHdF2ScDMwlVEtdSIYznSvmtxLRteXq/u7dOp6/
yrxC1e0tHdSoQyobd5fNjF3VDRmYH6sA0XsnmMhhAT6WUjajqao9Bz9x+2Yk4QPF+ozLPqgA1bfR
xX5F+IhSPcYimtCtJcq4DzwzBXKZjDXR/dGeMb49WbV7fNy3/ARFSDCCFKxDzXW9LS8cTFIjnjdY
orzbL+NhI21RK26j9cD6NqyATbhjXVYbc+oR6AiLuFKgjnBs/xSDtUlwqKstgLiY2BsPwBMFkFAy
Wosv02LvFHXGC1ORTUL3f1zmWmQlEJjl5alh9l5/7YLHN6HTxhizn0hkSF3U7ybG7oQ9Gy6K7LCX
aBkFuLz6uQDzqYcQQfA7wtROS4qiUNtyKqx0/MzFCSmL/H/ddk/cqZLH7fv8k6Px5m/70eVVNeCY
5ttJITrPYxK12qSVACv09dRXjwOrAEKvtRP8mcfUXzxPFJJ6luXO1jba6Erooxz8S1w4/duHfb+4
XKIsv5rGSkNJyqaDZTl83vUMSEFJ05cV9aKNnHEXA0n9bXAJj27V14K7f5sJcWEUeHZytEQS2+Tw
HZaM/1UjuYaj+JVsh6Kf6KoqgPXn2NrZdSsXEdeDgPnCWad+TD+KCeGMjGbm22YHbfNlWn2beee7
0/j0q7aNa77+ui+tIYnO1NlBJl+Hjb6euJ2xhZN89KOghDigtwsaZbZSJgtHAPipUMcwvOxqMnBz
IXSAZhAQgIeg1ZVDB7dTk8R3CoMuWArEnRe74BOW07HixQ1GgSbUfo7HAQPGZeYwyei0t4HNEJew
aP9a/qEKXNTq0pEA2Ng4KrJiepQ31cuFyXh3ExiKQh9FuC+fOkBJURvBojelOruaLfbN2vVuxxu7
iKlMhog7Itc8jggrNaWyevs06Byh0GW/fojQo3UegQj/RYXRNVZbackZbrZDPGUAhZnUuXoP0sut
Gn1uRTsnKAQ4xCJeWAkM5mXimbjp18yEEEZjgZscrM9lLdqpDEBwN1JmdLcLTbscSBbZDYeD+Yol
RYohA7Sau10NAkMQgZPtdn3RMeMXzOmNi5yyxvOEp67+lfMj5CnHHXziLgKDCqOVR8t7BKcbHC0Z
LBNG2bI4sIGUxHDgeOL0rvBCm7ILMbjywboqz5yO61dcdY3a45wuDmENjfE0IF/OyzgEztcp9QmP
CN2BB9fQhesBN+2TPxIEGJv2Gtr+vVEbzAmJ1ipOxA37zbXug/J6xeafUKCaRXSl949Uv+pclHUR
b+bYrHJTvi46Y1fdxEQ3kiCOX4mEqHmYUNxSNYmp+yfo6O43Bxmwb6jUumXd4V1xvaTST9c+7ykc
Yxp5qIYgngnr3TmcLxzaU06l6FehyqYo4FKf4tAAVRBpx7gbklTb7U4gRTnuzL0oyHQdgFliw0tT
nPd4+dXCJyuBjNpWatUN6FGNqmWAWtCqEwcA0MMwkyKHUsAuZTHQ8EIRv8uFU0b6rSmwjm5UbwxK
Jtt0t2j09B+iPAo0Osr+U8SfTVNCk62yU52JenW6bLaXD+U+v0cKjPR8hOnm8S1lDVdEEPIUjoZ0
esTAonHfNRNvm/suMytt3tO3eqDSKtfjtaRjcI70nW6BB7tPBiA9FzK6do9J7Qe+8tHU1Mn2Dk+Q
MFObO3IR5Qbc6acZQsP6hf/uprOIhvxPO3/DckVNI2jbdtCvOJBdt9z73ZHdVmRzHAt5DxEWyRPn
Od6DKYLv6OkmJHAGVJ3+Y/02nRbyDO4HbdilDQo1ODmAapDT5kgniRDsXF+CtxIjis4kwv8ydiPS
f3th+TrJbNkfU763wddTgPTVyoYV9s14IuvMpZhDQcQpAUgxAgFhAiyMY/Qmcmojob6HSp8Hw2c5
dzNzbD8cIrykivReJQ/kwgGrzamT89K3lxTEmGcqX1S12BwwkI0nOi2QhojD2gvkRMl8faB02u3M
bGkmCbUH2J/ejFABkPIUCRVn2nTts9jGENIRTDYjbVJBn7x7uST5zYvcMKhXGW1ydUuWAAzisnI6
zDzF/9fiCcKlKn5/3PsXMDKxlgyvsufiP9KzPiwHy1J/z3RpgL/WjTNim4of8yzzNxWyEJWdqhfP
oY11OEeV+YpmmliRZqzr5F9SSQ1yp//f/HSQVgqjj7abSVX1N95dmk/oVA/OJw5m2hyioRl/nlUU
N3PK4GG/C2nzXY6JvAOg16qXHjTsl4HMnkqjzVLFZrlEUHV90BCCGKg+vBttMroYxX1zselCjkkS
q3s2SrQodrx4swbN6A7ZeWLsMaNKx5mrhdTP4CpvRcZkTGR/sG/gRyMco209mTASatr/ZDDN73Og
mNCJzI7a+CFhpvGBFM6F4I/8N6jcfpa/Tss41/nGT4S7sfYjKJxSS4mxTbRmm7Tt+GLKOXerZIli
w9QuQwj/A8ta/iW/i5OD21hecQrvSJJyNve31YP9Oj6NWpwJWOtbI0JKPBKNwjhDlaXCx+f+wvif
4kT4qNnwfQcHVt0KBpBeDY491VoTkabunrVCB8bAHwvaaoZK2oYosdw35k1t8EWTo4NrndC0owne
8M4zJSmoXP87IoipfAte55y+qgZUZGfoQnFhTuFr/2cl7LLCbZ/f1TEO1DyqjEvjlijRU3Duey7g
ylS5Se5AzEk5sFgdJrOMDBebBBkzln+jdMFT94Uvh/rMlzow2jX+oW33xt23wyq+Jr451XqZHb6m
ld11cOugroQxYVPiahEkOPIH95OjzndGahlYjK4BF1+KcI6knCVhobw1TfXgVIZcAkMRYKBZw/l5
nUWGueKsJHMYp1YjrCxY5NmgYmi9hovzbWM/Sp0H6tfbwf5LmXqJWH10AMWyQIiiO5lNCbmdiabB
pNfHUpgaYXmCwzGKliuBt3mp3Gih1mGOO+G9dL/pwRe1QhLd87GfxvtP86rQSd7YpskCZmq4qSsT
RXPLgtcmJck0kej5mbs0VQYsfCTpNlibR3USnQYDD8l/4gDOEzWB8Teu42GLf7dyWbBAJCajTKPX
kCYGPHae9FvjnrdL7U1XKhF8BQGoM/XOBwMQN4YijrDqpAjhs9JWu5ZCfjL2ZCaD191HaIzm981D
hdVBYIRfmdoeOIBFvLQJZyBuDM+Oz8z+SEkdhCL5ofUyd+y3Y007X98N2APEwK35jFyXKg5sWAvj
s3IuxeV3LOe06axkl7AxtKhCSbK5dYSEhAGYCKUYM8ZyUx5wd0djWmBR3G7wQ2dVNsOvQDGNwiWT
eaT95QKbAtrJ30raMnxdYx4V5E8Kb8dCaiy2zzkGu3kcubDKVTHf2CqHD9m1D8rxHtvK4R2EimRz
NMOUrvRWuxJTvtG8l6WVv3Co+2CRJTXYbswGoUIXm2jTnEjqJznLH9I99mbN8aK7BBhSZLxNEOtC
gGdcShlKm90LK/Ahqh65ULENWFtblMTKDSrwNY3ziML52r5pRNcZZ2ZbmLV2L+U5Q5PNT+SNdoTI
kA8nMXY21b/XauaTzpuUtM5KFpa5kjLJ+XUCx59WXwyEv6Dh6gt09LHo/VLoMSgzo1HDg1RPnnU2
0lI8iOfcevFdB0dLXrHosBX/CZ8fUwiUi3qb56uw+7bHUM9LtyjVJfsJhFxVnZmI5GA+N14LyOoO
yKs8XWoCi9ZsvQA3Mg7oYB1/HOH2FVx8s78EBm1rKaKFDY6P/it+B/X4PsE5TXAMTBfTmBr5rlgm
9IKst1nUQARm/3tWKj/2EDAH/dkoC0PS9CQ4trjvp4syK2BHqVKiiJ5mzPxzlxnq2GTSN7s8Dbcb
n4nxoqIM/c+amwxXAYdZQWXfpFxbRUhII4H4WatH8q4XjcGWdkIpiqgCLHKCyFU3KeXquO6HRzCd
2Ghp+ADIkHzTn7nKg8AX4pVfj/y/8LoAWUnetXTaw7gBcQ/ma/sMUm9meATPQrPDVjKyDIHLe6Y8
YJ5LNtr7utdDD+tcFt+vUKERrJaShT20TS8YY6P6hcCG99oAPjS4SsVIpSccJ8ROT25Od4Wal1Dm
ZC+1GizrOmdSJll4hYsA1qmJoMn6KatxTNdE0p/dopH/pykxq0Rk5LHzrKYsvikfHlCPiBVwJelV
lcQocKInnDXpcHqbagBB30/PJ44PR2z/7E0WX819e7JOdbnAtGex18vPayO3e9H/pPRImKNbnTJw
SZJVUIw1fSEKIBuxFHimPVoIQmcMzaQ4ZUWY4ZEyofDBC3B0UMX4SVVZu11F8jIcb2ILWuld1jJB
V98i+4sHcbwU+RzJ0GN6ksN0E+qeQmSYmaPJFqEqpu6VXDPKObb2mQgTFmepQYwkhZHXs85CAzR3
EPKunK5ft0jSzgrVHICBT87yAEdKKzFa36ODz0I2JD5G+wGfB49mcAvRnpbhEQ27HdzEzQEI30mf
UFVv+FECHjzBJJUnaxfJ8HkNiWzLCAnR783DN9C6aZo1Hi+hnRYJv/xdR/7mPvmLt9A6fUnzPRWJ
GgbBLc8uNN+TrnM2CM5182bKw7hKESSjt1ss111LN79w7tWtK7nMU/ivD9jm0I9KVI97/HFI4ppQ
jVtLe9QBSpJ7ZiJdnEFVL4LYQz5uRpHdQ0+gM1uJAmWFqv4YabbVkllUsflGl4MnGKiAiQEaj/l/
xS6hBAf2C+l+UJ3yAaIiIRl1hh+eSXzh+Hn+qyRgfW2kSaotsJ5IvTvep4iD5/nlKmoPDs+51I7j
1qJkPn6NEjJR+umHzh1F59b55CJHpSlfCNkH9QfEGUvLCARg9ZSq7/0jCuPWR0A3Q49276aEoVbK
RpPkU34eYRypbGMmhWsjcELRXvTse9WBNDEw6sQD2bAt9xSFDsxGmbxCFkUw9C5bhDpOhIvR7O5i
SNcmr0wOXiD+maBu/b46rSyE/BFv77Z2l8WPRKjs3bvWFvMLo33cu81zcjz/qmUxLKcPifYc5tDh
+kr+znbT4Z0Alhzsp8qglve9GefXUVKr5KzpBEu0O4UQPEWoSOkMsaD+HLiNd9Y97qSS5hgFesZM
YIb8L0F49u+If+W7yvT8dvSYbqQOR8nCNnUbWdLUxY7OmrSkdSBZviGAV5z3+2CPpBAKWuG1yCoI
fslG/PjnJEn2/6YpUj2wlgWE+QYKUyp9To46eRdX+iOJbgcLZVTN0hvZSQy1smgGxE2lzNVzygt8
hf3RxeZO3F9AdrTOavPmgYSKQDPs1JZ6HcDDQ9GrDgef8Bpthn9bJzct+pDdedArM/TMo21BuYan
Q5ACgccde00XKJ9KINxzAbwmijS5lxtyLyUNzC2dVREu2KeTNsaDxxSwpD4g2Sti+xmF2QBkQVfh
54NVRWOHSPYbU1uZ4DujKM/KzvNthXx4GfSyh4hb5m1/p8ObYVwMkj4ZP6d11HHYc60MQDS5c55k
xRHBbjGafzBnLM4Lm/vL/N52MDYDdgJ61Mo2M6sex139o/WolZkn5enF820H50RujYeGC+AfMup8
FOXzPfymLA/BxtqbDM5LJobSkoLVx1avIMWvB2+DwEoq7k4vkRcP+lai8ZNH9yGTBlwqPEaWhztt
j2e8MD+gmb2wZEd/ZNVSMtcl9m7P+Y/RjXwEsLWLqGaUK+c0Bkrfw6TnXOQOjKi9jsVnJeb/ax0f
4iqpYNgILDF1x80sqVjHqAb7YQ9RLXs/+B/NP/h0y17osQ+q78r0afeSPYSvlEQc8o2XrAp2TLjN
O9fiFLSTD0UaIrPmS/+G0IZ4GIOzhDRCA8MldivcXID0j63BMezsSjIxTh2xATFRYI677DvKUZTO
1rmRb6v9/iixPORQqRcdZM7YnbUDQA0luXjX067tMwrtDp5PN4baPh3zbpu4PTAiKQ4rdehvzsAQ
8bEydXo9qxVk5iDMXg5qR9Ite1j05IRth8rwjaFPiJgXkPrIuzpMYkoNMri9jYldtVALtFQGrKhI
0LWdh9tqyBozO24hDX+DpOg8w1F/qsqqmbr29HV+/zyK7qUGf41ssrfcvkm3BMRM97xsRBXgu3Wj
s/1JDjHELtff35cDyPZhdlrqnF/JQjCRMnOTw4cin03qkmzYwUSH0mnnIjGbK0xYctRarAFab0/E
3mWVqsYXFExcEFvhYdOEqLRIInZbvfzoTigc/phgtIM0UAvnZ+e9ZvU960wMA4qLI67uKxPk/CqA
mVY4kpOHThVm+g0FHLITTwPhJk3naXOSTeQfQb7k9cvG2kA0WswLN5oHOqwAaI94GX215Vl+e9+o
op7byvVekkvC/H2hjyBNPRRy/rxGMEcNX0+Cp4XzZJimQQ61PaDBgcRWsiPj6RpA8YDLJf+vrRae
10JrFkvUJtcsjpr78AL+pqCmxKSqVm7hADIrJcaPKqLhbeZocJ2zUIeyGDQ9K2yCMZ0BQObODLfs
Vz4rixE6IfRrK79dwD8WZGp3oZlNQlRQBXQ+12mveF7ZX/ZnxOA/tWj9bLArGNkvv65XhsGg2an5
5CxaTSxBR/8+QA7pprPdDYRmuJpXcX1wwFvgAWeIrdUkv+YoWCUa9YnT/zmLkXXdXqcBfCoK028i
RgUf2/3IsQNcI+Dj+iwLayIViVW5oJ0/gKCGjhuk9QgOjRizZe4DJZzDQ5wSQXWxRGt6ZRhItTgV
jpGgrt2ekSKBRXTRhf0WnBiwwcFziyMdGVKLrF/VkC0gQq1CrbCpIdGzGCRBEtXu7OWAmx2fQYJz
jKocx2cNZBgtDlxtzgo2WISAcD6AWppe5w08Kyol+bFNYBng+1ZDoDfB07NXXzZ+/rmlcw74MZpX
MlubAP/iEpJM/YPptcKk4ak+K/zmdkYKLr7xnxjkX8jxRE2vDA415rckNIQNKQ4Fa0fKCkF+vcY5
p811JCpq5GMRvwZlOF3MZcUENcVdNS/IoFlAC+/2sTRmn3GrLIDLVJZRlnfQrHsksHzwsy03pJAt
9/EQHPQQ2ld3onR6n7hP/wsWwgI/b7XtmdpC00QyZZ+4dkRWqKtP42IL7teewi/HxHabvqWZMJ9w
JLUFDlb7jXkRanQB+WCV0xSAJU6WFQ2p5a3uk2FgnAEM9kgqDUcpwvyyn7ERGjh2M93lLyjC/Mev
Kq31Fp2A+4kOCRhIZQ4hOefZjmLCklg2h4mAxXXpb/M+HNQ1HQLQGsyHEYxE6jlFvhYZt2f/9sz+
riVqAuzskwLisAhnm7G50fcRbff0ix+pesSSfWIK5SRK/gQvuH1jhUqE0ikisvIrYmtm3f8wv9cq
hO8FPcb6BADgG0qfIBEynUl0W2jXQ9/ashBxMUbSgNg+dr/PMf6yKe+1M2s9lAvPUCiIF1UsG8C3
fn+2SgzUPZMIDWvQwbaGwfBYS4JOKrrLYwk4PR4L9tuT9MFGIE7Y9PLkm6wr9OLbTzR9rIT1vuzN
zWz30CA5RFGPdH35DsjB2X5JJu1kXO2527YZLyhFv3nMrZlVPooZdO8bSwaOaB00p3F4pgPZcA4i
qUYwPfNs+dR8j4n1uiEkbTQ23wpKTBqq3MhJkYf4BEawOAlo+ulWatl8MgFRdB1gC8vsHy3hckaq
u75IPRxwjZVboOarmoLA75rRR/YJPuR61ClFAabdtXd9dcUL5lQYFW3UCD7kHeEbFMozFdLPD21x
wTwBZmmrnMjUW782u0MppVOi/5dG7LPZVg1DbPkgC5HuWj6qsm17ci3RwCkiHCpd0f++5GswHvoz
HBgWB2/9JyrAkuQdq3SeeRdUPwzynHFYCX7hlHUm849lhxL+Maw+UvwEOpgiSOifGdHkkuS5bxHZ
3gfUUyYTkGrpEDyGYKguP3QBv2DFLrNU3upiiPmzEEHw52AuBxgVq6DTEDhqT/G4gGEon/hWfmym
cmWt57RYOb4XbVQtphMzbVCnOpYWpBgarVohViBAP/y6YIexSQzT3u2jh3tRU/boV+JF68BzM6/3
oeBKgUMcC1C7mTbryJY3o0bFPST6RiPQ8Bgm3yVETxF2gRa/FLXxphon0W1f0TiMdzYX8sK/Y8mI
au3xidp1Z/GSFe8tfk8PQq8UusBLZO68aUpjYyLrSJnFNwiojnxt14ZJ1QXnfIMTKxf3idvxoNCJ
/R4SF57Gbn+n5g6FHTsg9MXDvfJBXVJrSH6pacJaPNFZ9UW+Yk+016V3tT91ieDXGQRJv/otAhQm
v03Rm/kvVd2WwIzRA5f+qPgb1GWEdnbhMTTDhHwc+0QNzyQRJ4xaGhhYeKYwUs/CPurY1/czgdwG
UPBLkDJnRjYsDY5fprtrgzhmzrvRs90PJ1/bQ0o5TZL4YGK0iMdVwJTkUb0xg5P09tAJfrRFX7KF
rCt4oxhbaAPVnp025Wkr1iQa1YESkv7imQLaX/UG1iMa3VXxiCEcq14t5DPPnf3hxpLzMbQ9bgOS
OEOrrDzQaL75EY1J/KjAL0UEg21lCP6So0lHJZWToy+c0N01+Dmtc1ryfJEfqRg4cydTf09LjyVu
sCjARACClY83+xyh1VHPE0UT8UCFdc+NzmBBeHZ4gVobwKQjbDL36tk8DwZEcHINGMKOA3i7yMP3
cQXQzU9z1cCdChnVFUG+5lMBIGRVfXxqC2pDof7pWx1tI9aCCXMYxsutRgKXNpNuxb3qJEKKVXqs
HEJeiQH9qS6siccCZrXE3RB5UcaJV6iXMHvw8T84VJRkrD9fhM9adwEPoV7kuIprC7jubF34NZbP
bhx7mbSGxfbL9oeMWp0+diPEDoqbFnHaUA9XXbLzWiVRXYzVDQMeDrf7axoR8LmUfHLv6PmCzCgf
NZvDGCI35bysUan0PgCFC4UgHzrWszOHDDuQFQrXfUR+XYpbrKv5cIZiGF2RjQecXJjgtdTKKXII
I2AGV8MytYg/EZdyxmsuQJksGnCkvWhWduPg9DVyTBcwemL3mXh1Aqj4/J1Yqc07qfSgcu15VnOd
iYXgyo20fOny6jtLTL+xqWaLAHNBfhL76pGLf+csJ/Xx8QHmCKJMDNbqjBTTRao9THVOqskSTTQA
0UJR38rJJFel7EgsXpAcHO2/jTGNpjL/fyp4FSxXLDbeRWxSGfAgbMEqi3aUROGkd7q0++asgQuB
NLX1nmDBsOA2hj0vMXXpvRugl5q6e9ismNvOdLP2mbHRqBvwysd12ZgRTdLcCYW4SzTeyUA4K6Eb
5VLRrKcEIcMal7E++Slkv7T+PR3bLGiRxZJi8B9Zj0b/Bi3XU2Zgn2jkR2IaPw2xsG/IdTJrV+mc
EIL/SDEtXT+3tOBQRl0VbArq7C1XLG0iZcq+c/BhJWuwnl5Do3mTnfYXLmQzZ+L6TYR972aIUSr5
Oq0uSO8JKD+5D+OahL5qPGhAVseXXu4iB33hI+fGoYX2AvdFxDe8UrVnwLzBuale+yvGjdb7a+dK
3ESYfDZyiUO3kLcAz3iNwNgsjdf283vjkcO1YZpV2Zc+VK+9gayupjkhIQ7Y5NVeLTqeC48UzzsC
OZvowIGTWhEwQFhsLmPBnjE18sCY7pcvBxMmKeYCckbULQorJzU3H7epYsjnY0q8ElfFkAskuEfT
p6k2wx9kLJa4ujdJpyS/kxPrOXHIlwyBMkZUOA3Uf8PtwxR8JGa5pOsia61pm6E8tYxw4WYFx1Kc
gjFyA+9qBulFtg3soZn4UK38izU6ruBSIa7XMM+JWrhB7r8N9gaBUZzoZgW/g7Aow7nVDPaed8yy
s74TJyQrUoE6uQ/NAhQQG7DETq4NpXAaA9CHbVvTRPN6KpZztypKDt8GLWWCleIot4L8S8B2q1w0
flBwPtvbfyLwB18M0osfCsf6OoQboG4wGTwTNRt6DuXT/NtMCGW3gtdX1fDPUju5C0jWC8snY8iB
PcqvCOqucBzPzk8LUY/NrKrALgrVkV1msqwz0dWxyhuq1WQGbcnRySA5txToiJV74kdeA9h5TOQR
vtuEb12a4Nx+SFF6UyjS1U1NOpf35snsXcZEATASbcYr0fA56JgRJwz0eDVO2zPLIYK+ZDF8xjKQ
3KfdwCDgHnluSFzlF4bFneUfcoRoQo36mqXk1auTla9343uu9IzAr7zq9DH1DDv/LNS9x3CkGYkX
Bi74UjMF6zttZNPwHWVoDEybBkKtdFfa2GjgIP0sXcH7pbHIdORKCmpI1FjmXj6x3J5w3884xvHR
0ZNZPTCoyQ715YcTuyUrAAsCj1RZaGIZpa1SwHtJXA7m6nnGlZAKt4ln2uILtdLWBpkhOdWO1uFH
UX24ny8Am/DHz0HMYShmnHKar3mP5FMohaNAFnpGGa/FDoUmzB+OyTs4urv5hzqNyNGeveu/+bVX
wfN/2x6bBNHkuKtbL72hb4KolJ35Gf77sZjSta+QnTUbG4SrSa35GlYS15WNoXu5gIgcYoLESWrC
eTYAH4V3ykfmG5siPL8ZyPqyMDu0jcqT6lrTm+XeHH9MqNZBZERgy+fHyPgDiZevZ7BtTLWWJVmB
Uwxw60z0sFMOz4SnYInaXxW0xDbVNasW6ta5MD8XyJ4YuxcesQ0dcYWQ7YpIzMbfe1AX3/cCB72S
FctHtpRbsAOiJVwwj/ElUR9N66cmMNaPqZTpNKJSrGdQ5GSUJVgssO1uqyenV/tlMNyoiRaYGqf+
WBIMQMz4eVZX2Dy645ljm76Tk6POkx4meZ1zzzx0oGPBlgGk8xr3a2pgIYPLMBoOYhV251LtpkEE
tHcwOihzrNMJJaq48lYfOeI9J0/BqCkuH6eloHBWe9KCM0CujpFGgFGzYgc/n+B3k2ryOtdF5hE7
3VhzvtA3qAGqYaUQ1akoke5oQb3qoq9bi2Am4sd5L/mZ482R94mYooPpLJf5OP10MlkudfO7XDa2
ILr3hq/PuqWD4p3avJPPIbnSfxrD88MZ/ZCGIttcxjgSXCrhlgTmmBHuOYby7tDGXpuLf+Gbs40U
cfiSiaOPMgYUOg1hywseHiT+RBcjh3PZBufKRm4J6/IMLtXgd91EHEe3vf3PDnn74MxFKXyd9MKa
MK2c8Zvdj8PqWLIamr6pdpgYLqO8oCQdRWRdBHH0uSyIdWKOQ727NX8HBnHj6XewrHtiy+YEtes8
tghIFddzljRch55W5MKqgJoLTOUF6A9RpZR9HbXffTf+Z07LlLph7+kLcXKnRfCXAmc6IBwtjyfS
+xG+jUlKeSoNMIl1qsHLDHWvqjGM1gAFkB14Pk0obD9hCOJ0C+ZCfniamj4rwGXiDLD4eLhBVsVa
6ifN8kQWUWPWsibQ/0tMHLnxzuxhI2oUAXS72uGD2FBAuUM4/F0yKfdyT4p7ISMp2PrQ7ebPOSpc
SfV/sGD1IGvvZJyO0XvNkSlkYKGCdQfau13ihpbGpZr43OdTLmrsM5KehGsKRqb9W0u0JK9gxnUB
KkQdhKHHugWepyLv1G7ma+bkDmp1EYM0V6hHthV214HLGZdR1FmNTsOSymHUNnbsMldTudrj36D/
RmOd7dGiVZJ8wOiDuu85LpsgMRRGqOsibwCn9lVCcbP3tcnk6hmaTkk/U/QoAC3MJM2sJpWm2lif
7tW7u6AqpDjGOLGWzEELxRkQgV1t5KQHjMwHKD4/Y4nvJWrT2tVL6W8NnY3b/K2N7DWfOXWFVDe/
zT+PSsCHStwyJ3v1scyZive4DVfn1xWJqFQVhWId1hOrNDKFLgCRYrR0VM0KHPJmuCMeY9PsWolP
eWNgUWknY9S+rs5qYNTo8Y0cnZDppucXuV1CVPSg13MjPAck3XHPo68JM3Wl576+dkuxgQm9gOeO
hSSo8+8unf/xO3xVVNHXOkxyYqyyETufLiYfIdPRE4KfsF1iIWIWAtPmwEYefa+PAmsao4K8MAxc
WS1bznKrIdWk9YfyOt56s5YCBS0SEo2LDVcJV1zs4ryiRU1Lf5qA1bCpBX2aDKz/6ah/caZhGAFN
ieklESNgykLjs/+XbQzNbWMaCanlqzyKnfu2yX6ZFuG6qmlf7DHKLi1popG+heZmgdt9KhoF59N9
ngNrW2CezdiQ801NFFO9ANcVl63kzMZwcVDTSxQ9tmRNVYUUVrGx1r/tUFoUYKEHkxpY1982aIP1
Sih5g10rZZ0+LTOhOqmGEpv0tyLNQ75wiFe09zoKMU8AhkfiW5N7WeR2pMlOBKC4FEd9ytcu+a6c
Qb64xb1tPvIX34LWztIBZEikkQ/dieH1iZVdGRNCeTsds8TTB1hjO8BKccIREx+1d9tkp3ioBDRV
22tJQp2AStzkDjUmaMz78qyuApfsdrTC72mohqEbpB5/gsU3YY7hSwz9mw0j8YwrlQbDhJ0nfFqk
IYl3GN3wwXYlaDtRSNvt6qvmvN5O+ksOsJScZaxo7sAve2ejTwkan8MXgO4sNfnTgtC4rxTAq6bS
RmIxC1NlkqKzTSB6R72Eux675grDInxsVa2ZoUgZVsybXTy0QiB+KBKM29WwnoBgGQPRCfzW63w3
LuGve3uVMLBxG+t+afUewurBW3njR02iKmX/LNPw6uGikaCUxRdvuTFHz1BULZRBWyr9phJt4mwN
3A9yXW4DGf7mPBs/dg0KFpo7zDMAq7uy7hxSVos/dXXIfKCwkq9vNfXEQXFy+njZP155rNc0Q0Hc
oQF0zD7c+TLGXYmFqLKSzvv9/dEGnxoXGzwBACJVa2sGU9B7p3KH49Ns+QzzjrJ+xgTvo3IJUfrM
xQq1H/RmowmpsHOorJGP4UKKksF+3/yfdehAAB4oIdkp9UffJYVjXwDEUjZnTKsMFZ9SfR8JNb0S
4ECZKkw8AS9rgOkYt1+Jv0oejCNGVK705B880i6v+5QuUWrosFp90UChTkX0zaRn3riP3wq/VN88
eeeYom4JmV1dgGPWcuoOuCn775D9gYsbX+U98B+2Dr/9jUZ5PfrRGMKw3c1VfOvNcvbi0//LRmae
n/5kcVIy9HXtzzK3EKcgBUDGx5XsoFBLsDvmkFLMupoWI4HXS2LpWakbSPgxBVcH/W76TGcq0B93
DXsUl6693kt1BfkForDTYg4Tmj68ehGUKsklQkG20iLRXvlytRPZMMZfrwwfAQN32/wICj9yZXWT
ybBsRWGebQ1T9E3b6l6EZtMUteWyCvsRrYJzyN6nkP2FMLDkIYTz0GSaf03seNHI7rlGRkbkKz+b
s4JPH9Q3i9OeFXwXOrYaWDvMw1AEAlMWh6Udsf58w3Ur0+xO2IovK96nNZjvDijDUg/OrjEVOztw
m9emqMfLT7ip6JXJ3/QiA51k2oU1XmRViglEahgwmHlhLCIznbSWPJn9sDYcDxCjZ+o83cuaHy4x
G1Ww8cjieiMyBVW5zCWqFdQEiN/K6w0C23VYWDFe/vgOpGXVhScQJupv3Vyf76aMjMZXGZSSCW1u
LAFKRs9ou1aZ5tekgPR5hucCZwHU3fDSnKSBdvTW1QYeDHaNBudCq6/3LBKYpiww1rSN7vcWISwe
GnFCISLdx8NmbFzhIDIk2LtodYHaieOBfkAEmzMBzhU/0TcpHU+9Rq5/nqsul6HY/p9h8QHUOauD
VjOybHqUvhpH76VG08etwngA4UNt2i987/l5w/iUQWsb+9uPRoJoObvqVXKT9GiIVFY4okoz9/fV
aPdHYZCqDf+CCxaIaNzHYGCkiBz/GYNYg//JFIfMP6y2GvSl7NybdD6DsgBvifBoXSCquPr7m+Rf
smRh3Y5Nv1Z04NsmwDuItlmp4YlVEl96Xc/BXx6IWflXpsl2qEyeHkOeCuN5DvudB1IXzzWWQqlW
UZFdwz+oKSs8hGpdTdMN/GsLAEqdxV1RxBKVfdAbgDaTlpjUD4Y8vvt3/rWrfVacjHr6qHbrIsgy
t4AxiJZcrHJsvF8zyR6Eg1czRRBtXZfilaH+JbFS4fEU2Ri5n/5/ZWvkcbFx4CwiCbOl7VsB0Nhl
gzoQTaZlOyo/3VnTUD+2m17D0SeoA3xz4Yq1BClxlZb2PwFm5SIqul5sY2ntaeJIuQ3FzBW+xiLg
jkmPCNvlePLoThS6OHYzWWxzR/kMIqid709ee1c3RC9AB77ghhXFHpg8KXrCkAgHAEGi4avBSKu7
XgrfGTbGLguFse+iFQHsFBAnee/0VLveuhZl8lxR245GPoz58C4DLtzrdG+ao2aCEXbHVsP6/RDk
9xxSTbpUTUhfRDENr/qy3OPrp6N/v1gpa/4jS92Fl4zK5e8Z8rGEtdubExeHa+6MwfVxUeGRSwAm
4tCD6peMByYWs77NO3y7QTbZYQ8d72b8bYUYTB7hWtlGWOJimjeu+KisbLHvVpNoQdMBwdCiG9sI
aolESI495SkrVsVUZWkQaAM+ZSYe55G140zemmBkJKNPRZD/+68gSBgaxvNAZtYNibmhln+//+zk
eu+M0Cqlu3JNZ1fmPAvPVoAFmOTCCPTXWH8bz5QCa+NQinrjnpUd4pzxGm3E0WgrsBkV76Z8nW0E
9UfAYG3mzgDsMgxnPlMvPOMAiz9wIMeU6wA3MIq82BDEli0GIu4iZbaiRymNWaTt6DzCpzfbwrKJ
qoMkBbvHaND6ufJ58V5yG4srHyYQwrugXrEFeMGkk3PTYXq7e3AGKmI9hGRfr0lsdHnE5A8jUGcz
exb2gYZyqIq6BD9RYWiWoDOMVzgz/CLOVlJX+BN1Q6VGQ6R+1qed1wfIZi5IRiqAWpkvljk+4oXl
oTs1qrdHEOIO4UsOeW7sbmrpFqDLs5ZBF05RY+6n7NoKfaFJ9DTOgfegSJMDQzJNKTw10+HH7YJh
Ww4jBfUllyob5OrQZjZhFaZqfCXfnERHQnzNa6Dzmdqsw+HIuvSwjgdZyqTpFStz5VSwOSzpRthe
WVZ+jMKFKUSfqbHD3bHJcJsZzye4zWaO2cPWzhNjQ4DH4fq95xH+fRNR5WDAG9dYPbgEd0jW9Hf2
kb8MzQIxUVcKEb0A0E6tRtFJo9vU7Bn/+V4AIsS+R0IxP86fJVu2/TkE94oFROVt53nw7m+iY2Pe
iOVXoe7u5rIeR8N9bx3eTXbGsVjoSNjL4cXn44KTf0heNhulvVjsdTRvkBT9eTmWPNZ5YVxADHEQ
w7dMylyzeITYKxTcYYZK5MWCD1YWfTb6k4ER6FC4PLu/1XwJAugT3BARglw62Qp2PcWMpM2BvohI
WPVWJRg/J1G+m1PMpDXpfPBGRVLBJxk29LGKCPu97CcTf3tpuIw7tsSOVxeXdD8ozlsnieYnXZjp
aXXj3yIXGaXjzLpH5xBnjWJSHa/HCEtSfLrMLhHOdCH6gJE47Npet7WFgIZB/4Y8oNIYbvnB9xTS
31ZFt++hlkGD3Zp8q2bOs2lYZkvxpQ8Pst3wTmBiyhR4ShxX9AfAIFkpCMRatJlIxwfDkRFvmsDq
Myvuj62WTvCdkA8M1GqIhG/KY5hKBO0DWKprxa+t7+N82i1wcr1Is00BJidYq9Dhe4+2DmrYN5sS
bVKlCuUX86wg/m8OwHvB9CX0tYg8JEp2hBgiASdIZh90LXFKDcLesEWQe2KFyJ20uXTRLRVwQ9L9
z1k37fbVo3DAPBgxWIqu2N3Ar9rAJ66qBG1FnETSLhIsHYeT1YYj2pK8AECd+B59yW84C7ycpHlW
RpyqRbrcUqiWoIZmvmirEtSUu76gGGYdrncZVCldXS9F9NDHwHzw9jslXujxFFwI6h2rnWRpoCDT
DOnbAIs9TLQ91zSv/uD/EEjqp+666pzNT5Aae/tAThaCl5/1H5I3cjapoTipJ07EB0I+x3zZjdmt
C2uO4S5T/alOc/zlFmqkU7G+IoVSEwFoLp7jAvi9uGOpzOkqQAqBGZ39YDQETkC8giomY5iZrWYC
OGQOl1OorDq9r3CUkXYtzmONI6isZPgsY6kycHz0BnDQZ0CwBICXmexN3JpmIqwg1AfPf/jBDUv4
8O8ETpaVSWRXkOfCubd1uJlR4z58fIoTMfcUhIg1XG0Tdf02GYoBwhCJEMBwOkramWjtOlX2LoVq
DX1Pnxuj9ZuUoGfIyd6+Og9f+Tt9Wjg9rxOFF6Y/2CbYcu56PiTvui4aVjnP+xouI7Zmxb8wqK6W
jAReard11J/dfDakT1efhls7LcvKcsVPXkV2Xd//56dy3zPfQ7QTTc1IcHHgfUi7iN5Pf+OQ4Wo9
pepcH0L82vGPdFE07LdQPoT+mFTGe0yNuHMoFS7f58jxImOkDKcyQ/3g2A8ASrSblvQXlO5vd0aB
1PrWCU4+woeMOvt3ptyTLt1LIAkK8M+9P715AjVqki+vo/d5jZHYjU66V6kPit8APUCbt+hhf2t9
0CEV5RRt7dj6RALJezeTMty7QseHIj4scKglzaMEV7I/tmQ/Exm4gOcYYv934mgnoO36QiC6dABb
dfkZ2bNw18boH2kNJPIGwmblaKHuexkQtWaAPkS0vS8VeZsVW9xGlmvjYXF6qth6f8ry0dRMVyEk
OZIdZZlVzLlZsohS86rREPZRsDZv98KK099ENoVCbtp66T6lSiJqwWBM2A6zp2WHCHdYTN14YAaF
u/hdqtU9w0gXmLXZSgetVLktXObUDj+Rpz4ESlbw8OSTBL8hRm4VVD8rg0SwwtBmwndjEsonvBnF
Cw5WFjPZmsiivXGokAKqSDEg2mS36qbMqWc7eoerPKkVGYsdGL3+G4NHWjGHtH3zFArnyG05KbIr
kToOao7UniOGn2TcbRw5nPQzZeC1HjN5xm2GwWatTCJIz//GL3Ir62sbWqr54jlrCOqlp01++yzD
iKFwWXbowwjV288Kfx+fcXwVonrWS42rREF5oI826aJq1typ1J/GG8cZgMukimlektFeb23HZ7An
l43L+j7LKmtjT3PhyS5Hz5jMMJnUwOtd1DLDqx8JTxf+6f6o8VyroTkhYmZBeDNQKVfx7V08ICEI
9xi6Axz1KmKdyx0H8lPUmATMJESPimTlLu+6IKYKo607sXiGidq1kToBoONfeIfQVPey2Nz8+ooq
dioHdR+hPSG03R8f2b/sqpw7e4ZBxIFhbArFREUiSsNUHvrEls6xgl7JEXOywfMQ/0/w4T6M7ekM
PovHkB0CuVISUyUCMJRqy2Iir8x6wg3k/VmqAzNnLGwWfL6Z5xApKZRoJKLUlfraVTY4lowKLwVG
Gm8vwvdzUnmMjgvTRkrWAPAfMsKY+6tsffzFZSiS6EhZYHL1WA7S1SPdDXcaHns2pSM+mEefG9RV
fyCyVRs2WcDKJ6DFP0axG+cOm634fmANbJGxNSe258yVxJ/o603o+fytKfFUVRT28AC7/eMFW4CO
00+FbkQ4n3L2aWYBNmQnSHWksdz2ALKd/w1aIp8ktfjcDP62hLlFyJqnGRAy2HYYeaEzEgPAb8oF
+0LVR1sBLSFLsfQdNvvuDK7+USP1Q0OixKhR1aCuPTz7I/JqxpsV8Vnps2m8ecz0itcusBuO1grY
FcD+j0TizWT5vFppNfskndAr4Kni2lGhPkSNvHiUgx39sckrX6OMTQ9c+AcBBMiFDkm1Mp8IotPJ
HA53qPMOpVmJSPXWcxXawlyxnbtUB5sSnjOxKsnDeTEYWDnaP9Od+DQaI09X3FcnFfCCeCtB48TN
CmXXDmY8X6ZKZBTEAbDPnkKej+zqiNJ3RmFJJpAteaFVAtxw3h1El/7H10M0Xo4b2wEFFTV/HEXr
D/rT3gA/1JMpFB1EilIcgtdvZJZpwJb3ZBjSQdfXgOllMSZnB1Q0VyjMJlvSnpXppDR6/LAvG06r
9HPB9WW/z7w5/8Y/V80jP9gj7cIRbccPP+57NKQmKThDNnBdg30TZnNt/K0fwz8kwmVn6zMlDQpV
WIkncX2yupTiF+3kHymxnae/s4qVh5bRP+eytJscOJrHA0f429l4sJTkSw7Ymq7PSlSH/tvMZwer
5wFXmtF7N76N3nZAuHgX9DPcpuQ/1HxKnLJCpefPyjJMNFR+7F08b3HIVzIJ99IyxZGnVdmP1dRy
ApsU0WsuTgDSVuOeHRGuFW6h7NEmt1F5w0jvg99DQwzND0iA7TRNXdglLSZM35J08cv/Ccsbw4Fm
vO/2+C54CLdaKL/BSIdEg12pcyppAxHtVfzRIeB2QIYsru2xVzGbrO5jv4tbIRCISePr0249iqBe
LgdK9NVt1dwcdhMQmO7e35vXOVJtj/XfxtUxVBihv+v5zu1P3lFjY3eOTQ8QRWKv0vlz7pFJZxpQ
GISZRcWUBZ9Aj1M+nIV4b5TsgSRU5LCasQ54HJJj5whgyX5bCxBlIL36ShwI5EHF0dP8ESLLYBfL
RU6ZH8JJEpO8jGiEPwzKhljIH6xL0TMpc68J9y0hI5UyTKIDt4xblRAYuVSd+gdeg1oB6yauCIcz
wuIOHVJDNh/dfMzzUV+1hK3oKzwyhkyq+2u4GbgZH9xe9BC+7qmFMq4k1OnHOpU0ubsolBFI8XVn
+qIv3SunaMAd5XxEHgUiF+q6yldGdlu6B/1HFYqWYWM0qw+6BVgz0U94DXuA4cC4l/kLrbLKtYn9
Np8QaSMQ/tC/yJgUoDlfKhcM5zoQjOnQlrDxMSisspY9bOT/JltsYBmrMInshcryriUzET3Q2Ko4
YownSdr4VYmB1pvWIaqE/JcvaEaWDbZnM0mCXuVIVD3gdOBzKdgpKjUNkOe8Hvh4ugFVDsJOJLKi
TwdodMhWSRJTOWLhos9lp0Ns+yIy40osJbvta4VYYOi2Onr+65FiVcxBfBAi1gQy0SAZv3t6+jAv
eizpLfmDl+fP2y5Dqlwj/RwpQCWG8WuVkfaEzd7NNn9Gxx44ChM6c5XIDt2OkidoGwfpw+btjNvx
v4fq+F+jB4TSPOqn+guKUx/gEQQ2MZ83MjfBOp3AbdXuxyXkqSVQdYJ8B8ZzfaBPV/Y9cLQqso71
j15kjph985hid9sFZ66JuHQfCjRD95UnLVvAka3Ke5qgddlDO5O5DJM/0A5WBzlWHSyvYFten/hc
/OR4SL7SyLqnf7YRI6dpEoEq4wfMR3vvFteHLBP8jA6bonQJGCwKBpNw+G2qC/XYb4CoHMQ3ehY7
vYuh20FlxddZ661wO/2soY8gV3Hz5+6hxwLKAigTS7NvRnFxr2JytxwDGsZlHhE07uJgfArBfiIK
y6nW5YrNTtvSEVrZ/+aRt1cmw1RnDsprqwNx0KH3IBd6+3ckwHowN/6LoHq4r2Xu8porcRG23nzJ
kx6MknWSMVFpApvrkSZP0j2ojRmkgVBB5Fg40YHn9rVCb9KfqLfWkIA51tUoI/Qp48BZUJijlL45
2r3YcELzSJkIUXYZbQa+aHGU7kJdQViyguq6wTmu1tkmzard8vpzuhHOLJXlhfuQJFKtM/4P38Wp
AS2yj6DgF8ckLUEUKvAMwo0OAXfAXbgZ2DUu8z2WHmIKGEadBIybLKj12HgF+b0JIbgpcPdpC6Ru
1/wmgDYq88cXu0gAcAfqUx8WQlLR2P5bip3Uz8ogcGPHOQbXdkxLhVRxiEyJhR6nMAsfT3yGKPIE
8GaeRCgnu9PHf1RiwRort6L/tbxPXgDtkDrfOAHtYNeXjkLsExSC698J9pZSntJQNe/WveC06Ohm
Hf4VBcYDR86/r8PKPsW5hkQt3wmGtFMUkmdZIxuPyxIYxvOS1RH4Kh70klPFlgh7JY2ClXlrDIBX
EskTLX2kgJl2vBIWrS/P11ti1jKF2jtPhlD+tXN1wkEggx//QMAC6mcEuOJKmpVMtDN6Ofl1wUHx
mZeT9GCoRZi9ZBXBINy1uyiEp9fcm4MhWuzlSypNueXAcSOYCNwGHWMoXPo068YiIe/PZinTkK9K
JKJ3YJ/0yx4h7oTi7ksw2OYwRqxqMZd6EirV9ruO6qFoGjgqonfE5naRDx+SMeR3pTm+nO3aQOYl
R+B3entFbU3mg/2+/kIs0RY4m7v4rSrymw0PkBImwGIQH4v3S04M4KjbGnK6znJOh6b5UaFNO4VJ
2xTJN+nJK7dSXhYn6+Ouu+We/oxAvypUg9fB8cUpwABKzUBnxFrZYUKWN0J2L5a2kAeRVsETWVeq
ECxlBBTbAmVHA3IDW7vfpIuE2Wm0aseaO8gXVxoQMo1G/Gw+ojVAspke6yNv0Ods3ZI7Qu4+GPt+
OAMUzMOL0RFwbW3Y5JpXsYCwjXdU8lUAEuMX8t41bdCWxZ7U2tpbcvlANHBGHw//Gn3mbgRfmR6B
/HX+vM3polT2efJfxN3WZP6rLcfs7HtsKf4j+bnzdpmDMf+gRub3jO9g1BnpYJAZCNxnV6/bNZTk
jCGP82/h8JijpxEJ5pEK/1D8dcKFDJcY5k+oJL8FMLk7KSDusTdFq3phj0S53xEoYe785vHbSQ6O
b1Pft+NQ5gMu2JvvVhUSFYNEH2KvOsTLLrh8gfbay/ewje5SbzqH3Uk7E/B/Jp5sbzt+gViMv8W0
21n+JO42RGoWwqGN2YaF1PqL+5RKlCSmWGCK/cFdD6FcUd+1aK7ZPeEB3DMQ27S6HQUwddCYb5J6
Pg8O0orD2e0KGbWnBmuICahh020JnGGO5UI3qARjcEHRxDMt6pwWBp3h94krpYvKBFALCau4sQuI
ZQFrap2LrQiF3Yd9UrpqNlR2XK8donAae9YDUx/a6RbqP1M9OeYwbW6CQI9LGA82u/Z5lFgWafP3
jhba0zTGaBJbqjZJpR2Q5se8PtVQNMV27S69/7JzBqQtwML6aetyuqalfkO39VI5f03il0AO3VUQ
bMeWfrk5eahWt1oGKeo9uwGceO51/EiKXlEr/qw8D4CfIqk1//rUn20fACxRlr0r+Htd+/LOeI8G
BjOOw4nP/DFLIpAd+v7Boo6i+nRl6ZN1ukHE/PVGtYVFwkuJPksllx3Dv5m1z+8ACW+/uqtzdJa8
xDOhiwkLaHbTjwtHrHxZTivy6x3ZIC6chm6XVV1RckzGOk0g/AJZ/rRlKkM6lsJX4r/n1Ucew4an
kxyZByAdL2EzKnNTI37sAKPdPiOsHe8fmdrJ9soY0CVUvQNfyixYyO0jkC8a9tSBo1tt/dNqdJ3D
vZUNEOOwBaYmgBPUS4+ELE/S5qdBxgj+u+qSQW21mmCJDfiiIKA9uMyEcDrnlMkaPnWqFvSIedx6
i96CFpLqaRb6mxdMd85/8U74GC6or6GL0mV4nTmr0qtSiQ4UTSI+rFDsTYYE4JDjQfIJdEmQ7o5P
8nZ9kn8sDW8fLuI0O58zpg915irAj0BSG+m8ogS/JFywYBg7op6Hh0jiN5pdA1DEYAGt7xP+QqEb
l+tn4M7jKufcaV43x+fQFmqHq1/UUW4vA6xVMQ6lzGLI3tOKjy/L8tttuahB1+LoWf9d+YKSi1IQ
6l89sZcF1/5z+0Jk8OkpuO8Q+ygGgMrWf2pFo6k1oD4Fp5V5azejrz46KiuJIgSIf8yuMJ79rsdF
zp7zY6FFPz0Yv/Ul42K99NQv0qx0hDYp/0+g9VX+ABiHsMCnLhe1DHqy4zrKtG4GeC3jHgSVil5Z
wqEWhYugAFpU1gi4aM3qz+ZnjHwAMWFRCHXeAlHdy7AbtvkkgtkUQemxEBMdXrDIqXFgtCmw2ukR
ECRzjodzNKP9Ztru/zAkWKlCc6ysNw3XU+uOYt5HFapGulZh/giXJ8WPEZjadROkS/wFLh4HA1TO
bGvEpwy54yDcLjlsy7qOeZWXzQ+28h9ojkS8nom+wCeXfjBJB6x1T3TnXibeRF7QOZBieGE3nsep
dECtKlJ6tW9hH8K1qNx6/rgkliVPb/UipdkNYAxvWnnukOqYPaolNCV/4eHFlOSobLKBgfO0j45S
haakHBPMUrci6rBnt6n3QuVqEpHjwim0+GEm8L1NPXaSVF59zc4FJZ/+AZnZNSeNhWNk6SDii6Xl
66iorGLg7WrQL56/+S3aTyXsZVA1EuCRpKZkBeChjp6BBx3yx473h2BPe7TWT8otzfGuqTZ/4prU
uEC5eNcwEOIF/bB+lrL6TVVceMik7E9j6FEyRAzrAU7D6TBiBiH9PSYd2/yOjlW5O7lsK4YGYyKE
puFfyVxMHaw0t2p1v+N1cFRKnD/yseugra+67IcM0sh/DB6OCBUkDTbezDuk5vgRS24rpNc0syzV
SNCWRzBCJO3h44t9nNC63pG758lo1LOAe07Z1ZygrhgTLN8ce8mMwjwAGE7xR3GOcoGy6scTIVTT
Gw1UKunojzzR9IG1pxIjjxb+kPvCVQ44wR7ZXIHa8GjTGkd6Ux3L1bRZJ5RSHCqrUrm0huSrDWUy
c/0AjV8SCE1tc/RXJ0nPsg30VHxmWf4QJIdrrD98V0dwdGSNYQeYiWhdF9fNOwiTvC5dUE2yd+1B
KRirl09Em0+ONPFmaetDUedx/2ahVLrVDmTKsh5b795xN0ub1+XzRZ5sRcsqxM+QwH0P7KluW05l
QWQ/anqFo3r3VYeDRZyPdeqw2B7lgC+AMbky0RtmEvM9hHBtbhlBZFWKvG+K6EU/EsSI/7REtB+r
ceB39bikJ970TM9jIR6d6DJi1Z9rntQxyV/JsqeuJiQgtWT6ppU9yOD0q6lHfrhECkYD8j1KsnWD
GS17N5m4CPFT6pEGIJwf3gmzfJaOt8nLlzrxnlKK6hc2kAYTjabscJ0d9PMXkfpDQmcssrkfGVFD
ZN307EJC6Q57vIxHsZpRgmk0hEOQNwors0bwF6tQ7sGfUTJcDQOr2YTv6yhjNQqeRQCfsvFmyqNe
bpVUJ/+uCqQqYZwjqYjwc10rX2vHD/KCMwCDxi7DXMV0bFFo4TMalNXa6AceGWmV/V+ftWaW0J/y
Y/YFDRYLhG6wiiNfyxc7EOHpZcMKiMALWI7UzpE9tqOKVb7aUQ8lLhOtwXBdRVmZKdrK2VUvsQPh
x2NZUM5LD27BA898PxZot6Mym2e1283tOvGCOSn2M8OKETbjjSmcYuYF4lycc8YkpUpQWvwW4nb+
PY9V/KpJeCOaKOrh7TbTtUxIs5uY8pIcRYSWX9qdB4m4F9Vir+4CRupzlCk8H/iv+sT91oOZTT7g
1F69kQUQvZ3UocOZtVxC4ulnz2JHwTyaAsdZDquBfzs1fwkD1fM6HtqDg6THG0WznnHDujc8OA2E
zoh1UUUJRJg5GEZtoQtlmnwLN3QEmkgGKyvoCLgoZIGupF708tCllPcxfHaHFp9cKVOCWbKO6lQ4
fKJB+M6oGBQjhNDVQ/uFSMmI/5S6YttA4JhZJpoJuXJKaVq1EXNl8r7aHvOPl1x86cNaJpZdiqL1
4GARLC0z1Ex1WJrmwoFWyEy8N5Gk+45HM7pyrW7PHgYo8I8VXNECDr1OB4dtb0MChwQrW6VBszKm
8jVdCoh39wvvzvSLHF/pMz93OQhV+J/Th83I0MYY4WkhXxRDee6RUnyDlplafw8bMLXtVVvlb7j8
nKaGXsM/62cCLXa3dHEPmNsONUqkxXnRCecIFC1NINGfBDIizQRoRspdHxr1moel0zS9+hZM5ImG
/DorZuWw2X49fU7YH5N26rmtIlSRq1ihb9uwkZtPm6JK5zf16v+WA/GOEkCM/b2e0KCdQtFmEYqv
9JBSuqIIjVsbaRXLi4OY17mSwaKPaSF1JmHn+U9GQxOVrjfAau5thN9YAG1R/fmxhC/weqNNdPM0
A2+1cMUcfDl5ycXASR8MEyDrXM/uSdMGA2DpqSj26d0LZYIgOJpfzma8NQiQEfOPBNxwiJV4oFOd
lhc7rH2he3C9lJD0I0CN3L2vqMVLMKBzxAhjs/sWC3KVSEmB5odWaq3ZecLBiZrcF3KHQZylpn/X
NQCUHaoZYwxszKCDHMjXFpGr5cq+jkNorhTqH/BsSQOMAb5Q8ev2vVJHkq3ulR2jvICcQxfBtskq
V4vCTMfG4eeJVHe3Akr6yST9i245AwGEhOumYW0LVzA2TqnpDNiBJ2FqLueaZRIyZ2BUaMKvy3cE
4CyMRe8BuO2Eadnna4acN+d0FYBb3ca2wz1tS0ia4Di5ET2sp+r775TPlXiAuFfDt3+jKSl32UC9
OD/8dJV6WKIbVL6bXpMt9FPvuWncRkGsNwEjhpVGg29HkveQgdKCZXkSxO3EwfqrHw3l3q+HFfhO
y5Ydx1PTcLmC/YQ0VoW6Z0UiW6WKZIdX8Sp4YrXLighHKW2YHXdrXYK4dxPXLmcPsTQLvx/Jf/gt
q+4nZeC8Lez1BcOFk9g7C5iJqy2KiZ4kwqTPCfmpJKSi71ok1ZjXkV+fzNpg+4yJUjk13aSs6b+r
hb+ry4wFkL5Zb4nkBkyMnTBNLrzbBape0T6P0J0S+fxPMVqwhJuTFmj8xuHzmD3WDnpOkUg+nyYL
hOJOZc05bsja5hvUJ3iBZ2En+W6uMJgjScIjHY9Tp68exhd+XsjmCkBlE1VoHilbzlIOpNg9WVIn
UHab4weS6Aa6iJMwSy8WjBnrrM2BKmG/RlZipYU63UDg8ZhBDBjeXf4vkrdubKtNgW8HKSmhIMmC
8cm3v6Zf0SMIrbHkg60D+P78Lbb++T5GSnGFRqPYcm+SRMmRon5knsb21PJmHI6a9jautt9yYSiX
tfoFSiHO6evuXkUpA3nmkZ936USoXT4o4P9y4u12qb1ojcypW6hQKiWVFyu2k77myLFEsM0Dbjl4
Yo1cbM9G7uyS865+vK+Gm9wJ0zJ93ZC43cX/NX0kJqIufthHJ8lLRLx4VQZkn86P1yotWcInqiJj
tPiY6tj7wzw+QXQyFFm4lmcFSflLMS0G7P/UIJxIneYkdOiburMTR4gjJWTEdo/+AGANlbxwKMlM
9jTBrEUspMEFNeyXSf9kKYajzH7/6xBu/UO2VHOlEk3QY76eBYeUsqS4cFo3VDpnE1Sj2frpIeUO
8L1mBX2U2jjtDv0zf5RYIno1tgm+GNqB+5LKcO6q8wifbFqRztmyoSTXZu8Wp9JisK0XIWeZsGFP
xMTP7ZXZ+q4RLvVflU6WGYhNLu66+JV+0IuOPohPhnIikUGNohSajNTEagkpDpsbugAJruJul/xp
580xv/Ks95YYX4e4HiCzcxuFvQujqOI71VZeAGma2uGkZ+ca3M8Syq+qOaf8EAPOtaVU8306OcaU
F0kzhBFDFcyeuknstoCyIvU9SzMpLjGpsD/MFBXQNVw9huDPkW+qVJQXQrkkPeTBjvoWS3R1cbG5
sUodPfIu6c64NLfEw3kGZx86Cj1iCigCpu/fFX0+XcXLQfRjBSqrIkUwy6S2njp102ETb5AIPfOY
Abluip5orHXSyDXMZ+XKzyQiwz7Uk54hJU8uSO3+jICC2gW0od46ItAGErYubnwQcxKIZ5K7xYHy
SvsV72zrCTfodafPW/hxGGIl5pG37HlbKBVYlKeR0krlVhTBDK7LmVQ8zv1Wgi7BiPzEtPSUgb32
S2yKIi2ctyDEmXm0LaARaRK5kCvhReS9duyOV3D9yYBauKb8dFrqQtx7Urrk/o/NN5E7cJeurQaj
EYsK7Emch9RgsuPsV5VAWp8E997xg/Utn0VpENouPeas7AB1MCcRt2JqETUPTtJU/R5rrACxgI6i
wWk+VwXNB2N2PxXNIHWlf539eyndwBDoE8bAavwKSiRZN8QwiZdwuRbDhUFEV8kCQioSlV9p2CUV
mfOxcEmlYI6qpYtQcsn6rhcxMkz7gBNxh8PvF8VvwwMMwM6GHpHqQ5FgRanbI3jpGm/fpDlc0l43
hPAOKjZcH6eG65IOyUEZSrp+tUn2OQHxvnhLoQgTRs0wwIwsB3FVMVGeONoR85caOPje3OEEmym4
lCtoOYC9g8ar/amZ6GyKYf6YR8BZrXUxuV4Zm2iARjrnr1YgTnwsR4uMrAKZqSN5w8n21yX0RYSP
C6q7cKkfHQceKHOdTKduu2rY6aMfRBX3WqmVkVBlRW2bp2sV2N5n5ViQbH6tlflxi/BrokjooBr6
uS4Mu2XlMC3Od2Z08ogP9OXKE/r3BwAH160rXXgSRmZHFfDYC63gl2W2urkTcWQD6MkCiPzXSljm
QJfv334BDnlKrnly0WR97waBPnMdA9cMqHcn+MiEBFYgQJvYb63FEXtc22B0qP6OaqOFSgZj2S3p
smXvC6xH7f7T5zZxh3Nko/41lmHFSyDVPbjdAR5CM/Gjm5OzghFgtUqVhDukjRRuzKTLj4Zm1otR
OiR64MJoqHS48TrtBCHV+k5qEq8Mr8VYC9mAkObp5IET8/QpweRnRmu8fLfm4e3EafDEXhl3iriI
+pIOBg59o5CMcWJwYBGe6d/V1rM3413N3oLmpb19qrg2StpbtDcPxS5Irh3+r/OIUFWBjzDT2GKv
Sx1wBe9IUXN8TJaWv/e1QAYFIBTLvA0iKWTwWcDCGVmchMwzxZdEgZ1pjNqRjp2QWKF+HjaHbp1f
TA7zblTG3bTbmv+dXaJIgQgbBAdG9oFeLAIJsynj0iKt9qSDKvN16t0efp+t7UKQlh9dIon9BEWc
/S8qHn719qZ0Q8UHTf9bobgNydakDfXf82655L8wxXgDKJY3NJ2pPQ+nieiGz1XeL4kdAHTNc9zv
QsQwFTWgEFhUVa6bJ8cnnKoMROtSelLPuA3pcLMvdxrECl4mjQZ/I3GgCkjupTfkP3HK/bP23VPl
RxfTfPPAW5ofOJaYH04IgKdlusMZLohdg4/fbbBrnUwI6jOZGvubh7TZCwpvv9k9+EbztVgPXig3
b+N7iaUWFg2Kr3rkcDZJDhV4Vo/saPtjPnEoKLbdNCdKyGtCOLfb1Y1kAznSYZ2B/h7RXvLf3lMn
6dWhuMWXkmbhOnBwPvO8RH0ZIb2SunwBEs5D/+5kHI2uzW6gZvjmn0VnCkZJTq1k4wwqrZ3D+eYq
pGKs/wzvjuNmRfH0PHus6tdblPwEnZ0/NemO1mnFwFkHgBqdhZIwEHsm9NtjAicjMW5fpkN+imyH
xDfEK8bGgk1DwTeH5EaSsRGBeUxBJAucwEPi5phwIHH8/nsCnKzFZVWFfdSuoYvQpRaU5Jd/pc3D
ToII/xo4rQQzhkuCr41RZgERTAFifFOKnTz82sFqUmsu0F0vE0R8pyZqg5UYWYIub/msYEKQ7nhp
XeB1kYWwQIznGvaYNf6d88dbWJ778crkI/aul4HhGrPUfX6QwaPvyHXpOZwZ4DEoEWl+MPvTdk8x
PjkE35CUwzru43SeC7ckcV7HaeZ7tsIh68jLoKhgo5P6ZCCcv2wclD8LYS0oJYsxIDvZuJ4qotbF
WMSrEBkBEV5lSW9DAnz6TuCU5crLGGIqlBaI1oQxM29R2/1hYOKDE1YryAVvmT3wtumVYK5naPF0
MooTrZv0Cz7lsYNnWX24vlMGTi4zZ/ZecPdYenUaK8ly45jwzBZaOQQdC8kMysO1EH4uEg+UHp6Y
AEXV7rTdGo8PKpJbD/eFVZ2PKJp0haV8H4KkiBGvEk0CSVSajASzXRc6ZYjzyx5UwE3PwDu1O/tf
pFW/0Pp2tj3nA+LGdrH08pLV4I8kindecspPR4F2TgHNSRUqv5ttQ9tdH3UggmYRkjqFxGyhWdLp
NjEpTiSA2DsaeFi/u6kN3hI8XOjj3uh5yJ/AyC8U/cu9WpYPgrlFUqeT5Es7vPZlnqpQ1/dNxlhS
bOSRkzlWW07zz0H6M4dhJ7yCHZ6DvlUUqPJ72FgG5+t24wldcNm78isC98AmbI6CrRteXMwEew9E
yArbA7XIH3A62lCT+V0TXyKZ4VGnzEbxg707579+M8RBbSgwunEKV7XA1LuW29Yvgh+e+nHOEPk2
r0M1S5fsHZLM9zGyFE9UyFqXz3HAXKj4sfqcJwSqmxXakW318IJ75Y4w2G2sTWiHXPVDP+84yu8S
K7jnbPruYLDZIFqsEgwZsdOz88yQPU7aDgTK6srV22DVJlrx/NcOA6s/ZDW9cGpthGrn6PEiceyx
AxZq3d1U1Fg1RCykffDTIPgv3Uj+1hAwp0TyFQpWHoZSOTQQT2vaBCVN1N5SlO/Y9hCv0jdSa5Vc
Gx9/XaKB0FvrJCM2dwaq5xJW9zubMt1cgTiQxIB8AYC/DoKbYy0neVxrhxUBMZXFbbKwu/kom0G+
T47KwEcxPZpUcMsaDMtaBe33u/Q5Ju+ysXGBWoz0NifHrGvBfXhhElJvNp9WOQkDKbA7+/ywJM38
BeKVfDuUTq4MwiXtEnbhFFf8QaTw0wcaTyGqZS7JqtMhGq3e+4nkK3xHNTOw8KBhMCXmRVtKRa4j
StgdyQ5qQ7MTbQb7qumKxwdOshOAsxKvmsG2kkWqNZafRvxDYXVONH0+tqQiOEbYToqeH+/858bw
N9lti5nmPUrF+DA9vD5MJhNa0wAqfv64wwaFu1TASyFEhd2kGQhKYwUBHroPheS4l1Xm1btqNsMA
1JhecwDSO6NEc2guN+56pJa3u7YMb5239J0UFOCv2JEB1Pz5EHYH6bT714caGNbMxQ1NNopkGYpG
ItoKvavjuav6uGnwcPML5i5SyuljjzuyxEQgm0ACY1rnntdjhh1atLdm7MIWTOJolX5G7xA1gDrH
lIotpbOdeYVfUuDbkW489lu/6+Jn4L1+HnCrAH9n2II5qy/tRKYqh5GuujxmT3tr9tT+bBQq4qeb
qb7x/KnF+7Lc9IZ1aCi6B2IpaJxwnZHIx5MyIbiIcuInlcvzNfx7xBZnBubzxmXubQU2InE2GI/M
58fIbJCdKCNTmvenDq1rLxsOGlSb9vh9xJrtMAqS6YeAuykti4FfDEH+wxfSwURmIW8OEFKmW50F
LvLDvGJcqt0z7qZFG5pR9aJ8/EOFnPwC2z0+UkrzB0UcCFohuXOLTRetG+TBKPqiJ+x3Fb8N6gxQ
q1lixAg7I5Uof9gZC5+iRKdVOkorn/ln6kFAvA40gyyW5rypa4phYBjulNB/1YZx4wtUar3XyisU
qkl2tXIbMf91Oz+kk2SssK844c8OBkFEj/AnbYZ1SI9QXTpX5i50I38WSZQ1OqbExPTgw8E8akLV
jac5HHzAYXpYtelKI02sPazSVQInqsbupMG0rwWP+O6Jno3r4ILC0nXINpNKZZML0wNtE/JJqq2g
ykrvfG6HE6rmNp11C3eKdAU3USkT8TdOKRWui2E23JN1f3fsbq+zjwa3CcXaZi38WT79E17oP9l5
DowAlwaZFBB23TkyEGX77G8qaK7GzRCV+o26HL+JLTwxQFHuWf/xgvPJylK+3cMWTpKTKwxJ6R8o
AVd+MPFFtM7fdc+AsGt7ZA1c2MDXEzlPtsChlOvG3v3uY7vND2PQ9LBtysEE73TcT19AF9DtWGE4
UGV+PYEprkKXxFJRHqSjCP//QgSe+K6G36co0cmLt5q6bmvcKBDsJDvYvzwlE9SMVEACcVKf92LZ
YPmD8fDvjNHr9zNCaPJzlqQ9n/4JQXkqt8V5e5SoMacBd2QU6n8msWOcebXopDckBhkqtZsV3HVI
5x4Dhkid9guPlTlXeRI2XYo7DAoCd/k7sU8fs3Ias0LqUj8XwbeZmlIPnGijnwmhr04bNHUQFyYs
NUoFc26EFJZk+dJbjaLa4dH7SRKJHIzpZao0xh99LovA+sp/ZyHgt0iwBU9qGJrJCaH9CfnEdIKA
EwpPgW9CcJCD3NcM0hhaPWVOso/H7ZnkENkuQuGFDcxcX17P7aBJZpr3T0aZf8B87j2RQwm6F4mJ
Vd57Y/fK1fqX3ZEfJ+T1mRb34T2NBb+1khcxqsONCPql5CTHIubM+qbTF7QsYEDI05CksWh6L3ga
Hevh3VLjBQFRX39gCzQlFOn+WMMtREQsY1MIGkuHqwP3VWLhM/GHqv6bHs+b353ZEra2VK05znZw
OU/+cGOfUwKi5Bh8RJ/v4bqBpKUdvOHg7UdYY1wTwHXZkAwbhbWaS75/CE/9Gs5r11f3AEtxF+/H
JJStSPbPkMbD5iLF/RMhPlVcogthS6p2XRjE1H6zPgJ3VrJOt0FzVMqyrcJ3sv4Tm9yNUQgjJGwU
rKcYRNNtIZ8oUBVHQ/yuEN1nGpzqIM8FL/puVZLJj2BwGvZI+Ng0GACMnn9NYnUM7gNSaaWge+ND
xI+kaEZuEBR1klLR+HdZx0CkHcJlvGwnFCFY3OPlIvK+EiecWZ4Sr2An0/GTINQgjdQByIpPexyG
jf4qaUNuY9TpozhwmPYxvXb52xzvYTTasJoKf+YQLY1zA8VUgsJVN2GMJf7kDxMdz44kVERRUCVM
tPE/4iip8/500VpzMqdCh33IweoRByUssVQdgfSVXdqv+DT7mkyY6EyeGxeFGjgSb52vUgekHM7i
OMhSZsqlsHZAkg0UmcslgONLMKkYsIRTLL3kWoVpmbFvQF/gve/ndwPtdf3s01D7w5iEPATs8Iuk
zxBxtQzSrawDabuTSKOKUjj6F24T3EfdOK2aDJoYktcrQ/sludR5F3erYPHIbeDqPkZGOUPywTMP
wyksC0pdRn61SqSo4muHPHkhFsGUXcSHuiVi0arM0NZr8Laxmj9xV/ZxiyFaOmJNnWzttGslhJtS
wwQBdtCKSlChbF2+z8ISo24gs6YkDVucudZaa3uM4p515VOqlLXHPazSzNTkS+vlAny2v0moKmxb
lThaKF0fsqgPdn0ge3gofNya7/AC9TtrvUKAyQJWqugF6QBFoLbGE9Z40KzoEmkOSqpgfoHtcRgu
P79ifVwSQqJq6Ih1ao5sGITKzXXdBS9gbE92OfItfPssMip2m5SU1fjK3tiHBMMuHI5IhAzKu2MN
BI/phOs17dhT24Ns26zChtSDlgeZw2hyGnRmi0pif8EYE8fUo7KPssU3ONa1mDKcyNK68ODP7jzT
/62VrTwXbhaCJwDHElp3yH2jmXVDQmnWu3Hm4uqiUFZE/aeiAoTmkK6lItruUPMplVNONG1L0ubJ
dtGmWDCtbCQymXYDhxJrGlfmYGiCU/QIU8dffg7r6k0rKIpqOxEkN6tei11b1GMNMnAUr54PPka8
JFpqbBjqAvh68qW3/CvbKWpmkkn+fmkGKM0vOYi1dE3okHfDL+Q2O+nh64WaTCr4jcxRx50J/TwF
44LH1MmmdxNX6k7SHa2GvGyzcoV4aHAAD6HMzk44hefTqyQmcp5b6/V5OOzdArHU/MalFQIK2MXn
GvUErIDP3MyNFt4TcY+hg+w7izJ4tx5bkYwVUhc7C2wxrTXcQxnfZ1QNwbY7BORqVMg1GCLTCHFb
rs5aNtIb6y9tTKYUvTVXVba67UHTG5pTe8EpXFgDvqogvyz7Gbjpdp9iDmlVgMQueiiBQ6ZkyIhj
nFVKiiswFNEE+uxWpR8kWxDV0FE53/Hx7pnuMrcldedWAeYKnWh8p5lnxWZrHVqieLLwhvE1h+/1
AeVfLeVFuTfhZ9NfNxcWjmjrMVvXGCupWCteQRFKqR3YqYbhTCZLyTB6bz1lzNuBYlXsSkFuByC3
wANfKeR4hVEEkqHVxhUZAojolQ2tio71gemjqQj0u7EeuDXyHNfSJjZHmPXDJdMIcCvR4lSphtnP
DPqZaGJq+a+yeLZfNcgBExkm3JoNLSTsjtxBq6XgyH/mdOZ9n1cR5iVItPnblt+DN8CzhdZIikwU
PXVa67wDxAM0iSvgYnkfZddHiDtO5z3lgh/fxmTOdWAjtdyGVk7h9gyxZpy91Bt4jCvPOdWASbZN
lwJKeHBlTahxec1euKwYWnb3WBkSUsTZq/vtWyKf2XgdtNKEIfp2HRHUU/wH3mlUmUNfCBt9TjGs
jymhb82Axn4Pv4VV6nFrCOcGlyz/1LFpiFMTzaUpXS75Pi1egLGdwwtHwJuU6LQglxVnCTFSwnIf
l775qNrOknFEOTVSB7iI33qdyfkBYrWIZyZdLP3fHM5ylXC4qaOIy5Kq6uXUZIIQUtdlzQrMIsTX
zVIeWVJZDtlrQhS5O9Ubot5vOGaMEpnf+e7lsoaEImqFGdZHN0+1M2U70pas5Dx8Di9uRUb+pRnO
onC+AJhuiRHSpimfsu/2YbBiahPRQU8TIzYEoWrZ27Yix6aIRchpqsV1Xe/sCBTDySe1fGRumLkC
bnIZ4jjWKJguBt/BReXlsZY3ZlfqTnHNRrJ0Z7gU23jXN6N5rGL8EZ+iZ/4NxxdCLUBBzNoeK3r1
PjMf8vU3AoenY37IZ+c6X0FN/NcGhDs0x8d7GJDvJocAsXVSMxK38RGxecQKD6lR05SNIFfpcR12
aGpbHNxvnNuRNhGJFKnHTmg8wI0VsG/QnYZKf/2EltxsWmM82CEslrl49/SfIuIvCw64qjzq69s5
2P8y8sC9+tDvpKcpccyLjWrLTU/ynwq2veHPDl4L0hDGEkKsUpwOC/P4kB/fiNdxbBo3Yk4LPWBc
ThyBhLu1JeGzIbVSZsV2q4ULifAQo1rMQNZ8Yo816ucVxbtZQ6P8P6yWk884p0VnTwNWZfB0KDBD
38vmc8JQ8e/0R6rkhvqurqZd3GJsYLx50bgZHAL5bPtX2jxACfyWa7FMccnXH86xCYzNuaWpJi2T
h9NwVA/po5epFuh0LE5W+IdCcP+jyKgqW19wlhRx5hUoBBVPjymqRGEMuB333KsQ1QVJNIntSeS9
0sPWTBzIdjLRg/AwlQbmeMo8Na+uQXg+JoBvUpzJnRNuKxN11TG9zhHAcLhvTVqZ8/tWGMJqCvqO
YzYxAKDYGH0DN3bu7xz3ASp8NeKn8yFoyhh86t/76Jv37LKGaDLdrPyuUMlKPiWhzkiLt6r7TXd6
GGwIqGWRVBXj40xcFPP37rktxz5SHzRGk4TkHDISUeCqacjmun2A+EUZO+u0u/edhKqMzFu2GYH/
pGkSksGhyGmBuKR/UZYLCzVWrSSxLKUUyTYZfzv9hG3j1lvnLiSR+rWbDND3zqLGgmoCxBy4iDev
pt1uyzPr9q4skMzuX/POi/IaVTOMf9ourGtQ+4StjrA65W+fjfVQizu7nKUTXMBY8WHlP39kRkZu
ZGC7uRD77QE3EaOCx65hTGX2Je7BjjVIeYpiZwqZi5UbgzJ6URMCJy1pUpTgIbGXIOLET6mVTBeY
o8yiKtOESRe5xqmdHHRcUDfRDr+TOOkD/1dDFFBtDrpPpXLWsxjA16gA6po0rr1czY27YisBw/S+
CcEk1iX0iyM3cWY66HrokbkB5jv6sadYoJA0Ab+Kv0nkUNxZyfEmXhuysFaPvE6W6Y+wmxpAydMY
w8Y7WxLhFNBSIveG/ZvCt8JsoCq3cgJfxuUgAukS5UNebY94jmFpa/n5HrhiQotpygWtA1H0PS7y
uWV+UInYzTZCM+ud7cZ9M7UGDRZWaBtiYT+ElzL9I71x6r9fPUezPqPGAP1FAwS0CjxtkiecX78P
0SEJOryCkR+RtNryt9gbtVx0byKuweb79DLIBV8vdf9DsPI4kPTA1FFvYniAc8pyEVTS6fzoiXg3
/0ODOXJlAmeX1rjSWvsCLON3j/7yau44Ax9XajBrRHGsVo4eV3IfUQmfpQjCsjJREucsCYiP9zgz
1biAsKdkL2XA5hlffIlOrvNH77Dhs4LO5BUE9kKB7Unz7BvPwADkanX4FDBJciED6qyqjOEHHduH
UmNtngbwKayIfQSX4+S8jmm0JSVEYt9W6fjH+xZydp1qCJwFzVP7BamucgqH6WyivvItHXWqltiR
gDEC6YSd2ii3K63uQIPE0Gw2C7SQDh+luVlrBThXEzQ/6jfJvosewV6vEtw6rhALqKYOcWDa78Mg
JTw/JY6AuD7AQyBJJhzrNU96Zbo7Pd+nsiru/ixH2L31lRSZWJcJVx8iux4eHFcLjMt43hA8gJo9
w6f0BTuzAZze6QC0cdX8OBJO3XFRH6oVfSog83eM4Hc1hqHuy01tl0OOq4ipbbyR844nW7t32rjB
WfD5DZ9+1HzWymDpYgrtBE0aquh6oBNKos63ljmWVQ58z/DYALKs6FDPsG5haeAogG7gE0NvGxuH
UJTBdmqQ5vfg5ePOp4neYebD2yx+GrTcbhsa/Pg1H/AhsibvTyc2zVBRKyCV3l62fswQFadL+Jlf
MSV/RSDQVm2261Wv23Z824vSM0xaq6b86I0UdB2/QhZlbs0cQLbHHZcw0+0nIggu+y2GnRVx4boW
LEZ+GFCC2yS6/Oe8dcOnjC9bPct0IGGaSIk/2WneJ8B52qlWE5Ak0c4WbJ1S7xYy88PhJQVCCliZ
xjS1T1nfM9JVWpnQ3rXmn9K77IxHoNAkcl4KIDDhp+VDuyslEgBTCLcBvrFnVn+xvhorgWmxK7lm
ORWuUcJUaYBnr4oBPGWmpO1Vr2HH6/1JFe1NU+bpfAyHPIKmDMd6sW9giVYJ7v4ATVN/R2ZtcxAw
DUA5Y1F6F/uQLIgQiVif7kEZRW/eFB9IoLJ/cV08jbqNamlb1L6tv+h0L59fhqmE4Ruu7yJ0+3pM
6ggReYbxeodxaAT6ClG5TU6WcqZLQF5vAtMJpMfMXUrNmI4ZNM9ZnOywYUL3RWq1p462gp1LFSJu
usXcvrsAbyYp03tI3PiVZJfpZx2WhmNpBWpT8C3n/ZkH+1T2rcz/YW39imPL3Sg81v+lv4xEKFTc
Rqc1cvzcZGXQalpxs6zVTd7jdjXOR4xD154JYSqauSDNCTximjfvKocwgrJYQUG8DcMjONeB/JYI
DVkI8xI4BeIDUL7+ODFAqVWGcqzC+CccdirSxZIVEzP7RvlAcJV6mcKRMNsn6NhB4tWk4VAnIONJ
hJDMNlDAHN6KjBE4mYRB6c/mkqO8M7V1F+26vxGU2kUNQaefADnYTlPbI4hnhHIwuB3AH5qMlIUI
lLH3C+732Yt2i4EkZ3W4RRhWsEUTKtz2aeoHYON+TbqkDX/PvjOuk0LlHzY7an9wdkA7zhu+Hoz/
WzQh+5GXFWQZhrE3iX7qSWXsQgOF0u6hETOSU/q3F+LRjsSfHCdpxdnYyCFODxPXBayHnF/h8qYD
twg6cqGJyEX2lfvUrL4Blr30xRAmOLZ5ftkhJPpAGZOq8Tq9KoFGlobHavBml8CH3HIaIclMqGru
JZVby3wQ1KhfJPQHzj2ygy3FYFGhLionj+IFrQKa31Fz+ERMK2JjRUWitAER0u3x6NvJgJAKppkU
f3x2O/KN8f2t5TDn7A7BKgTktJ89etJERl6zT6tahTjLU72Gkw8RVDixPVLQ0tJqKWA0+AdPlylv
o8lhemsQ6DjJt7Y6OHmmJMGVtEA8gbEhaWlnkjOnZRMpHN7q5nffUsI+CKag0Ejpq3Hzhdk9sshl
JttOdMP4oLHp6lbmLSWzVNKk1qwXE9F4tyq9jt5J7aQxEWkrdcSIm+ac7H3YX1zK37Ay2mWU3WA7
CIOBv8PdMgpAPY2gHJ4lgO3ocrMe/3D2diXWHRwExHmZYem/nJtRkOttNwRPSj5x7hn4quR0uGiR
L4BO1A4I478FJtiMO3RnqiC794BdDs+05SBG1sIZH8eSgLRcW2M0IDs4VZDqVjAMXG+qemk2Vb+0
NWEPib/BAh58qXyJoY44ezuaDHqdmOHX8qmYveT8zz6xQgr5HvXlFL33OMuuChJg7ZMjL8slukSS
lfK/kjrCexEI5NPeO8U8/bYRWpZUpaPKx7uvbGyC0PlKi8TKDpFfHRXVBGVGuhpNvi76h6opG9Zt
W/SraOiouzllA5FEDMzn2qS+/8U34wNoI/nC9jcuiUdvvutseulR8aZjXpLSaE5y+M01+H/OiWlW
cDIAI6HAwZ2NZbeWEP8Yy6XgZwYoxZvCbpReQBOaxvRF1Bai4h18USdR5RM1HjjEwn752BshhCrM
krhbiRMC6LdYvDEZTbPOicjVyC+ikwHycunUDX6zBYSa6WPWwzsFM9MfHC+2SuLc023TuaDcUCiL
vun3e58/snHasGeuEi3ZVM9OUchVuBJYLMLQe9rU1M+8gKRGA/prI0DUtUAzD42b3ORGLeEWQrMj
RmiodMsA2tDPFgdCrEEEFehul9bewZv57HaQMuJkHS98Nm6wshPVTXFQse7fAx1aAQGPSAkWc3FA
qEfkhnOG7tiYvnH/LOvlAV+S+p5s+BSEXNEEVDd/4mP7TUzY2WBOsOjLdXWr1w6zl2skILEsiYUV
m6UBSvtraxWk7FRSFLd6lVVyG8KriwPYoQJBVkv4vVdRVCSUuJ0daw4oS5LrzHUOTygcsaawhTxb
wViOkWZ/taJJtYtlJN6fw0f/0Hwowb4fpRD/MT7vcPanlQ4wPKYr449qgdHEPzT8L7oE4xqIehJv
5l2Wl4YOHTIvmfL8DFnJrvqcZ49JL/b/8BKDPoSicSKfxNVqPEex5rS7mlkZruyifQRrsZmlHFXP
r5V/JHOag+qM3IjZN0twVv9Z782d84lS4f8kCHoqKoC/KzqQnWE48CXFheazMTCiEDjedIhU6/Cj
g7fNdCGGmJub780JK60tTjnGtnu/KvwkqO5VnpzwwKfofoZ7SW27HDIOq1sbiIkLniteZ1nPHDEB
rhsisO3vqncLYZ5h/F2rB6NzgmAcl//7zczHbIVHsCvb2bXaz++OWYiOom9EulB+FOVXn0SunSIo
5dqkf0gdAelfUzWmSZpE+sJZ3a/Gb2r+QxUJQqPWaXjQ4kBPmc+AskCNwgC73A/2diZwP/DRPb4q
85cBsgLPscoi6+TjawlLZIR9OnmM8t4szHC4/X17VQNvY13EJLwEYPv/wPEtRkRlSp3ftzIEXK3D
hcxI+LwNUlFC7ne2lWjl6O255S+mSVJi9OYvr8Z52hnFpnm5x5ZJbzKHJOvInSe+NnP3GjpmINCt
B31KaHzKFiWdaEVy6IlWbAUVyX0ouTIAVkHtPmEYf+RIZFKLdFcv4k9bL8KRO/HVKT25/uslGv6I
iUTi8x51X8Yn+59I+YTnmbNgxUOaE7M5ShxKDEINx/jXsHUiM6vAnHHqn5bBxugDnsp/j6KtXPCV
muQyAF9+aAz5BiMHyRjLYGJiqTFTMQzh68SKNIUAL7c7T0eSd3xCJ+BpeNaJFhF/3I+udg+EcYD+
ZX6HVNlkr5DAIcrhWTT3W8dYgbnj3zYKL71MIilKaPadfRpn/L/swdMt+tg2FPBdQnf6JMuJOCun
33MyOOX1HfuaxLsvELkYaMJw3uX+r5W+4pn9JMvIXsLHm0JJvko4GVbACKEQ2QnKGb3tWvUYTlOA
3ztLzXcUiOhAsO0E72b+C9e5hfxKdNX8Hn1bVwCCvCc2KKfqjjKACR7bl+2jGvRvQ6bOK9PMzFQh
HfTCJuRodcePiFC7kmd2SYGR7tOYwi9au2AlsoXiFJxBhNKtNTFpPG6WazZ8AfD5zjbcES4hrwSW
7chuXL5zwEyjMX652lp6uUhr0OrAsXqxjknU46XmzyQJYlf9UQjHm+rRt1+TH45cYn9XXdjbunVE
8RHGTJptf8gfwBJ985+eDCBwhbtNfdOaz4/ngLATT+iIqyi2sckxqW5LkJyVwvKFj8ZluHI8vJYA
MTn3pqHLtqEiaLdTATmATTyaQwaw1KZRBvDU0reG3KZ2Tme4yZCL8E5OKaAWStr1cPgvLeHjmIze
yq+aKj8IlMVztA1zKzd/1ZGI/6O8xS5wo+wyKF/tpp0eFFyEMo0o05+csd1bkpOwIqH8uQrtJwuV
3zFEyLeTnr6Cci0yujba+QHkc5WZKHdXznWAL6ymMYYKBBAOx9kWB9SHlcX8OvbUnnZtwfyThcGH
KW0YngSh4zc9g2TaXgs+w1wSwMV2JQZYMC/7CdSbCfUGdZEYFtZRcTSrKpOYNR8mgQnTU1P/2ceA
sx0VmlCJQ7bD4QPchqYsTbEoZjuQIUnjMQbAewMx6OlFlToyfztHBw2wtvX2ZxY8YgiNrnAHOX8B
R7eHK74YDR5qRllMg0n9pRH/QNz4uRO9dpeQrBNm791sAkUfPXvuO24/DdMT//KEcEZ9oQlBiaI5
vloJ7n7fvONxd8cpR/rSlF2nfxMmM3RUe12TZwE9qU+6kzoV+Iti5tffc98xzsORBP3hRXIajnws
0m8TrruwwrtvftKoAHhz/ON7q/UYNYF1lyAqMkLv31qnbDhdCuzuiOTyk7IOwH8srRyIMpLNVqqi
SwwUJOxeDzqzP3QFGH3CHmB0l7cy01xu/9kBQWf2RVLfwDcibt8h2Y7C3Dno2dwmKuRS8rpNsmsg
MDzGs4J9aSr3DAQVqSBL7gOxE7XMFwjaTgznBYmuuQZkKX1i24RfoiAR38ON0D2Q2d/qsa8Zc72B
t1TnJ+phyPjqmBkiTArWwmPTho1NNfJAAyr2hiUU18X6qhxGxP9GQklA08Cmxdge9mCb5R8noNOX
HZvlrJgVkBa0ShgGM1LOrkO2y+z2CPBAsH7eXtzO3o+UFvGGzAsMndND5w9swhZBL097EklrL1Lv
o8E8cdgiIbeZUfpWGtW66AgFRNmh9JZaJBxITniMJJZab7W+DaJ4Viiv63FA+EUoV/RHIo90TcTY
W9/iRPLwpqIpY333dlNwgHBRtgYL41Z0tq1RQNtdfI67s5OuFCDe04y5VE15rkgr7DpbWtdwgBLE
ljAMiXDw6jGMSpPH6HCEZxv+N3FCIZoX4S/KkQpDU39rKffXYtz39OfmawdRevKuHwQbwywNaQ0j
EsBYzX9Rr6EVOK0fd93TteOE140LXWu7maM3guNa7kkWxlKQMXh/CLrViR/GLdsVBs5Vii+fVmOy
PgIDMPf7rRRvTUwR6UJX+qatjz0zyOVwp/iYTphDxYWz1t/jz3rJQKu4K3Boz1b65xK/y6/auGNw
sRmY7m3L9w3PemUQsoy/kzeyHfIZuaCi+CnEkrqIwDPF8V1Ar3EL70IVZW2+rbmoX65WmzTiGBV7
995tnylYNKmtGP88PMdLRIihpECLqowLnLQrKR/Hi/8yz39GkeFm4YTR6Af9r5KIawhn1W08mRrU
5RhQX87q0rkccooVzXP9IsVRE+isku/AYfozcRPmeHJV5TYIZKhSGaGRKO75vVAYbFaRLLskBC+O
6iKejlvj1AwRyCmHfaiw+PiQO8h8O91s6HZ6WupCHjzDd3mCf2jmwC7coxU5/2g9418ILGRYMsCO
IePCF9zbp6dkXgWDAr5GMeJBqurwIjj6R3m8LN5sjT3rriCRbXcpXPl2rVNQkwKDP5qqqY3Lg3O8
GsQAQuDM4ccnnda0MuCeAro+fLLk6nAJqR/nOExxpZP6VZ6x60Np9kKOuo7FNGPLuVmIgsgt1jgq
qZMOqc1Q5SDvaA6JI0KmiYedpLgWFUhIz0kSv+mPJuTTMVXxAM48ZT+k4yvn3QmBihjwS0h4dVlJ
zJOBhg0i+9ojdgcsL242z1laqYc9jTpSMBbjCPsPiwsB1Tqy8ab0sY5P9onMLbkClYbKl8RiEPeP
RVDD4Q6HzYB4IuKgcfHskY606R68nmlhp6z2F0Qc+Qs160CF8rLnCWOCUDV1DmNKagYfogcEEq1h
OxXd6tW0UY4MdgIgf8pC0YDfpFXuA7fp5J504omdT/ZQh7WfGSHmXWDcp991xTAXSxuiAMMSpCD1
r1KZtIAaj5UiFOozXjy3VOhWV7sj5VVpkhjCbtQfJKIfMmvtXy1u8wQPakGKfQoMvM1HRTPO2sYm
QPRkdL0xoGdNSJ/EvPV4L6YsjMqFYQknWPqdxcEycC+44UDn7/TWD87U9KIw2pJLM2ajq2CVVK09
4JFpedY1ZLmmkGFJb2lG70fuHm/sFIzoRASjEbaSBTkCBBw0/KI5KgrrRay8neb5B7/8K8+9GB2N
Eifa0OKnNfRuZRzJz1P4h5DuDk2jHdbjB2LmkhSW/pKHfEn3DXex8/tg7CgNdfjtwKiAMA3HBKR0
ErKIMmsWjz2I3daF9JUy0oE/o5jdPXNoOJxSnyxnwDZPKgDkxrfCi2/EVicdXdzBRlstDBjzaakW
/1BFhCKnAKWRio5CtYO+lJ0nKpID+0TaLCbRwUnPMlyXC+5Y/ShKUIaAhs6+oT97l3eDRfzwx2NR
z3J5l/J3C0k8b12H3FzQe4jvtgOThOM58NLU/in9FpK6NDwzOwtPBKD5QF8jX9prAfIGJNfdbJpQ
xcov5Q3eIww8a+VO2fakykwXBQngom3ik7o1+spn0A22YA9ww1DGAkSzCSoKaG5C2h084Pah+kVO
SDke6Pmhqe3FQOYfjGt/z+jsfsW7/ecRTO6ngKtu2s6fD+K9pQqfFBWYLxw5nwQnme+ktKXDNj8M
+LZgFFm++GdLIspPOPA8V/V4LpQurQl6xFzhMUwU+beLCevT5OSH5jX4RyGvT/w4vZA5yttRoQ0G
9S9DEnN4wM3dGPRnWi0UlmzJa8f30wXeVFWUZ3ohfoXkNvH4OclFXaqCvBgjLpkMfcUER+weE2j5
bAJ4p2LQnAxdNA1eBCSXenYFlSjoZh/LTbf/a31uNBjpglmTZmXvb88Kpn37sPrkC3Erl/wd14qs
s1cPUEUeYO8gV2MYzkQ/dcn84OBFZsdY6iV+61gBOtbGik739QV0VA+MN9/48JXUcr8QKqCw/t9k
o4txy4fLrDUJyut42MaMrYp7mEY/PHAGRRO1QCtMatqVoPFMIVM9FmQNdJ0SGmrcL/5Jf7ZFjGcq
/bzWjO7Dxry8tNiG5mGlwkRn0reIpD0YzIHrGENjPpXPvxwT5ymr9LxCfyffbZ3yB2wsnlAq3ZwT
MUMe9xnOAIUYwV5gig6T4yKhImwKmTRgE7VjvgC42/szr0P8oAMTugQskRREWBFd0MJo31mRNbBV
Dkj9bPTfny2EUWgxNIBm6KuqJ8sZufK1KqN98w0f3EG/Y17ch9tT/dxADEVa+Sm/drF+Hcb04wRn
j3DfVzVH7xAGi6aIfQfvQuPfSnuA6XZoRKUDaMg522bw1w2f9yqjMWWKfwZR6NKNWRWjpnBm0adj
jnT+vA5iElcevDebAu0o8wqe9JulftupMdM+2TKIx82OqfO9vzg232778fkxiXi484n6rTDbnIPw
Dxrj6NF90wIwTSaE2k5IbvPpcv6/kxqy1wmTU180gR+ZmwKCENZXilxmDVx5s4jIUhYE/HKpPzor
uelfu+xW0ttRqu5psVyZYucJ6ecm19L08vhcICmpoPVtNq05aw2Kjh7wO0EWqmOBSJhq8hsBh2Mv
RqZWU2FQLULmzF6cT8HGZ9j/uov8Au6qknDcZ3yu5+zD4rs91MquwkcrNmHyNgN+6H1DBeroQ5P2
CD2Ydf6HTV0IImXWKVjhvOy7fU/OGAGVHZVHabi+/lwEMMrDvUhPEI/OBEHDkPLTz4BIPW+7ypfc
vtHnK0aTuBRTk//l/CbaLiYcXOCgF7NGv7okQ0V54mk6dQGuF333V2fIX9o23l8eLTvzHX31HXTh
dntf7eqe249kPUBn7unr1HWyaA8tvoUjmD/UBCgadcsZ13PM3vlzmkPzsSF+Z8vWI50n6QdCAuB2
8RWEnpj7C3QJcJfKM3CSpQCrCyWKgY9NqP6VpWuitheaSV+s87PlfbCSCGY2iEQFSzCCrxYVgAPG
zOD05IpMlTRz0VHrUnII1L4Gsxr1TN9AxyWJVxLnmhNkkdBEzcABegBuTX92RTrMJ+sUGYV4YE6e
i28Q6GT5vrBhB9iO4qe6BYdS/HNgjMeFn94wZX2/FPGCMtoaipL1yd8be48Wqbtu55WdYi3Tc9Qy
4JojC7oWaAeXrMJdJd2dQ11fLBZm/ZLlMHUysECAUCqAkEGkQ4N7TauFmx51c45Agdgv9ALo/ds8
V3Nt2bG+Nvps8pOAdFRYKo00NEPLiiPrR//UxBFtvnasjKtj4kF0jpne74He9bfaMGEeGudHZQU6
pY2n5idPyk3xW5kzw4SfwCd/N7r25Fyibsd9RtsjwRaHWGQ9xbnvpoC9WW1HNK2nVtUeGfQmCC6W
Q3Du0xVnsch+MbgCAiTxijU3yfv0EQzdQCF0k0DuHuz+d75cytlzBMDiTIfwJbmL+kfGgbOJCKeZ
c3/OiY7nQERKAU/IZT2fQPKkET0IkoYKIlvqX0upgUfgdaITJXbFnqFCOwToMBIl7X0CyX8GaH/Z
8TrOQqwwrsGIYaVf6q2138OsxmEgpGmoAzqaQLlmCiHtuddeFU+6XlqYL89CV7XI5RBE7lUEMtLl
p9UNmdIerspNDpW19y4mR2PJP2s/gx6r5lV/h5zBMS2OwsmTW7JvjShnq4ywj0wg4cUMJdf3jU9S
To96Drt3nGMauANa5jVo3Tvgzh/IZF1+r/2uJCVOlkfkLfDuxW7uWCFKjLnRJ95NCIAHpicPerz8
SU7nHKtmjdd9WkxOFoAhmfTo3wHzHx2xD5xdahi/JMuIjzXFJw0Tea8PGqQ+lh06l0jyN/QFnoIm
+B5o/cdbW/6tKR9tI6Wl+BAgkDOHjp3292yHsJ6C9NQKtfV5BEciOc9LJXFe0moO09CzsLQSoFFA
Ug/2ygRhQLr6S4ySup/7NRsSzFRuvS08zfnoSnMgmQOfg9DO288ftEb45Cdyubf8vPdcL5AcY5X6
ATpH8pts2ZHuJGYhpBO+3YwDJmKwQSGN/9H7ZnrTDSyfD4SHNAA4mE3jL8o8SO6jcJpW7Kcbmy90
xeiYLWICchWbS5i5ybDlgsmZJLSIhm/arQXoL43PlF+cxR/5dAv0pcSqX5UUzUr73E9auS1/Qvk8
v+RgpXhBLb7iZK1WR6NhjJNrRKlSWBvcH5eunsryLyTWPdSFzyzWuEmuJcoFNspMcTnYfG78C6qm
5+s6GcGx6MPKS3Uz0ndV0XQk5Ov0ZZJOJGBBw31SvuFF6nvSwSaRm0whk27S/V3np2hhAAbdIqQG
NfcjeIUE8YH6eT+Easbf8V2f+99bLbhOEjr56omn9qXvHxOFUFbZ5TnSa7TvBYl2AWq7Fu5bP9/B
7prZoHBuAgweWeaZFP086eKFz6tf4Thfmqpw3v3hE9IlpIyJphEuyzLnPFUgVL+zCWe77kgyHgRJ
vC5geaI5HfhEN4fuMk3vF+1SrloVHhXbFbwZnq9WYQrcEfEg8WVuL5HAhQTaNJ0xbI783dhmp7Ac
CXKZ6SpxJN81lCbiOdr4fOnlau7YeXK3Ll4gRGIUvtU3EfYKbGH9qeUw8IrJ8mCTAxhdcaNXqDoC
uQ5ihBEavj/Kx2/LjTSG9wd1BzEfWEvw1/V71VqoMBluwukHE5z4sr9PzngNDwcxBlIdzmya45R7
Y8aHyZS9RN39KDYbtD2zmxyOioFhajNPKxurwiwDYSy9gXM5KHlHfN63k4KdnHuXv8kjPnbLIzvT
yrsY6ShNZzd63SNwMfKRuHY63TRwyKxYwZbURcF/+f9m6Af3oEvHl62T6CaBmlDsatFqdNDi8aIy
9ef3Fks5AE3CYQDx9+NxGXAeiscKck2bwJD4rT3VvJlbVvVvdkI4lNF7ylKJegHDCQu65SYqa0NZ
Wm+nHm9Hltlro/KZ/XnNwvOXRY29aeUGcdUEVwnludY3uklr2Gzm6vSu74aGLEKbrMk2dCgXb5i5
GN9+WFHYbDe9o0l6Y2jXFRUz8Y9KWrldmRAVPwoWCF1ai6w2t+CMypi7W7hPlWRXpSxOHwKninzt
gWUz8cvxzNgMi0X7ZA3Ii1gfgcncsmuzp++FR4IihQ5ZJz6KN6xjl/D6tRaL+wn9bT1rLxIYYL1a
sOTlC7axXhpBMna3S86OxaO0yndgS+LRv0WIOKVerTiVwvIK3lJ9U6sV+OXdsQgWV77ePdjtFkqZ
qjlmukdu6vO7ikBM+6KiA+WP/uJT/Ja+c2Gc6e9nPYOCVggEYOVLinoNCfZqaCFgKNPvKkC2I4Jw
HswLLZzq2P5OC4iD226/XgxGWj9GbRAYKbnETlm7f+KsteoQzM4Wg3VC06dZ7DGn4WekJNHMaiGt
5IXCdubby9by5LXQnVUJqreOmyrZyfu2ebMiGDzIkYNKRIxCsw6DGR8cEtQzW4fgpmsnorXdDC+x
YhGNsKZtiFee2LrAaKXKacB+aT/ytOY7MkNP/ppTFEcYbyyLiXB0xt51aa2ZR3tWE4BSxN9z5sOx
UMeSR8+UtB4SJ1JofIY7uXDdrUXWYGpKSsUaUev03+rznjgMzIN2hvl9H6uop5MQfKPipSPYq9Vb
rvL4MLq2Rcn9/IC1liO0UOKDIR4DgOs7n7vwg7IAFf2HiWjDimrrQG6bPW2sEJIXDWdycxATbqco
RI2jjBwxLoiUL9/sT1tiqpU+z7Uuxbt4WW6GNB9tdw+nk0yWDcB0oTlL6pfkd12rqQAXsunm0Lhu
M/CSLpLh0y1S1U9d8Ub8/6EsNntpSL+5FvImAPs1G95Fc+pf3h3+59b0fdHwowl8xyH/NxhHj7s0
jSEnEijiSGoD1HIrjuGb30UsWaAOFLHSaAngfcZnO9+lWVbX/I17Hi9O7pKBCTb3ZD6PGLcIH4Lh
PUZmGdaQ031tOmoopBOFfxlS1d8BdnNRBlnlAcLoQm6lHc6bB2aUYGsTSKxnOShJ1NENBRK88xBI
fcsc51leBGoJJ37x6Z9JQ8zW+q2l4gRqM8iXidJJZuGdNLqzGvzAQYLgOe3SpQdp6ARZcnWXNVYi
F/Nvp2noIZRapi3nbyLdzrnGEGcAcINIzaq9n5eNB8MuJVxPxKxONs9/o0bqUBu+axUwzFT0WBNP
CFejpRgaDhHLEYRauGpjOaHpgUZw0uIJSfhS3SLwuaNDaIaZx2rhTV9WZtLT6NVPFstjAKIsV+Lp
TaRZlEChu2Nz/YA9hpVxLSzXPAPmmFyotFbt+HI/5yPHQA0Bu+3hhMBcPLvAvkO/Y9qbZd4v5L4R
B2i3RBQsRSWUDOJU8LBSMVyFbO+bQYCJa1AZGVIGbU8Mo/zFfzGP22k4IEtWKJi6R/RdVVycURBF
jtoPau7r5+I94Xy797DavHsK54/UxLW1rObkt/fielpm/nd08xOvfo1/xBc3n8StJJf2qTUCIYMj
Pvz195OFmMmo5QHHKlgu8Fb2DM4ba0GmJ8QIDsXYjDGbI1WX4S+N5PQLCvdib6UuD+ONQ3i4okQr
givKopzUFB9MjLx8ckvMo0djmxDoEJeygvXwQ8QTy5kunuyXtuLK1p9FmCeZhQS5Pp9Gb1lTyfz8
XaLYfTunZ9NkyTXU6ZsmCdcg7HnMmmr8F2QxLwpnw26YIAdMZ/Q7AmzPPUt6czfceWcUa2FLW+PT
ijm/iYV7n0bEnQavugRvY8OoEz7fLSZWgDlLbX/lM4URkdZPo1LsThz/lKZ6A6iWhuS+P7ENxOl8
4nTgulxAu2zNYj2NVVcOUpVH4c+4aWHK1xbGfay0soNuBpcvuEMhetRDwNpqmK/T3bftVF8IjTO7
GHkbCmA2pEQE3IXSXik2aHKH2WhPO1i/jl1SXWGCSBL3JWHVjexGgGLwO5Ei0vaQyBVic/+F41f2
3GlJLTIzX8xqGr3oDxk4vKOldV5IdY6RkCOZvp5ayuV3Ul+D10sXq1l1uuIn5sDb5R3kshbNcmrb
sN4bNhBc8JcJC1+PnlsUkUFVpeds1smrURgzoTu6wbyS7t9BWFzrPJkeyYZIwZiOfUX0pW7qLEJU
l9lXf5jyJO1SrMyCzRIvo2huic7ziU97D56tbHjfdNERRsB1b6st8p/FV3Az/PkA7/qT0Hch/dUT
hIS+WRJUpyzbBo93bFg7KbYCCOXBVzLwcye6/Tc5oecCSiprubN0jwrddMF4F/Jms8wqcJTMZLNx
7jfDn7eSm10+/8p2mNMT7J9nc2dmbg1qznS6hpQxPB8R8RO26BCvnat+PUb8JQl1DgqSIJjJq1UA
G8ODtc6plrfc+YzOvdxfkPbQN+fTGx9vywYdxH2fpqwMEhW1cvLqQDXed9eS+NKs7FzC5XgKXDR3
8UItqK8NbrWpMXb9sE5afTNVodQLon78m2j46OHtRhuSk89FWIKuEB3jsw9QlL2qKg4CgVKQBRMo
OthtzjHJZwhZOtgtWzhopFArX9QQxnSXcno5gJbfu/VSjjenfyj8erpQdIDnmFfxoDmzL5gUVP9/
Ms4/p2s3/0e1lHOIjkVpzk6cBDNk+h9XOnNzJRAOvYXQUzAVeNKvxycHgFMQfeTdL8IQDkUDM00q
+0LjMrnzVXL3Q4RONC6o9GFmXQBLnH/IFqlCzWgRUF46VgOsm5T0aFwvhsayLUa5WlwnR8rWa07Z
ObVZ9s5jIx5xFdY9FgPFanQSS+U+oXZEO6VcuDBKaneM8ki4ZMFpOeAmklNyQp0Xn79R3BSmXpco
LIZAEh0CiS/KysBEVP3GD4pDn6RSW+1IhU5r+E2Fbi9/PkSlwHj5grpRp48NGX44Pv6DaGR+VMMj
l0swlmaA+sRfBdSnLP7Rlhk+50UIH2gJKCt9vIlKmxzNwUqYVkck7ve/Uben4+inwMt4rnOwC0+v
XRD5l98g8vRf4VOQNncEMF0nQJtyyJkR78gQ45FOqV3RVwFgUlWI+IduPLC4R8DYgnHgAL/hOlGt
9PCRX/lZ0uZpdHoUCcKU3NKL2YCwbxh+v2m7hhoOuZ8g0qwNVzGmUc962sa752zjd/5APMLJIbWe
5ESbsdU9VYp/EXzR4fSAs3qZwHFftx7Tz8U5Y2iIM3JVcy/tt/EZuMuORB8vAJcpYMJ8k2onj4aK
hOiQkKf8Dv/mmOIg8Mn9FksxXHLJ/azWB7UF0PwaZjgYSnIHrb+HUCcVvU2VC3b9x+ntRDbVN4s+
pi9tZU3snVaPmUhAkOKTBsBIKELkqbHLAQMumZahrFZDRpTDjrF0nXyI10NL2hglhC8O6spC/0Mf
zOjk4U1HRE+IAO0jGdIfpKrdyoRHmXOs3Ks0p3PSEHILOmQ5kjJ4XFoSjQDMU6mAL7l94VA6f2Ep
/O6hYHYSejjW/5yn6qHv9G887UYsWXelOugnACFsbXSGHXEcmVWTP9l9EI6XJqJ9i8kqkCnUP2VZ
tY6R4lhTsUu2vovy9BJxa1SR4faTw5wYY4pNY9h/hAVg9ngk18FHC5ZYsCuWcgBc6FIiBAJLirUl
tqg7bMuacXGXLiY4V5g9l1se6xKmtP5ljdt7O//QilokMMAo2NI9+dNajYvgWxgQiaGtWDSFqvdt
OKIsXxtYbQhEKetmsnCci145jbJi6WL2bzEQW4REXCKYZG7AhpMvqGDc+C+eC85zTLa+nCP8pvVT
ZnlEuGocpGUOmiXvCk9yqbX+goX/zuBRZNMj08iL+PmdJV3ekDveqaZ7KIbjRu5Z/DUcamKn+eYq
lX0d3bpMiAt7IYJ90aFcKDNmUZY987zAaj0a54u7zWvyFhguyXYb2gufXPh9+qcUeCetkrCMOAJj
GmmF48QE+OXslJhzODGporiSXPkZhZljgz7guHtBltj4bbh47uhamcHFiAqfl3kZ9mbJihduajCX
+LSiua4+8yxuvwNz/sksdg688D3ZW7bkpX4zoD+Dnz1efryJrje5aVCFVathvhOnABqIzc3oW2sy
Ta/qUil0z6/MuxW0uMBOINNvUdBrV02PspvNdh1CtFGks22ev7M4QlDJh4PkhPUZYOK4awYyH4Bb
CxnPRTrwc/tdzKrs8u8Vbzg9cVLXOT+erPNW7JH+WgXNsitA0DoodLHzB44MIaHana6sQHYLjgVc
BekUm5iRpNHKcfkPQSvuzc0gHuXn3eFJZJLItyrdYV5A/J+mOzYeL5cXd+ppIxtwXm9WF2CmiRNr
P2GCZMJFabI45DGqEk/VX1iULbh/hqU2yHIHxhG40pkVAREicAVwOgU4OtDizxjUoZy7E9hODQY0
IuQoUq9WNLlj8sG7V/x/L3uhXIwiEUxxQ5lpk55K4aTdyj4e2UKMGNjXgMOhZaPORR7euWF0Z2hP
+ZbvC7cTzKC4raBdS6M0ZejkqwnNQaaQU/mGd2MsTS3A6mk3DwDb27Es+tgbnhLGBmI2ExcjSUJ3
4+58wBPE1iA4adSbJLToNGaOG1YPzuTLw/I6Q7djqPiWLNR7ajcXaxCTKzVQ30bht498SNnNPELb
N5ye0PZ8yqfm7MXgdLrkm59Wdlj3s229Jjz6sWUGtgKkdcMaUVR1dkwRpBRl7Y7DWOYk0Mf+fIdx
AaWbrp7PTEq6g3hG4j+EIzDyLEoF7IdCVFR2Gbhk7LksjxVVbK6aaalJF5XfliTT4Wb2Pla8F+1c
Ui5fc/PoTgOFggcyWRVsRyz3GoEfYHdbvIvOmXTx6B/1MTLuxkgLN0pRI8nBPhc8JMIY+arg1NPR
GUOwO/67nwD46uzkUJZuwcec8Q6NktPLyPxNvNx7WUWN2O5p2aEojyc8knFIgPyqJ/80Xf8BSKyg
bOFhHz6dfE6fPNJVD/p6xVXpDJC5935FD+lpVGhd8JB4LFE7ngLpi4iqnZJXHoVhmPIDF2VvKGqJ
ee9HvKZ37dKB8Ll9Kg+ES+GwgxuSlAWmhpSvyJwuO0pJSl3f1Ov+3F6nZ+zpV069r6XZHpedq4T5
NZXPdfdHPYMqaQvtudJG8c169faqpfJ+JYArJShmMnkroLItMDy45+20e4v5d+Fj2IQz2xYimdge
K4snfRU1bc2CqHoVe2RUvAUpAUnLGSEItkRqcPf7fXMUNMJ/AVBKsLS47P8vZJjRWBnTa1kjFUAX
8w3lW+eVfC+sRxW4ueeTHby+1QlsSF+qIg7i1DZpt4FitIAjRXgGn49hx1rQeTZuRGxN7jEZoKIi
N7/f+esNBmGjqcHPnF/zM16T+wfXTkWaa7h/DM6SZs7HM/i19W36oN57TrlQic7KZqi+fldQxePu
Za7Fw+GXjN97M00IPx/+q3pPFHWB0PaJh9uvZLufvV/vmHLBrvj4pLECFgIB4chRQbCiVAM0TPRH
QN0XwKBwuF6L1pB80Fyj1mbKdQ64gIiB6JYDInJ28Nq+QrlQlxgxV1yUv+SxZemG1T53IFDGspv0
YOG/gYc8kQYL7uUj74KTSXjQlQaWX0qECBSCdVimLuZ+KbZGgQJ+jaOM+tVERpjwmVbPsqvgKr8Y
zneh5gBuXSqNY98niy37+1qxTffjtW1gLL3hdHgK2JcqKthP2El5NSp+VRF4dsxo+zNlQgX3WpuB
0Vx8IHp41WE+8IHqofwv86zLkmYt4RF0JG210kQGQTLvA59YGduJwlNr0nsyQj+tYMO2ZLKFYNZ/
FaOU/7yrulXrOnQxWnu3u1sPShZTLB207aqOY/u/+tF/zrNzYS+CEucdz9jB61VY3AM8n6K7+6hr
vQoPh/yVuRUjm1+mMY+3YrRsGomazTqMnmVkRnQw0zVi7FPxWXpYTeWm56Uw3SdAFs16W+9QbXI9
r2LwmmLa6fdHTGF2Ko7TTFa6zdZQX6iQxApOTNbZ6fxiB+0CXq7vP4GYyaJChdUTKzVP/gJQMocV
iUDMFHQFWyjIh5ceZDEGkzmoabLHLATz9Y2X5eKpWMgePn1YpjqSTTajNyZvbVl7ccdFlukgLS/D
Vaps0eKbA4ouU2xOMqArXlX9BR6aekcdyMsBas93de//bwIWlpPmFC5mNvtmekbMqtkyJ6vW9btY
cz3Gn8AQHVhwBQaO5OiV2oMK2rehRQaAmS+XWgpixAWmukYKlNGvfZ9Ug9fsOH/qJYtrcc5V4Ynt
n4+EpF8lfm5LT4g13kNWSkCTlsxtU6ktQRASjnqMNZPeBy7xT8g+tHSHTIelAdS5138mZTWdR0BT
RO9PT6+OM+TIfeKxBsPE99RoTnb3g/SBomp4EblLPWLxYgE1ZVPIFwugpRBPkNJVCwFWlEEhNp1f
31t2VtXsVG60eREMUcEQr4uPJcnnP8WoWmi9lCRM9bWtbS/dy6BL56Bil2dKafDEqso34z+7RDAM
V2Ww4xNi+5nU8aFiOB65XDdVukQWIfCeXXSe50NvtkdNc2LQXOxSHeVrrfpliOeI0MWh0eZTL+eV
q268vsw853qmwAFpzsx25+ZHo0pbb1dLJNUIEyYBr6nwaG5aCCkZWt4aEJg9Xw15Sa22J5Os4cff
0LfhiKcLAMNP8W2SJt/ZB7iiEckvKSM91PqqzVXgkhFMF7tKJKhKFNm7nb+EOqCG8jP9ZAm6+W/l
f8mVDFuCLNRrKemuFfOBK0+H2lnM4p2tC/a7qrNOkCg2wJptIrbawN/8q7/dXJo+pJYleJ8Cb/46
oX5/z5WcVM91XGOiovtIhucPTXQ8GsKBnimYfVFnDlyYE3JOM81T+ujRDEWVNTrxBu0IOqOYbzcR
6yn4CO17sNs/+r3NrvqMng+nI2Q63ie2HK82BF+J1HPmo+6MPws3WnmKh/L0GV8FwAON6co6kxvu
ngbkn3/weAzaFYdISkgAd1uoZWznyMJ2YK9BjAnAbIFOGw5pswRFBZ98163kgEsiZ33LAeuBbvcD
H6ORCvtXrOLiesget9eZW2avEm9+EszefAcYjK9gjbGss/10Jb/6VUldFQ9/KZVUZOA1Z0HA+qqV
Vv4AvdK/Z1c5UhVSuBGqB1k0rHTIBT3qXR1Y1qBvs1RYF3IPUGOY9yTAK2DUb/UiBDKKD62jwX5U
IJqDBGdM9LXGro3p78gzMrmm9jKtFmvOFWbrguoPa3fgbBJy3kjApuxjwWzDz6FAziMJDppb75EQ
kS+h7M3LFfC9TyYBL/d8iCMSDY2VlrVNRexhSa9IJRGBEVNjivGQGQ2Bf4Q9L2l9wnxSN0cGqYJc
9cPEa8JwnKQInosWZtvEwqvLontqZr/EWCs1GPLgzb07IAIvTMqJWvlEZIhoM9WcgQ+iV7fhrfnd
hyl1sIuve8zqB8j1vtXwH45t3EArCoQGS1Waf33Dkc3T6+q6oOACGOGz+cWLS6CS22KQugeggH5M
eDESa9VraZAhZ8fzrWLzRTkgoD8LVEZHsHiDm/bvVoLB2l8yJXaGTA7JF51rzvHm1iJ1YrnUbCZY
k6AHYkk5sIXxokwIXeQU83hvCnK0P2zb81SFlde+2PUz5mXrs/3EIy/xBGwi2ABkBlw33LY53SdC
TXqV0fnS+RP/eDXM/FYpFGDbZvIbThSs7Y1ECZLo2dfvNDBYpBEy3cbiXIrhIWJv+SoESxoOjZLz
6Sp9FB5SfUODOQL61r/LqQVaqmcRkp1RNNcup1RM5y6kJcxph0Ak5x+gfE5XK8JUyK4FvHctJIKx
mnJuceLlz5HUsGLF4wfq0TQ/EBYRdAx+JnqF6RKbJCoxIVBgEb/eK2otxeP5vrZXVvB5kXcwoDrE
YbEuZBssl5GKulm5DCxzZeiJUkTaidd+kPNVW15zABgeoFTbRI4PaNmCcYBr3g4hqAiW6oMUJOHF
LN49YNpMsz+BhAflwh/yhNoK0SkBnhEgRwyME1TdbvzEDI8f2BEyNj05ulYviHWL2l3mu4yF/q/c
eZBGgN8uMOq3B6PIzTaIxTsTTQpzoxRl6T9e4X7d9A+3io7Fqi0UNxChkapIahEpfpK6a+QXVAST
pVQv7vK9FBECtV1H6v/TlYe56Be7SmnVomywS8QHfly5wL2L7DCsRhsuDjS8cQzlCTWIAegcpaUK
ul8M04vF1SYOFsUUdEsZH3DsFGa6zke3NvSLQcM0JangAwyTgJ5au/Bm8obJcWoMG0cJfRm+62P0
OtwHdynemb//e+ZEpUqKGlp/wo23/wt7U+ZzOJ0SZ31hdKZXgYNnodE1f73VqytAqzDI20/s3ClQ
yfqt4YVpluLrMEu/zxUrqurYL6AKexRTWAog0/msl4EhyPztUAb7bdnMXOnrZfhlNy1OnxlOCSP/
U0vxX85jXsP/cxSwmwZ2Rf4GZOnW2pv9u/qLP05J3YmkYQ7JGuqdcSFj6S8BBU3WjET0h4jVRhzq
Awwjcsu3V94OxcqLO6cduOFez/6olgDt0QUpiHQdWBfXaFpQzny4N93heOk2O35LMbbI9pfgC0jE
1wL/tjsAdSSUXKxwdejp2k+0nDX+IU2de4/diq6RhMxAGB9D2XJq0Sc9eo8fYwGv16GRFaqpQGZ1
4Ey6JfcChZJXI4PNpbCFgLQzbTEDB1KJvhSUgHYPfrX8M/te/6W2+v5G4s42zAI9EdevRs7E5rAS
F/tnjICaabLf6Ashs++pFvB11q1h5u+MLsa+I0C4itcJdYPQk9+1psxxd/TxSSL0uOBohmhM6oqF
9asBa7a2xlo6X0KjhIlhzQP5OFeQVacsOMnj/4e3gBBeJ/fHeW0cv4jaUesc8cuc5WMV1KhSIVDU
8bcMaECmT2mxc0w//Ox4wGDGFLxOnstJCHotph0P3aDh6gP8V4wFPdWDBZdk2viYyyy07xM8jfaK
yomsgEgtfJwOkr3+o1HuuvPHmh3oYiLhMnPIWlyjZM9eyR80R0o+YDPBUkzpdQ1ysKhCRj73A5P4
CUoU6yILcwT3I0rRNeGQj6VfOPRipyscoXjz1L9t2+QxIRAPdjUThHE+gFhA+v/wNCaDl7lMkQOL
YdyNW0gMiktArDXpS1Krq/4Z/wlX67AzKgjwSZrqVfsIyovqbuhrpN9naF5LFHFHScNrOL72CE5S
hfZc5KlbExN0XIus2JXKTPBlFYDhFin8UfQUh/2dZuE4/IVQ7j1+f7TeWG9DVb3gUdjG48NWXRON
7eGH/Z/3o6V8ZDgmqY08nch/IYj+PRMbfpcYDNOpfgT8cPYEgt3TQ7XH7JX2MCBGCBFAr0YNkq7s
vxS/aFO15iMkTGokbx1xQEMCIX4/RGRsMz9XXqa5Tqn7vFjGyMvrFKC6txDzFdnIgwHq/wsXdmYm
GKnJqF++G/8QVAhOzdgNZZaGeVMJaXy8fX+YTfyfzGZvotBNhjsU5fpHmXEUpqGGQerqS9xZ60/3
2z0gWmashd/XAu5T2tBBZPzdoih8wDwmOQKRg8eAqn7q1eqx4DMPAa8iLicrqLycIvjzZib7FwJm
c98V3iIWY5wyw23iWyRGLAnbf0DUb0oouzhSr+KHG3Oy1EKb1FyjCXNgg0FdkM1MHJe9lOxZ/Gnc
rEanSyDE1qNAD1UQzUlMvAUPmRCBLdyrZK1ip/rSconQZriK/ngA53OCY89hbDHwqh7tpQX0z09r
RKDU2tT0tUFVgldRqp3OBNtZmN/lwxw2FHS3L6PEZjKXlU20nrN+gBA0hUXAIIgFVcotM8hyMZvz
pCjjRsD2p+ZV/b8LVuqAgNBmnK/JDsKyx7MkDvWdZywpcF586GKJmF/mCab7iOPAYJhRzmuW/4dD
sLjtf1/6SuPbA9M88gdkQiQPCJhf4q7+pi0tFDstTblqwiNrdmvAe/OnYfBJsAS+eKNCWp0c/ylI
FVFO/4TyryO0wBdf90ajFOVf6M/hIKBND0Q/boxH12g7MPPL5+YTyluHpijGscglNfsI/iNgiwxf
TiPuBXzog5rIH66b6HOXSU7msUCyBAIHdwd/kX5SDSWYnk8bVKqEF41nj55N0ZYjVAmsLe36xkVr
8yelJ+IFE+THxXGQfA0QDhGpLIcSnVxS7e0TsZmKcXYHOjhJND5jt873D2VFro56kcD8qwKzzIi1
lrnA52vsXB8nvieytfyvcpDRY9+bCt1+l/PJZdy9TO5sCdA+nyRYfgMqmPMMlldrFnySAhZPbWag
DL9iXz/huPUzHbA6SSx+CqY4PZGbR2KCM6Yngu/XKZflFpYWWc5VNEJQQkeYX0ZkE2yJMDNqBWBX
RZSLQImxXchivppfTrvjMByhVU6vGCzi5D1NLCmTIZkQ9HZs9m+7N3Jw8VHD1QmOrEH5Yz37ukxM
DSuKm+feAlrtdkMuHOt/a8emYA3xPnd/itTpOxyFXB8AXXqHhgOIPbu0Ki64rdEumVAlqp2JNRD2
o3D47E6yrincv/FogY9ZiENI4v6vv22hkRRhCjFdr5K6salIPB+YvPf1nt9OFGjc+U1AYgmOlp2D
Fvf8LHwQt7RKE59hOs8DOd8+WcT+dw7/igFJchJuuZ9fujSIlR4ICBIXOTCsS/UU59YQ3mNM3pUl
CvpDTMy2XciOkaeNwk+7LqUQVaz5JbClWMsp/56phmjPKXtRz7IGNoMgeBIj+kKiEJsFO7v2npvk
GfWYICOO6eXkx3aROaQTUMwrpZilUoXz3KJyYtBfcUrBpe8WyKdEkn+W2zRCHH40KvF0msUgMZDm
dwKtlm/Yt1PPf85EqYlFoG/BYjcKkgCiwJEiNE2fZ/OHCHIT7vCR9v8fPKlS47aDZmNVWBFYQsk6
9U30W/p8k0pMF27fFoWTFcQMh8XhkENNvUfYpIRvoEOriw+AKrmSWku8/KnBF8uqIDluTpZOnbdu
mQViuo5SYxUDQKTE4YJ1BZftYXxsMJdFKXTa1gcUdIgeNw1iGlxNn7kfT4Mi8h3ZtsYlY2E2rjdi
9E5q7kvpo2EDzFAoDBkITJbbSlZ+f66fDm2nkLsPsvi3CVqvCO5YuBKlexyjqnBlaFXNv3VbsmWi
2+qukuj3nBZHZSyNUaW4a+i11FIVy8Rxs/LX9Ck9erRRu6nhoAjD/cKgXV09v7a0wsDI9d2ee46u
9VU9zqP8n/gmWA1Rn088+H7muaIsPOD4ePQ38diLkKf076Yq2FlQxR/8MMIlmKHbzNnDdv+gomCS
fFzW87nM/sgb6aBIORfDKpjWxLnoYO7fRIU0Cltvkh/sNfQZzW7wp7LPV+q77kC3rwIvL5YrcPYC
/CfuBtjukF857hLarBKUcvwCE5oZ2SJkcMowzko5tXxUDX0x1uiqI8YVU98z/koLiNBfiSmhbyyb
nXf67PgJ5gaOQHHe857dQvS5fwyHaX6RlDswdFFYx4vsSsDZddLKJ4Xqy6bbKM6GYZPTJupQngNJ
JhzaLp0A3U3jpMw7tcKXMUDkVXyQctuJTDYEipQSABvJO86ksPaYAcGMsAHq05nU765z03Wv1oSZ
CB+McbI9VX7F5TQMFUWWx/qZjmwejSIONkUU4vuiJSbi9XRhpT0dX+KkFCsx69qTRvrS0BbezdpV
W2HBPCHUntCpIyBwoBM7Zqv7JyUhbn2UFXFkw5Nij7wGAbnVbqMQ56sYTdQMAsmEgSbuCMQhYp0q
B1P/M4OdgnuL0diPhzU5t3En1Pqe/b6pV5RXFL09BT9qXx3zYwj4U3A9EyyBeHg+Wjn1HABLdHtr
rjzZPu2LEdHuC5PqelhF1Ds99bxw0ADnypS9Sa8cBvy9kdNSe5LOzJo4JrmIFj0YJeTg1++yiAEZ
IaSu/IFjKNBFF5MyKaNRh6gI3/Q48Tczfj6qgNP+yJPV+8JTg482BqaD6DQwaCDSxUb1otpwwKk4
q0gkMXYHtSr1VrNlfVybBzQycV0j68D2AJ41u5e7pCHqkhl/zaOi5Jbj3kqbmHJoYIny3bM/Wbpp
mEsUasCEe1NW+Cc6D+CH7BBZMUNkT8rmaujHXn3zT5wM/eJ6rKACsXTcyfgMqQnB7J0CH6Iv3Y76
ha9vS3TJYVmpHljOxyJU1ITaYguUs7v8a/n/71KmOLMqg7KzG7oA63MKmsvHASkU5O1yvOl5irMt
pTTeUwqFABp/dbGXy6+8IVTTsZqN26yBMnABAotGLNOhCL3cmnONrfuPhyE1/O0PRHeQOKVjjNSr
hLqlzhsAUKiwtgjhI69OmlPxaEvJTdVZKzHedMqYsmvC5wHTjQhROr2iqH2acQz+b0FJ84Pm2LJY
iNA1a/QIIrRUBmYVxph7sU9C2Go7yGxZ/94WCF0RWvP3lmDsrjAMCuCLuSZ86mEoiBMZQxsey+Cr
eHmPAEFB32aIq9TKfZvmeGuhgZCTFRVF5V83NLhIdz8M4MVvbPXn+CIiV58klmvtyyLh/Si1TeRt
9ZwTXq8/5uh/6/FNvBN4TJmeQqQi/3ZvjA+ugiztPJZBVgtuQVUoqxpD7fQjHVtCWavXzQluzvI8
0cYq9621JMZ0vOdlMvjKAIggx8iW5K4Bp36H1HA1y0vP3RgrQeuPHJfltrOm19vArJBg0YvGLXC+
vtboX+7OkgrxT/HBmUN5YUW+T0wL63ZpemxTFRJT76O9kwq6Fn/t+qVYtak9fe2OWuZa0HBTo/X4
f4EBt7g8n6E+fnF2AzhPSCbuyN8ECFcVMDvFZOdAB/vTojb9hZPPG5pdKyNlQ257JU7fmiwO+SM1
J2VIBSzMf/Ekt+mQ/McHX/FYZlAIe0y8SX7OtkJ/ILnJcu326qgwXTl+Mu3C4JE131acULnEeVDW
OUfUzuIQFHt4uo3aMJpHIgG4G1bo87ASvG40Sy0YeADaPlsY77gUkFTJN/PC02uoXScFqosesAL8
prFVT4S0JiS0KSRk/OX8J0khgfOEUo9AHqb8kBJ301RD2pRvQfOE0sOUN6IZunPufHPZo2gyMmbg
H2H37ePxqMMlXwPGuz1LrhByR/tiNRhK8e/xfhBYl76q7bxUeR1aVVYpYZEzr065Fhbc8O21P8mt
ppR4Gw4vivuaz47S6jhD326F/XpWBhASyw3hF6THoJj4sXNQGJN9jYSDmyusCQiV5GzwYq0fkNyk
orwRp8wydTXL3HbLD6fcGVV2I9Ufo2VFtw0Uv6crHbIXRily/0kIR3NSkZusTyYYfvktCXkGp1B7
bnPETYUtRy2TfKq3mzny/CLiALxPzXvy3TomzNB+0t9dt4oqxqpMJ/vIUJSb+1o1ZW/JkXfR6dkt
aKzLCzb4IKbEfDLRPEt+cx34ha7ep7GnK3JWFUMCBq2TCuIZOO4jvnWqK0DqWs4U4cOYB1jzQIWX
rZevf1AI9AatljN64vJU0haYt8EOTh3+izH1AGl8+sgg3Yyi9sicOFOkHFX5G8AcMEO61Ieb/Pai
2JEEIEN5Uan520DIQq2tRbtQ5K0rAbJOP3T4F147dPqbcgoxAMEYBaocgG3ET1wAsPpkocgpLOXD
ujzPBtB6izUx3azaV/6ESlsZ2tFlUb6vLK48611hh/BITLABXty682K1Dn6yNs96R3hmf7rgtRqW
W3CF1J7Yne+YbUn9ENHcKYC/Kug8f3avZVT3/YPMLQhgaJd8zJE+oVS7O7W+OsGe/BDX2HO8lRSJ
utlKv+mE3FU3oyIPSfD3ONoRMQKs2KCARalxQwfIvxNhPH+16u06mq0fxCrB8q0aXT3FY4Ah/3Bo
MwVzVvMCxRG6YFBP8kqTWam5EOtXdMXnDfyyAP6C3NEyWAJ6qlHOuZos8hO0FMSwNhS3rP4dJkZq
6OEZjxE1xKH8WDUx5zUuw5WQ5ibtV1O0R8FJUk6ivdlmiihOMpxrpeabhf3wnAhT0niVCRE9YlgH
8vzUghmWlsbU+Od7oprNilsGMjynmN4gzKGGnnQ7k6DeMaUCK8x9n03xic/7DWQblXK2QqoKEy7x
GfK2738OBYRSxtDh0Yg2mS4MpiwnWtPMA8QpEnyDDMvCTrMN87ETME+4bxVjHPbICuao3ERokz9H
d/zsg9j+ZRbwP9fyAO564KtgrH9NJ0VQ1KueFnw9dZ7pCrmI2mse1qQj67R1bj9rXDaqGopCr16b
ntWO07pvjLjDwks/Ld3B8NMr7aeh5x0KQqCZg0zRwz84WM1ITrFaHgIyTR2/7QHgr2HjoXEquROy
OrEJG/Hav/dN2hhJ9n1b6Lhvjh6NTvc7kXCGgIVluNt5PeBGqB5OfJBfk+qR3IdnZjyxeJxwggQj
T48C+rzjwnPLH9rMhYhzHLrl7kBK9Zdk85DmBcEs4Ku+gdJaZpVzNP85gxt8c9gGEwllFVLqtVkC
qxh4I1+nxoXoPYTfScM15W/fe/9XOEvNqs07hefZcgyFNCOFi6gYb7fSymOstXP++m6Tl2HB6SUl
0/oT5gICE6RTmyJutXENp8p+ZBASO83gsch0ARyozcLLCSeJmwlutMbLzO+QCWIZ8cW+3n3VHRYn
IB++MNXOzpYv/Fzuv0b4htwIweWP6+GM1/USryquPqOC/9d5TTMOLOU1tTUcOcpLkEZU4YhBkVN5
9exgTWRh/tRD/T6gZjUrUOq7O5CBtBAhao/VylHXAk+RYpc5uvdY60NA+QSboZqRhya0rZGSKpcN
QKEoblvfs5IaHre9dvLpAWbIfOGYlFHarjnTrOtPfTHFVKx4mq03bgUleDg6VFzlFRd5YAulaHLK
4uwSd2o3gItg72zafSfMYTF+gdp4stW2xWtl82qdHm9HU0OHiVis2xUmKR2WszVAMlIQOyP1jH4W
kbv9gZXnpcHaCkHIZEeq0ERWB43dLI8TuiEud7PjnzxGf2rHBTm7Pd7NUCxVAEmwLyfnyeX19boO
ZxuvdmOmnmw31E7N7dVpD7EI/TheA8hrIbIa+OfAniJtP4yo5hfV97BXbHrrkyc4EdDqwWPY0SPo
BXHYdLQnJM/3GWeZ9XdrURIy6g5iJDpsMLY37gEiTQsKdsVsvbsXB2o7YXF7Sn4WPFVmjqo2Hsrj
rkmSY6h/WuR8pVbFeTPQmZx/iI1ruhIXfeJqaRPJLVOcv/KF8PnbKPOe521KQ9shylq05KIOxAdJ
LJ+cs1B0qTfx/04J9O0wHYWD4Na4e51+0kXagiVbe5qPnMqSxaOnFiEmMSDGfl2PyF3r4OOLHFBB
eWf0u6Ty7WLUAgmCEJQKk0TXVK9kAscU8XZDFCJteh0yBQl1KN/LBNqLE/cxMGeOCRPzo1bg78ks
VTh3bRlXD6EEQSpTFgmB9fYvCqfhFA+veBHogzMB0sKvmSSZljlW4yH8YfezS0N0eBHzrohFmyiK
E44QCZJqF1cEDQnMsds6q8u+8/bqWStB0PWEDxcfJNp92veLMp0r2iHYXuviscoA0pafE2ukZFMZ
1l6FWP4yI1mIqv8JLrIjMB6cbHYjOHlFkQ2w+Bok2SJNNADpO/nhmU44O/JdRVZabo7arOfvn0x6
awJ7Du+AIHtpBXwN5dHGQO5z2r/Lj82WzNSZedyLSknY8dx0dGh8ceJLf0Z17nxgu/InKNbNAEz8
urBwwMJbgUr5xRDjbfv6RcdtiEnwhN050b6TUd2w0772siuBskeCyy345XjOCK2NZVQehkHoReXO
R4IGAYCHYbltFuOKkQoL2O9sequJXBcymrQifEW3OY/AAleeXZPIJCrSDmi3ZiaZ/J1GVq9nutTT
GftR+3RMTZVstp2ctTINMR7vKcMBE5tv6q/FvLenbfhmIadACPgVCTTzVCJtExmlJ7dnzhSFeSbJ
jl3Wduchtg87agtL6cXh+UgiKtFM9B27andOjtVHXh9g8mOxrP3JWQ2f1/h2aStb1YgmYRmAt4r1
b8u8mkck/OAD598jqdCP808gYcBh1xD/NtyyKD1Cv+zLzaLGO385a98qVm8P4I2NxruAckFbXkkC
9o/sruN8W1IbvVY9/M+v4xB7hBeTIQeytq2LmGS65R49RKKwKZNQGJxbNzKtQtACItnPscoQu6pl
Sz1TfQ+Zg0uZnVX+fAEGE0QtqpT1Pe3HkQIbP6BoBI5qIoaOWwFRDDrnRpBAX4e/DyU93jhlylxN
ysePlFISJJD047D/EontjB5RVCuEeG6pg0rGHpEyVQJkfU3NmNtbyx7aOlsPmf3m/hkMwnOKDGgE
qJM8MmhgxwlOqyF3zhhjiCr3MovXQzfcStZweb5SWNyKUUodD3du3PxN21hGUCPxq31YwQDPv58A
/mOhYnk2Pu0YMgxGcBT9lX6nMnagzFIl0PZN9wrBqQJFXS3Zpg4zZp79VX1MwNgethTZ8kI/qrMa
h68G30gcCQua0KhS+esXwzbxwBNesmnQUWq5LcemGClA7wXqIWf66JEQVB/JiNuMLyW3cARD+DKA
Ebttd5LXGGweDli6jPN9vK/+oirEbtIYOFnSkFbTFyH8jTyZiWSWuPKdVie2QaIEnxU8BS6A5zHF
/3eyL9E5iw5coETWLJaRAxejyO2W4BZHr1exm37dwGM9WO/Hnx75FeJiP2bE2I3+/Z/wgePlmKik
KSD5tr+2I5AAFLQ2ugTJ5ef43qu0S2dtL7IHQLGgG+zeEZy42twCs4Q2IM30Z30Vv39H8gpbfta2
anyie2FeJ/6ODg/yD/e0qVYmKHD2sr3blCWoM5udH2YpJxZMZQ+Op/IP1OaxuvQtmODa8viJiOV7
DKIQ4kDkd4TiSVlLIWiAraFgWcI3nrbUq5EjdyFoj4GpYAEaZdTjPciaND4BK1yFvJgedDir/svb
oW/QkzQyzYqjKbAMaCmJ+NL3YtN1SsV1/MjQN7P8CtFf2M3mcsUkD+irJ+JFqJerJQU/kXTWdBvJ
f0/33Iq2hERfJtyRezsvbQOZz8zWohQ2RBixOinR3Xt9Hw+PVgQtdcZubf18DQgXQ7ChQ3lJrw84
RWRgfXD3482B/kKGtFSj/La0KETCAtriaQhynzIepF/YuYafW95FtaG3hUR3hkNB4zKDV95zTx/H
nWLeEvQVXLEhR9tryGSPjTBNuoXnj/HIvp34EnCHlVi5P70RSFl6NRNbSoAEY5QQaPAYTnLO9IDz
RuH9An8/1a8Zp3zm8Vb55GvaZ0Kaf4hEkGA1ZYrELeA0OhXsiSqcRePs/ipV/8dEjV92fFqEb0wB
SrOgYnY051MSLG5ZkNWy3yeV12DH6wpUSPa51z0vWQiSHkUi/PYmEZmVhJopZBZws9qY7oLOWi0i
cEXOzXp11vf4UFYAceSLvkq5k4hacqoqClwPt2ALMxC38KmWSwW6Axdi9UXQBke8FG0P8jKovHXn
IkOJOwljcuvOCHsLjtmwk7GSFCXkoW6L91UODbuNT0qbNFUqKF1IslccB7asUfH+wrE7iJ5g/1H7
tW24pEAuaW3G8B/ffcZdQ7wN2NXo7R/NIaAcx8tJPx2hArwatEherZljHHP9XQ/G50ZAMxbYcItl
QB7Xt2rHyMnduaendK+VfbYovKDLlFIrSYUmDa8Ob0GK83m+KDazADA8h4vR2a4+NjmTl0WnTxKS
QUOatfrSS+ovDY7IyFduw5PGyBWuEjgTOgUKidlcOZPpscNYgLER+BOm+Ya6++EHiaZqdN0zz2gm
UAU9F6HMbgKcb8R2KKhEuuGYBHzx0XrHi3vvlFhKn/BgDv5XY1CoCrfFzqrNQB2/T1QQNzD3e0Mn
rlApIbjz3nOa8oNUk7HTbJmLEmpHRrdqK1AqWqzMFwQylQNabAa6OD/1ktyns15yIroOsnKloYb2
lw6o/afedKvYinekpaG31W6EQaU/qLO5en79lFtxo3kxYSeN8M5ul0Zlzt3HMXuvBGPxOI37bRdQ
XS5YIM9YQy6T1vl/KCPMf6iwOLtDewK76MVG8pM5etdERgSwcKilkOjb/zxcbKbkPlqmv2XQEdGB
GgEuU5o0efszPTEI0owABF6IzdWKSc1GgARYuN02ln5anNhdI5n6xQxY3vH3KWQor5y4PgrAbcLn
xp7m/5g/PbO96ddkgbIoA24v7lfC0mUe/Lc38sd3cbLxc3aJrPL0bbIecNwdhIgM1lOMba3tO8jS
2DjydtGUujL0fyWDhbAydZAFODE37VueeaD20Mk6lrJN5jm0ylEhxq0DDPdDmdiElXreDm8D/kCB
Sf741/rP4m+FS/CFZXg9M+3EMSEMl/oBKUsKlqd7SnnFoo3NNjbwjO/B+Zn5xFzDtxKBznK9PSmQ
G56Fxfh/SlncQHfdarjuxDbyYO5UyymhDZpaOEdzz+wCk2weVWy0qCdurKevKPb2n73I7mJGxN3R
tUajC8X86VPmdae/hleG/wrS5xVHEzUfC6OB+fgyI58K+CaOh5Rptcjqow1R2T9EpYRw7hHF2TEq
Q546kUhQzvgLHDPoy4BY8zZufxcSV7q4zZ+RyZ0/jpZAbFCjCi0EfDdpBrYsDst+OVfS6I8be/pR
xdhuUX6E2Dz0SkiebJr/ALIaRdWFtW4OyZ8EKymZthSVML5TtQtHNjjzl6HYcZBSunVvPEWUR2LK
O0XF6xTPCiCtawc7FjsuEesSUeLo2OnfI01YHnHc5HaNO1d1oWAVR4W83iTNT4OQtaZGL6vg6mSu
QhDuvaBe6iET19upi0nzHTBHqaPyZytS5sNz0BlYRN+zAWI4mabn7AywspbmXtHM0OQB/WgBY3os
QNxoStc3iwEmqKQOoYkrYuB7ERTq47bBx0mF4gD1KXTMJLU10NdPff+E5q6GKykCTR2LRDsrisSe
onRnxqz03sEN61ZuYCmYL/Qv8shyjj7BsLosm1ChchJYg6SBWkzc90BbVy58dIOBEt1eImFwxLOA
fj1wfpGf2q2LqZxPvconxG+XAd2AN9Sm6OBF3t0qPh6l/C2cwZKZhvyeyEc2wH7d5BHsxO8MuBgo
mflcZYMMKGTP66STl4NqlECvGKftD67JfHAFhw8zO5is/ws9l9cVuixKRitLD6726WNMk/P+3ZNm
XaBWX+teMQweiQ7rtdC5yDEEcSN59hJN/47pVILl6YUtgm0J42o9mHrwhihhuy5uRIuI0QBxNZpO
chJrMlCj8qOPHzc1MVuuerCpshtuVqz7QkYoC8udcvBuH0wNW4/ncZ6sJ2SQltuf6ogyiOzMdIcO
Xv09VvoA5OqtofRKPnGYNZprkZ7nVL6O+DuBuxBmgEcC658v3FqzVsJmh2vIPdv2KNTNuGT73DWv
lpaqczWHzPHlwb695+APi/7M9juQg7/fwx1Q2gzQSE5CfEEuFeiURZ/MPm8FYtgeENGkjnt+Xc71
OGLISgOG8q3UDLwNGBRvB+pwzwJIPijrSerfcJG/zWf8Aqx8yfzq260S2QYCCMBMbzwL4qiKbH63
3yXgT+ybBH8fjzP1w1z5YpOEansOobDkh5Xf0AyN16DrtPUxN+A/cXF8EaZobgh72kSTraL19+QN
bAybJU9t7/we0HEDH3MIeSTxfnU2oCjaqtL0eiMjiCnU7S3owv51J+0RAOKGJBJTPEqzdtG478r/
ch5AbOMcbbEi4tytM8mYta9YFQ+4yvO2HZ9IytvKoFjashF360wuLDtfj1mSH06HzR7mGmVdY3ov
rfpoYaQLU0CavjE5YJe7wQzCwNz1yUAbLi9KiMnu70ex2uKhg88xTBVZZDfOAF1yYFUFM6rFQcuc
2HF5NX3IMBQUHlRd9JbRy39UPgvMvmiPmQpElOTjcrVoZ2+ifhUKVU0GazufRfCiw8X6Mlz0GIsv
bBJv/C1NvQDhKRJHTMxl7mZyE0bqmwWDizR8//uEbEUVnHJGA/LfX0AtSUpa9l0751vMuUrEu+XA
l6VjBBzPlwTETJLFS9j+yADFrIoICKwIM9EBqtTu8Ns1+ZZz3gWJysEWuTgE1KsnWLQ63z35Tqqn
5odm+MIheOpcUA7/m64YLhMhXyqAUiogxMESlGr1iHfOfhXFSH1qLLeBWvBjRQ9A+AO3ENkeqPr5
FvewfaPoQT0NEejdhNLIVUawTl9exKgTFvlJdn8HWrw7Sf/MFTG378Ot9M2L4anCuRehimgDW2+Z
miDVlkOuYKwfpcTGZ1oEJ6yJp/Y6EgPcgFcwHPz9emZOYofXuVwUIptdoiWu6gmFqeHNWIhAvyPV
zuezipQOffcguoebz1rJJO5/AZfk+b5b/i03xd8e5cRilLseDGb6RtGUK2lPp5fhUsbbTelrlDVz
wr9KfeUfeDmcIQFOLprTShQQi9oHAwqpFf2KK6t/am3CtCrOI+FI7xltFakkRdgY9IVa14kz3Q1h
aIKg5b1v8KPJ6PUj6/KSo+yGeNkObaZVkg4N/+SELdCjcySn0zGwgX+kupRf/wqZIqmAQtDn52TG
GBp4k7MFDizEyKQE+9d1cqIMNrZ4eZ60NMoXgUTiXwDUnw6n9hEMsaunSrkpyptX0+8XDTxoZ5w8
KS9Pyye/LXh1jGiEn68lN8Iq4s7TpZCP8y8/lpSXm/s6/zPMekj+aayBVijUWLZN6n9i9dg44qaa
sHO9ugXUQXtQsoPvC1xGMlBeGVmF9d5sg5PD9oETiBbScvO7dQ4oqg+I1p+QyZQri0/mQ8N9ihKk
QNEMS7TvqWgjQIq40lzZEZ7San+UtwfL+K5QFLoU9+dCtvWQ6HeO9mXxfXziRBGki4inNG3Sf4sh
pslaWCHXVPIofpukdG0EDTuDIzLnf6diFonWe/ga8sjvPi3/eHjpDFKA3Jm1OKPTLkaCr/qpjCJt
/tjzIFij5/bLJ9rK4ScMXF4TGVsKvtWE7PXi4oqYrIQj/4sUT9vV/BWSviZOxA+lqt1SDC2ykNdw
4cnz4Pe1nkUPMNE87VgUMmdI75i43Wr7BWBuPkOwF5I7xX05TAOmWD81Rpw53UeXCON+td99hPX2
PXO2ZZGy3V5tIABLi1rS+xWc8VgoXGyNYytyutfDMuXEmk6ODwtd29lODRvdeS4Xt4XzAdasXiic
IXpswthtltggjXN3nDenB2eDO0TEdNmpUqLMvpGIAkkKrhUQKCt28U5vVlWPCziLriaTRxZMinBF
kcZXqRVZ+Coirg2OWCjYPCjlhdXp14eZhDegu++tQxIo5N+TFMhfVm+japkJjsfIAiRVizVkvhVZ
/C3SS/eqKDGHdS9VClYRc2D5umYJhgw/TJYa3GcTFC91/Nyz/y+wZLMUPEN8/9+hkfybCBLVjuWG
jtUhQDAgKd64Tevc3Ok5Z7mLOH9jhvAAVWZfmkMbAIAeoJTi0JaH1w9lavbVdvTyKEjLXN2ouFJU
n/nflGAAz+6Rk9RQ1mAs/dx+NYrmHlDGap2yKTMHP/f4WdPM9SVK7IMYFQOQk56Vyf7L8KXZBUvq
MQQ0VqMw52VLx1iOGB6XzSmfNnpj77sO0VZlj9yyjnsVxVDv6/81FnXBJxw3eR9wky0DN8Q8Mx3A
2Do0Bx/A4FY+jZfsLmEYkJUa5oLWvOlDkgEcqd4SmWewgv6n/NQujQODYkXMEjuZ7113T6u/prEb
F1LsKjPnw6P1W7vfyYFdVEMVb8dMjvV9Z5vK6o+Vk5GfcC4hjIZBZcEDPS1uKT/WaoTv/LT4lZuC
xa7Q9AbaplmxZSqGrhrfU+JdpxoGMbJFM5e0aOZUrLm3J4yAUo5UdmRFrGhN0/XsxbnfJ38WfgcG
eFVtO3N20OVTSSsCH6dGe0y7C6LoqeaCh7dD824Wt7SKrkIaBrRnRE3i4Ify/tOKbL9NK77OXHtn
IX+gychU0u+fPjy1HUkWlYFaKIl33AiDF02wSwCjc/rOB7dO35pAC4aH+OHk7Tg6vooLT6WLR92g
psxGDFH2YKAm7VcH9ReEWASVPJmn9VRznlTQKTKl03lFOyxpioNAIrLh0DYwlCBjXYGCvOiEzplo
o/y6aOK1eb/EQ9T1eC8B63xYPSsKADoH5ee8yhxmVALTIA1dhn8qp8bBEvkrQjiZSCZ4mxZwSyVK
GNCUjDYUHn99JEgcl/efbJCV3+fXbg7IA6sKhZtgSqlWRZlvDZww6IGR/7SjvUCijsAXauLARHKD
nlMIsS7JwIeIDzroDbpoHVR2HM9aL/zYMdfQSOGpXmJ51curblghJ5C//J1xl2HKKc0AqTjc1RQZ
Sb+5WDZG9gazyLmjZEkjYJeezbnp2jQJZfb3J9cAXAXm04K2QJFEb+u/MqYkdwMBiBSOwcyGJDYJ
SBFC+8fW6yjbTfGtUMAHGWuVy8TzTJrGdA42ehOn76b+imspUZQBtjZP0BVr/dRmBWjO/46m5zKf
nmqs7/f90UhQyTOXFtVrTyRgRTRkfYye0IQAcZ4xDT9BEtCumreitonyZveTSZPl6FKQwLAcqQ5C
icMahU+4yAyVI7uVlusTY/+SAz0eBdGtdZAusDc7rAntqcyPnDP7PWjF2C55w52pQNTtQJORgEhJ
LbB1yokGDfIYkMDdsAPL9nhLsv993nr2eW1BPBYJlxSFHfboT7exS14vZMHhKp2xLS2E12KJYCPC
0eJYTXE8YEXUHMdYNfc2u0N3499lhhl3BdR/Rqw2yLykp7TiAelS1FrknIi+YXj3GJsEgy8goxnG
7Wf9DpYGKJKDGxGZfa27iIeN23FAOp5lNRWjsp8A73c2qUDG6AzMKy9k8Z9+ekwlW4yKkdiB6hR9
z/JO8X+0I9G8uwv5si9MN7b8N7vx3NWXjgz1mCRBEGCgGQb60D+asBnSMfxiiIWodIHdf9gZ1JlE
pV9aJWuY8gYY0BDdiheW4SGgJzAKaeZSk6NgKlHZ4EEF3OtUvFYaQC8YKbwqsakJ56ngg9H+blbl
k/2fW974Cvkp6pkk/RLuqNDHrMHhlon3iv78gdhJNmZhQU7sXi8HlmiRFkqbuAPDEsZYrNOQohkM
jRSEWEWFV9DtwoRyk2fvNhd6epsC+C0w8drnVN/ywuq26uyPolkw/5wqPyQQUzqnUX4Owr4Py23/
WesZu20aI1zExt+3xf6XqLmRnip2yEjcuDsTiwtOpDr7ONSr73EvqzS/FTP9rmDIadv8V5s5XPIq
RWK32uvkHDJJtJJd+DWwmlvmLN9STs3f4Su84N5+XDMXsUTqCwApI6EjC3RV90tF4Cx3uYO9qne9
INa13/qXumjoVldcIf09HQ8HQV2ELd5NEJNZSxLH5yKkPGeRffNCAP9OcDleYZFCX3x/8EjRPMJ3
RIn0c7mxCBIoe2ZqUJf2EiQKF1rrRTY85B9akgfOThM2GwG5QWW5wiUQvILYkMRc4ibegwkHcBod
DdzRiQh8UcjSnP+jVsZ8iVXMc/h+nX4RBl3uDGPn+1AfdEnIc0tFGo7CGWiHwXjHGB64S0+Q5ySZ
l33jwe+PeYx5KfB4UI3Cd55fQFcG/F9njdpqKJNsPaVItN0G3cLaNWYa0rGxPRWhpzUGN/N1m7RX
UuCNWJGdV2k4OdqTC6nIAkx4c5HxRon+PF3ugM3B3T810kzcxxaldqPwjPmvMRo+7nd0bSIik46V
F1pRg1V8Or2y9fkZQsUnoHUdINx15LkC622YmD/Jn6NjFgLEiXLAVST5jxasL34NG5QOaHiavhOl
FNZVdcHuRgP7g9ZqJNuEQ6KNQ+T4pMaKBAMZNipc6cEaeIV2XIPLKBoyshTghFloqd2ksJWHFfmI
v9LyURlzDdk1CsX6gSdfb0WBzQXeD3ZTSWOCu52BcAgxca5rCcucmBkmw5llTUzXdFY0zhuv3gpd
e3tC32z3BRrxosKkTajSg3RQVF9HUrJPoRK4CKaSviYFDB9f3cnJ/GjN4MoZFAtEr9QG+uPVf6wu
4NzoOKqxPeFDm6/HPfFg0+3H9M+w9xy04C28AASUa2Di8pIM6zKJFK+TisIiwa1nVQ4l+QhCGpcQ
gjtXcbYEk+54wB9+l8yxmO0wFGufAaX0VgkKn1+VEXw0scKKW/99CnBavSnLFxyn0pXhfrrnRF6H
pJ8vIOnoq7w+8x/XMA20bpwBLQJ14yteg7Vo6PfwcYAzP7qhphuj2QQS3/wYETPoYaNgfIIsa9T0
QaOfaiohClErAxnmWFJ+h7SU+19fkeKbuCkw0NV1thXEU1Ns989l72i45JvQwkSHrV8EB9oJHnqo
lyWnfRqXfI236dscHp5KTY8Wa3by93T5DQjqY+FuDrpwaRg2bSkIq5PSidq7WB0GAiBMdjMyIsLX
ZfuYi2Slv8PfJGyRGkH9p/Sze1qgsYuLsRmYzHpkNs6Vlq/jTA12jmXEf9mPqzfjk3ETxRRKpUDW
n9HL3VQfAAzV5zWAqabHWEUZ5iOPYkbhLEBobLrWcuMGpbxT/CRtFulND7FPDd9V5Q+tHDqoS1Aa
FHv8GKdB18K5sF+jAOZsll+LnD170R+9OlrwleAVYPmwXlst5S+xSqGhkM1l/PjdFqa+l6nATv7Q
qnS49AdY8A3ZYUWz5aEPp+gjshcE7DkyIkY8lJXBBr/uYZj7UmAXt/6ShUwpDtz2eNL8Tn9VIRGu
y2jqAKO4M9kqOYZm/2rNwn7ErrDuRa61rMcB3pkKFuP5C1MEEipWg1QsP/tj9p0Jibvy67UQB5Va
sTGUuX7XoMnkMCiML8tN5c5/Tb3281DSj0//0WP9vVT5u5YNa3iIPJFbbx+7SCGF6uoB5dlmWpDp
s9kbei8o9DO6YeolZav+KO/yXXRJMoboYGvEevHhN9L5cv0NYc15/NDV1fu9y8PdGvM7QsZdwzMp
BDIO40ww8Bvr+18HyJsSpGcs5myS/jEh4XmncoxhNip2bLACK7PCYd/l9o6q1938pJvkib0jPE7E
G+4ZROSbOjCNJZgyhhb2X1TJvyCt/T90TCYyJWta9zSaw7EBzooyOWMy08iPsA2voZ5fVvt4FPqM
rA8cV5ZKeS1nwHifBLBmaiqTRV4H+AscamtOwClT8/v9gR4X9YqYjTwKiNJYTyYsC7m6/rkR6Alb
c/Te2GtO6KIJjj/2Wffzj87hSuFLqmHbiE49eumOt8WZvYCjMFSryxism2yC/lDFUssIuGJMu/HR
dh6sf0QmF+ineULySJdviOk8hVc4xOz9J35/S7PKTdKpnloa4FkmJclkfkrlYaSn3RWbpJ4CnyUG
FZylmiMecVoba+sDtyI+5qJVp6L2I5ZucgJuyTp1OBZyUs3mndg2sSnhdEzff8SOlX6LJu1nr9/b
r9MUzLqkm19woTI7W1H61/aRIHEXq3b3jegOQIJZpkPtlhK2oG0OhHMG37elEJmazVYY8ARfQ+WH
Ory64f6v/NZfX8IyobbQT3VLKwKWnCTdjCOSaIOlzBk1F/u3dbON3BrRcj+OUlZ7k/IsWDHXdv75
IJnVi8SdQVYeWXaM/6cvbKymNP41spimG3zKL0JgdPrLIP3/6GtmS6TPu/WcQleSZ1ZotdlI5sEb
nox5CRWOR7WCfpSWWCuRriHRW3Jzrw9y9vJn6bEgnd0+i9W2ANVBqnPVm5r3rNICdAsdLsSWTEdU
vWtvaMig0iAL+hfCkHazHcGdc2MVqagvJ7AwDsDVFA9mkafV6gM2zq/HJHD4mGmLjyZ2qnBNkc9J
qSAoE+BFaRrBDXg1kX/P7VxnlJ0vgjZg2IsAGQHFVFzcYoAGk6gl/BC0cgw7yEsbGTk4cBrjlUwU
NyxWASDbHCrQpz9UcMr5ZgC2cHcs5UZBahWspTSn3zZ6Dut070dsttQmm3M2+Y+UEO+5Yfcaxng2
MVrQV5cHbhxd1/smWaH0alNhowZaV0sKKki0ij+rnI+PA1h0xkkQ1fN1n2W9eDfEL+OCfdHyRaPy
hBc8DXco0FW5pEhthJPcXQrJFgY15gHxOPy4oD8cafauv3XW2x0sS3eGeuquKfobA/Nqn/6XGIKx
aVV7xiSqL0lV30RD5v+zPIwVekxseeD6BxjWZXO0EEst4zZNj7UuwRgozWqNtWt/Ssr60jLVj+by
LWD/77HKjAGqT2Nm4SoKAFzFQGqWgC+0lh9GiLRAxwyH8sYqgB0PAsk26W8UXWGqooVFY166Zmwf
tRoqHMSkKaq2b+DWl3+3q8Qwgygm6bM85T4T2HPLXticYnaCgRLLDLmTp9AZl50rDr2QJ3M+ICOj
rS31MMNGNRqDXj/kmZAlG+PXQ1gMWIKbUw8GGyCk4vNspvzsfDY8EgHbvbF4zmxbx3BVN+sEsZFd
e3FCiu8CpaKKjpwm7eZWO05Vz4k5gw+NTXinhUMUQHV6kJXJJFOK52AiBX42zhyRv2zxLiKTJEyn
Htlx+ViX/cTwoD29nKQfNNrmR8SGCtltoFqPE0YXkoOnfqb66ufKngnxEG7y3yRVF8M4enQxMwm7
91Qh9eAI/J0oEK10iVQEF1QtZ8chDxT/Lu3FO7+EiIUSpzs3POR4QMUusFwvpSCMHSWgOr8VpgkG
RFR+NoAxFFxwVN3TdkuuvYOg6W0UbIJCt5+BZ9gj5n3k22zIOSHgZVHhAhViI7BV5Qugp94deWfB
I+BwckD/dZcep5g4he6lH2tYcFt9qEryqtZSdeU8PvG5a7wFtykhf4E0GvhxeK9rCJwJHPUa81p/
ez1e0/Z0hfiETY4U/SNrKIf+wsZr956B+ZYaapwe0r3ygFQhazgIhxmiGWMLC76vfhmjbh4M0xAv
+5xriIUTHzdlRQL0ubltCYM/su9HDYvBq8g4BLH+NW8qAAXd63/0V5LHf1ME1ubGYCiU4lxRLevz
2Q==
`protect end_protected
